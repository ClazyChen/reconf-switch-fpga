module IPSA(
  input         clock,
  input         reset,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [1:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [1:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input         io_mod_proc_mod_0_par_mod_en,
  input         io_mod_proc_mod_0_par_mod_last_mau_id_mod,
  input  [2:0]  io_mod_proc_mod_0_par_mod_last_mau_id,
  input  [2:0]  io_mod_proc_mod_0_par_mod_cs,
  input         io_mod_proc_mod_0_par_mod_module_mod_state_id_mod,
  input  [7:0]  io_mod_proc_mod_0_par_mod_module_mod_state_id,
  input         io_mod_proc_mod_0_par_mod_module_mod_sram_w_cs,
  input         io_mod_proc_mod_0_par_mod_module_mod_sram_w_en,
  input  [7:0]  io_mod_proc_mod_0_par_mod_module_mod_sram_w_addr,
  input  [63:0] io_mod_proc_mod_0_par_mod_module_mod_sram_w_data,
  input         io_mod_proc_mod_0_mat_mod_en,
  input         io_mod_proc_mod_0_mat_mod_config_id,
  input  [7:0]  io_mod_proc_mod_0_mat_mod_key_mod_header_id,
  input  [7:0]  io_mod_proc_mod_0_mat_mod_key_mod_internal_offset,
  input  [3:0]  io_mod_proc_mod_0_mat_mod_key_mod_key_length,
  input  [3:0]  io_mod_proc_mod_0_mat_mod_key_mod_val_length,
  input  [2:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_0,
  input  [2:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_1,
  input  [2:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_2,
  input  [2:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_3,
  input  [2:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_4,
  input  [2:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_5,
  input  [2:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_6,
  input  [2:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_7,
  input  [3:0]  io_mod_proc_mod_0_mat_mod_table_mod_table_width,
  input  [3:0]  io_mod_proc_mod_0_mat_mod_table_mod_table_depth,
  input         io_mod_proc_mod_0_act_mod_en,
  input  [7:0]  io_mod_proc_mod_0_act_mod_addr,
  input  [63:0] io_mod_proc_mod_0_act_mod_data_0,
  input  [63:0] io_mod_proc_mod_0_act_mod_data_1,
  input         io_mod_proc_mod_1_par_mod_en,
  input         io_mod_proc_mod_1_par_mod_last_mau_id_mod,
  input  [2:0]  io_mod_proc_mod_1_par_mod_last_mau_id,
  input  [2:0]  io_mod_proc_mod_1_par_mod_cs,
  input         io_mod_proc_mod_1_par_mod_module_mod_state_id_mod,
  input  [7:0]  io_mod_proc_mod_1_par_mod_module_mod_state_id,
  input         io_mod_proc_mod_1_par_mod_module_mod_sram_w_cs,
  input         io_mod_proc_mod_1_par_mod_module_mod_sram_w_en,
  input  [7:0]  io_mod_proc_mod_1_par_mod_module_mod_sram_w_addr,
  input  [63:0] io_mod_proc_mod_1_par_mod_module_mod_sram_w_data,
  input         io_mod_proc_mod_1_mat_mod_en,
  input         io_mod_proc_mod_1_mat_mod_config_id,
  input  [7:0]  io_mod_proc_mod_1_mat_mod_key_mod_header_id,
  input  [7:0]  io_mod_proc_mod_1_mat_mod_key_mod_internal_offset,
  input  [3:0]  io_mod_proc_mod_1_mat_mod_key_mod_key_length,
  input  [3:0]  io_mod_proc_mod_1_mat_mod_key_mod_val_length,
  input  [2:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_0,
  input  [2:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_1,
  input  [2:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_2,
  input  [2:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_3,
  input  [2:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_4,
  input  [2:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_5,
  input  [2:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_6,
  input  [2:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_7,
  input  [3:0]  io_mod_proc_mod_1_mat_mod_table_mod_table_width,
  input  [3:0]  io_mod_proc_mod_1_mat_mod_table_mod_table_depth,
  input         io_mod_proc_mod_1_act_mod_en,
  input  [7:0]  io_mod_proc_mod_1_act_mod_addr,
  input  [63:0] io_mod_proc_mod_1_act_mod_data_0,
  input  [63:0] io_mod_proc_mod_1_act_mod_data_1,
  input         io_mod_proc_mod_2_par_mod_en,
  input         io_mod_proc_mod_2_par_mod_last_mau_id_mod,
  input  [2:0]  io_mod_proc_mod_2_par_mod_last_mau_id,
  input  [2:0]  io_mod_proc_mod_2_par_mod_cs,
  input         io_mod_proc_mod_2_par_mod_module_mod_state_id_mod,
  input  [7:0]  io_mod_proc_mod_2_par_mod_module_mod_state_id,
  input         io_mod_proc_mod_2_par_mod_module_mod_sram_w_cs,
  input         io_mod_proc_mod_2_par_mod_module_mod_sram_w_en,
  input  [7:0]  io_mod_proc_mod_2_par_mod_module_mod_sram_w_addr,
  input  [63:0] io_mod_proc_mod_2_par_mod_module_mod_sram_w_data,
  input         io_mod_proc_mod_2_mat_mod_en,
  input         io_mod_proc_mod_2_mat_mod_config_id,
  input  [7:0]  io_mod_proc_mod_2_mat_mod_key_mod_header_id,
  input  [7:0]  io_mod_proc_mod_2_mat_mod_key_mod_internal_offset,
  input  [3:0]  io_mod_proc_mod_2_mat_mod_key_mod_key_length,
  input  [3:0]  io_mod_proc_mod_2_mat_mod_key_mod_val_length,
  input  [2:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_0,
  input  [2:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_1,
  input  [2:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_2,
  input  [2:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_3,
  input  [2:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_4,
  input  [2:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_5,
  input  [2:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_6,
  input  [2:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_7,
  input  [3:0]  io_mod_proc_mod_2_mat_mod_table_mod_table_width,
  input  [3:0]  io_mod_proc_mod_2_mat_mod_table_mod_table_depth,
  input         io_mod_proc_mod_2_act_mod_en,
  input  [7:0]  io_mod_proc_mod_2_act_mod_addr,
  input  [63:0] io_mod_proc_mod_2_act_mod_data_0,
  input  [63:0] io_mod_proc_mod_2_act_mod_data_1,
  input         io_mod_proc_mod_3_par_mod_en,
  input         io_mod_proc_mod_3_par_mod_last_mau_id_mod,
  input  [2:0]  io_mod_proc_mod_3_par_mod_last_mau_id,
  input  [2:0]  io_mod_proc_mod_3_par_mod_cs,
  input         io_mod_proc_mod_3_par_mod_module_mod_state_id_mod,
  input  [7:0]  io_mod_proc_mod_3_par_mod_module_mod_state_id,
  input         io_mod_proc_mod_3_par_mod_module_mod_sram_w_cs,
  input         io_mod_proc_mod_3_par_mod_module_mod_sram_w_en,
  input  [7:0]  io_mod_proc_mod_3_par_mod_module_mod_sram_w_addr,
  input  [63:0] io_mod_proc_mod_3_par_mod_module_mod_sram_w_data,
  input         io_mod_proc_mod_3_mat_mod_en,
  input         io_mod_proc_mod_3_mat_mod_config_id,
  input  [7:0]  io_mod_proc_mod_3_mat_mod_key_mod_header_id,
  input  [7:0]  io_mod_proc_mod_3_mat_mod_key_mod_internal_offset,
  input  [3:0]  io_mod_proc_mod_3_mat_mod_key_mod_key_length,
  input  [3:0]  io_mod_proc_mod_3_mat_mod_key_mod_val_length,
  input  [2:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_0,
  input  [2:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_1,
  input  [2:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_2,
  input  [2:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_3,
  input  [2:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_4,
  input  [2:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_5,
  input  [2:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_6,
  input  [2:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_7,
  input  [3:0]  io_mod_proc_mod_3_mat_mod_table_mod_table_width,
  input  [3:0]  io_mod_proc_mod_3_mat_mod_table_mod_table_depth,
  input         io_mod_proc_mod_3_act_mod_en,
  input  [7:0]  io_mod_proc_mod_3_act_mod_addr,
  input  [63:0] io_mod_proc_mod_3_act_mod_data_0,
  input  [63:0] io_mod_proc_mod_3_act_mod_data_1,
  input         io_mod_xbar_mod_en,
  input  [1:0]  io_mod_xbar_mod_first_proc_id,
  input  [1:0]  io_mod_xbar_mod_last_proc_id,
  input  [1:0]  io_mod_xbar_mod_next_proc_id_0,
  input  [1:0]  io_mod_xbar_mod_next_proc_id_1,
  input  [1:0]  io_mod_xbar_mod_next_proc_id_2,
  input  [1:0]  io_mod_xbar_mod_next_proc_id_3,
  input  [2:0]  io_w_0_wcs,
  input         io_w_0_w_en,
  input  [7:0]  io_w_0_w_addr,
  input  [63:0] io_w_0_w_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  proc_0_clock; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_95; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 56:25]
  wire [1:0] proc_0_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_0_io_pipe_phv_in_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_0_io_pipe_phv_in_is_valid_processor; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_95; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_0_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 56:25]
  wire [1:0] proc_0_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_0_io_pipe_phv_out_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_0_io_mod_par_mod_en; // @[ipsa.scala 56:25]
  wire  proc_0_io_mod_par_mod_last_mau_id_mod; // @[ipsa.scala 56:25]
  wire [2:0] proc_0_io_mod_par_mod_last_mau_id; // @[ipsa.scala 56:25]
  wire [2:0] proc_0_io_mod_par_mod_cs; // @[ipsa.scala 56:25]
  wire  proc_0_io_mod_par_mod_module_mod_state_id_mod; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_mod_par_mod_module_mod_state_id; // @[ipsa.scala 56:25]
  wire  proc_0_io_mod_par_mod_module_mod_sram_w_cs; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_mod_par_mod_module_mod_sram_w_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_0_io_mod_par_mod_module_mod_sram_w_data; // @[ipsa.scala 56:25]
  wire  proc_0_io_mod_mat_mod_en; // @[ipsa.scala 56:25]
  wire  proc_0_io_mod_mat_mod_config_id; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_mod_mat_mod_key_mod_header_id; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_mod_mat_mod_key_mod_internal_offset; // @[ipsa.scala 56:25]
  wire [3:0] proc_0_io_mod_mat_mod_key_mod_key_length; // @[ipsa.scala 56:25]
  wire [3:0] proc_0_io_mod_mat_mod_table_mod_table_width; // @[ipsa.scala 56:25]
  wire [3:0] proc_0_io_mod_mat_mod_table_mod_table_depth; // @[ipsa.scala 56:25]
  wire  proc_0_io_mod_act_mod_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_mod_act_mod_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_0_io_mod_act_mod_data_0; // @[ipsa.scala 56:25]
  wire [63:0] proc_0_io_mod_act_mod_data_1; // @[ipsa.scala 56:25]
  wire  proc_0_io_mem_cluster_0_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_mem_cluster_0_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_0_io_mem_cluster_0_data; // @[ipsa.scala 56:25]
  wire  proc_0_io_mem_cluster_1_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_mem_cluster_1_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_0_io_mem_cluster_1_data; // @[ipsa.scala 56:25]
  wire  proc_0_io_mem_cluster_2_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_mem_cluster_2_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_0_io_mem_cluster_2_data; // @[ipsa.scala 56:25]
  wire  proc_0_io_mem_cluster_3_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_mem_cluster_3_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_0_io_mem_cluster_3_data; // @[ipsa.scala 56:25]
  wire  proc_0_io_mem_cluster_4_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_mem_cluster_4_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_0_io_mem_cluster_4_data; // @[ipsa.scala 56:25]
  wire  proc_0_io_mem_cluster_5_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_mem_cluster_5_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_0_io_mem_cluster_5_data; // @[ipsa.scala 56:25]
  wire  proc_0_io_mem_cluster_6_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_mem_cluster_6_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_0_io_mem_cluster_6_data; // @[ipsa.scala 56:25]
  wire  proc_0_io_mem_cluster_7_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_0_io_mem_cluster_7_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_0_io_mem_cluster_7_data; // @[ipsa.scala 56:25]
  wire  proc_1_clock; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_95; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 56:25]
  wire [1:0] proc_1_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_1_io_pipe_phv_in_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_1_io_pipe_phv_in_is_valid_processor; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_95; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_1_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 56:25]
  wire [1:0] proc_1_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_1_io_pipe_phv_out_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_1_io_mod_par_mod_en; // @[ipsa.scala 56:25]
  wire  proc_1_io_mod_par_mod_last_mau_id_mod; // @[ipsa.scala 56:25]
  wire [2:0] proc_1_io_mod_par_mod_last_mau_id; // @[ipsa.scala 56:25]
  wire [2:0] proc_1_io_mod_par_mod_cs; // @[ipsa.scala 56:25]
  wire  proc_1_io_mod_par_mod_module_mod_state_id_mod; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_mod_par_mod_module_mod_state_id; // @[ipsa.scala 56:25]
  wire  proc_1_io_mod_par_mod_module_mod_sram_w_cs; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_mod_par_mod_module_mod_sram_w_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_1_io_mod_par_mod_module_mod_sram_w_data; // @[ipsa.scala 56:25]
  wire  proc_1_io_mod_mat_mod_en; // @[ipsa.scala 56:25]
  wire  proc_1_io_mod_mat_mod_config_id; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_mod_mat_mod_key_mod_header_id; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_mod_mat_mod_key_mod_internal_offset; // @[ipsa.scala 56:25]
  wire [3:0] proc_1_io_mod_mat_mod_key_mod_key_length; // @[ipsa.scala 56:25]
  wire [3:0] proc_1_io_mod_mat_mod_table_mod_table_width; // @[ipsa.scala 56:25]
  wire [3:0] proc_1_io_mod_mat_mod_table_mod_table_depth; // @[ipsa.scala 56:25]
  wire  proc_1_io_mod_act_mod_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_mod_act_mod_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_1_io_mod_act_mod_data_0; // @[ipsa.scala 56:25]
  wire [63:0] proc_1_io_mod_act_mod_data_1; // @[ipsa.scala 56:25]
  wire  proc_1_io_mem_cluster_0_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_mem_cluster_0_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_1_io_mem_cluster_0_data; // @[ipsa.scala 56:25]
  wire  proc_1_io_mem_cluster_1_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_mem_cluster_1_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_1_io_mem_cluster_1_data; // @[ipsa.scala 56:25]
  wire  proc_1_io_mem_cluster_2_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_mem_cluster_2_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_1_io_mem_cluster_2_data; // @[ipsa.scala 56:25]
  wire  proc_1_io_mem_cluster_3_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_mem_cluster_3_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_1_io_mem_cluster_3_data; // @[ipsa.scala 56:25]
  wire  proc_1_io_mem_cluster_4_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_mem_cluster_4_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_1_io_mem_cluster_4_data; // @[ipsa.scala 56:25]
  wire  proc_1_io_mem_cluster_5_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_mem_cluster_5_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_1_io_mem_cluster_5_data; // @[ipsa.scala 56:25]
  wire  proc_1_io_mem_cluster_6_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_mem_cluster_6_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_1_io_mem_cluster_6_data; // @[ipsa.scala 56:25]
  wire  proc_1_io_mem_cluster_7_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_1_io_mem_cluster_7_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_1_io_mem_cluster_7_data; // @[ipsa.scala 56:25]
  wire  proc_2_clock; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_95; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 56:25]
  wire [1:0] proc_2_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_2_io_pipe_phv_in_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_2_io_pipe_phv_in_is_valid_processor; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_95; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_2_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 56:25]
  wire [1:0] proc_2_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_2_io_pipe_phv_out_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_2_io_mod_par_mod_en; // @[ipsa.scala 56:25]
  wire  proc_2_io_mod_par_mod_last_mau_id_mod; // @[ipsa.scala 56:25]
  wire [2:0] proc_2_io_mod_par_mod_last_mau_id; // @[ipsa.scala 56:25]
  wire [2:0] proc_2_io_mod_par_mod_cs; // @[ipsa.scala 56:25]
  wire  proc_2_io_mod_par_mod_module_mod_state_id_mod; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_mod_par_mod_module_mod_state_id; // @[ipsa.scala 56:25]
  wire  proc_2_io_mod_par_mod_module_mod_sram_w_cs; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_mod_par_mod_module_mod_sram_w_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_2_io_mod_par_mod_module_mod_sram_w_data; // @[ipsa.scala 56:25]
  wire  proc_2_io_mod_mat_mod_en; // @[ipsa.scala 56:25]
  wire  proc_2_io_mod_mat_mod_config_id; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_mod_mat_mod_key_mod_header_id; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_mod_mat_mod_key_mod_internal_offset; // @[ipsa.scala 56:25]
  wire [3:0] proc_2_io_mod_mat_mod_key_mod_key_length; // @[ipsa.scala 56:25]
  wire [3:0] proc_2_io_mod_mat_mod_table_mod_table_width; // @[ipsa.scala 56:25]
  wire [3:0] proc_2_io_mod_mat_mod_table_mod_table_depth; // @[ipsa.scala 56:25]
  wire  proc_2_io_mod_act_mod_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_mod_act_mod_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_2_io_mod_act_mod_data_0; // @[ipsa.scala 56:25]
  wire [63:0] proc_2_io_mod_act_mod_data_1; // @[ipsa.scala 56:25]
  wire  proc_2_io_mem_cluster_0_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_mem_cluster_0_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_2_io_mem_cluster_0_data; // @[ipsa.scala 56:25]
  wire  proc_2_io_mem_cluster_1_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_mem_cluster_1_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_2_io_mem_cluster_1_data; // @[ipsa.scala 56:25]
  wire  proc_2_io_mem_cluster_2_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_mem_cluster_2_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_2_io_mem_cluster_2_data; // @[ipsa.scala 56:25]
  wire  proc_2_io_mem_cluster_3_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_mem_cluster_3_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_2_io_mem_cluster_3_data; // @[ipsa.scala 56:25]
  wire  proc_2_io_mem_cluster_4_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_mem_cluster_4_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_2_io_mem_cluster_4_data; // @[ipsa.scala 56:25]
  wire  proc_2_io_mem_cluster_5_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_mem_cluster_5_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_2_io_mem_cluster_5_data; // @[ipsa.scala 56:25]
  wire  proc_2_io_mem_cluster_6_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_mem_cluster_6_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_2_io_mem_cluster_6_data; // @[ipsa.scala 56:25]
  wire  proc_2_io_mem_cluster_7_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_2_io_mem_cluster_7_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_2_io_mem_cluster_7_data; // @[ipsa.scala 56:25]
  wire  proc_3_clock; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_95; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 56:25]
  wire [1:0] proc_3_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_3_io_pipe_phv_in_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_3_io_pipe_phv_in_is_valid_processor; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_0; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_1; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_2; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_3; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_4; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_5; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_6; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_7; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_8; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_9; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_10; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_11; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_12; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_13; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_14; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_16; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_17; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_18; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_19; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_20; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_21; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_22; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_23; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_24; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_25; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_26; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_27; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_28; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_29; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_30; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_31; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_32; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_33; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_34; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_35; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_36; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_37; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_38; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_39; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_40; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_41; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_42; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_43; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_44; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_45; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_46; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_47; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_48; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_49; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_50; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_51; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_52; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_53; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_54; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_55; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_56; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_57; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_58; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_59; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_60; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_61; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_62; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_63; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_64; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_65; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_66; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_67; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_68; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_69; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_70; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_71; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_72; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_73; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_74; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_75; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_76; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_77; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_78; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_79; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_80; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_81; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_82; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_83; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_84; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_85; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_86; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_87; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_88; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_89; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_90; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_91; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_92; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_93; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_94; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_95; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_0; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_1; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_2; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_3; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_4; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_5; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_6; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_7; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_8; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_9; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_10; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_11; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_12; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_13; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_14; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_15; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 56:25]
  wire [15:0] proc_3_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 56:25]
  wire [1:0] proc_3_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 56:25]
  wire  proc_3_io_pipe_phv_out_next_config_id; // @[ipsa.scala 56:25]
  wire  proc_3_io_mod_par_mod_en; // @[ipsa.scala 56:25]
  wire  proc_3_io_mod_par_mod_last_mau_id_mod; // @[ipsa.scala 56:25]
  wire [2:0] proc_3_io_mod_par_mod_last_mau_id; // @[ipsa.scala 56:25]
  wire [2:0] proc_3_io_mod_par_mod_cs; // @[ipsa.scala 56:25]
  wire  proc_3_io_mod_par_mod_module_mod_state_id_mod; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_mod_par_mod_module_mod_state_id; // @[ipsa.scala 56:25]
  wire  proc_3_io_mod_par_mod_module_mod_sram_w_cs; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_mod_par_mod_module_mod_sram_w_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_3_io_mod_par_mod_module_mod_sram_w_data; // @[ipsa.scala 56:25]
  wire  proc_3_io_mod_mat_mod_en; // @[ipsa.scala 56:25]
  wire  proc_3_io_mod_mat_mod_config_id; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_mod_mat_mod_key_mod_header_id; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_mod_mat_mod_key_mod_internal_offset; // @[ipsa.scala 56:25]
  wire [3:0] proc_3_io_mod_mat_mod_key_mod_key_length; // @[ipsa.scala 56:25]
  wire [3:0] proc_3_io_mod_mat_mod_table_mod_table_width; // @[ipsa.scala 56:25]
  wire [3:0] proc_3_io_mod_mat_mod_table_mod_table_depth; // @[ipsa.scala 56:25]
  wire  proc_3_io_mod_act_mod_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_mod_act_mod_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_3_io_mod_act_mod_data_0; // @[ipsa.scala 56:25]
  wire [63:0] proc_3_io_mod_act_mod_data_1; // @[ipsa.scala 56:25]
  wire  proc_3_io_mem_cluster_0_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_mem_cluster_0_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_3_io_mem_cluster_0_data; // @[ipsa.scala 56:25]
  wire  proc_3_io_mem_cluster_1_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_mem_cluster_1_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_3_io_mem_cluster_1_data; // @[ipsa.scala 56:25]
  wire  proc_3_io_mem_cluster_2_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_mem_cluster_2_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_3_io_mem_cluster_2_data; // @[ipsa.scala 56:25]
  wire  proc_3_io_mem_cluster_3_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_mem_cluster_3_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_3_io_mem_cluster_3_data; // @[ipsa.scala 56:25]
  wire  proc_3_io_mem_cluster_4_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_mem_cluster_4_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_3_io_mem_cluster_4_data; // @[ipsa.scala 56:25]
  wire  proc_3_io_mem_cluster_5_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_mem_cluster_5_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_3_io_mem_cluster_5_data; // @[ipsa.scala 56:25]
  wire  proc_3_io_mem_cluster_6_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_mem_cluster_6_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_3_io_mem_cluster_6_data; // @[ipsa.scala 56:25]
  wire  proc_3_io_mem_cluster_7_en; // @[ipsa.scala 56:25]
  wire [7:0] proc_3_io_mem_cluster_7_addr; // @[ipsa.scala 56:25]
  wire [63:0] proc_3_io_mem_cluster_7_data; // @[ipsa.scala 56:25]
  wire  sram_cluster_0_clock; // @[ipsa.scala 62:25]
  wire [2:0] sram_cluster_0_io_w_wcs; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_w_w_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_w_w_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_w_w_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_0_cluster_0_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_0_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_0_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_0_cluster_1_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_1_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_1_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_0_cluster_2_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_2_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_2_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_0_cluster_3_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_3_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_3_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_0_cluster_4_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_4_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_4_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_0_cluster_5_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_5_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_5_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_0_cluster_6_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_6_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_6_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_0_cluster_7_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_7_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_7_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_1_cluster_0_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_0_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_0_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_1_cluster_1_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_1_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_1_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_1_cluster_2_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_2_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_2_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_1_cluster_3_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_3_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_3_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_1_cluster_4_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_4_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_4_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_1_cluster_5_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_5_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_5_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_1_cluster_6_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_6_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_6_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_1_cluster_7_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_7_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_7_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_2_cluster_0_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_0_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_0_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_2_cluster_1_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_1_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_1_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_2_cluster_2_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_2_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_2_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_2_cluster_3_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_3_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_3_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_2_cluster_4_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_4_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_4_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_2_cluster_5_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_5_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_5_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_2_cluster_6_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_6_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_6_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_2_cluster_7_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_7_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_7_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_3_cluster_0_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_0_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_0_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_3_cluster_1_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_1_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_1_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_3_cluster_2_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_2_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_2_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_3_cluster_3_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_3_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_3_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_3_cluster_4_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_4_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_4_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_3_cluster_5_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_5_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_5_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_3_cluster_6_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_6_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_6_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_io_r_3_cluster_7_en; // @[ipsa.scala 62:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_7_addr; // @[ipsa.scala 62:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_7_data; // @[ipsa.scala 62:25]
  wire  init_clock; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_0; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_1; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_2; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_3; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_4; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_5; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_6; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_7; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_8; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_9; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_10; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_11; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_12; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_13; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_14; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_15; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_16; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_17; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_18; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_19; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_20; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_21; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_22; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_23; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_24; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_25; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_26; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_27; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_28; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_29; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_30; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_31; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_32; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_33; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_34; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_35; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_36; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_37; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_38; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_39; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_40; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_41; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_42; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_43; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_44; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_45; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_46; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_47; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_48; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_49; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_50; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_51; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_52; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_53; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_54; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_55; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_56; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_57; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_58; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_59; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_60; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_61; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_62; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_63; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_64; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_65; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_66; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_67; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_68; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_69; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_70; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_71; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_72; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_73; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_74; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_75; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_76; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_77; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_78; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_79; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_80; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_81; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_82; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_83; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_84; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_85; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_86; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_87; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_88; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_89; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_90; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_91; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_92; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_93; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_94; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_data_95; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_in_header_0; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_in_header_1; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_in_header_2; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_in_header_3; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_in_header_4; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_in_header_5; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_in_header_6; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_in_header_7; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_in_header_8; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_in_header_9; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_in_header_10; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_in_header_11; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_in_header_12; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_in_header_13; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_in_header_14; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_in_header_15; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_0; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_1; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_2; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_3; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_4; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_5; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_6; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_7; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_8; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_9; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_10; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_11; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_12; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_13; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_14; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_15; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_16; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_17; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_18; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_19; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_20; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_21; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_22; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_23; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_24; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_25; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_26; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_27; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_28; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_29; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_30; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_31; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_32; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_33; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_34; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_35; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_36; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_37; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_38; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_39; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_40; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_41; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_42; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_43; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_44; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_45; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_46; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_47; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_48; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_49; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_50; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_51; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_52; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_53; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_54; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_55; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_56; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_57; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_58; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_59; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_60; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_61; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_62; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_63; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_64; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_65; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_66; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_67; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_68; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_69; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_70; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_71; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_72; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_73; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_74; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_75; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_76; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_77; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_78; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_79; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_80; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_81; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_82; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_83; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_84; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_85; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_86; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_87; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_88; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_89; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_90; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_91; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_92; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_93; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_94; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_data_95; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_out_header_0; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_out_header_1; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_out_header_2; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_out_header_3; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_out_header_4; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_out_header_5; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_out_header_6; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_out_header_7; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_out_header_8; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_out_header_9; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_out_header_10; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_out_header_11; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_out_header_12; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_out_header_13; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_out_header_14; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_out_header_15; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 74:22]
  wire [7:0] init_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 74:22]
  wire [15:0] init_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 74:22]
  wire [1:0] init_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 74:22]
  wire [1:0] init_io_first_proc_id; // @[ipsa.scala 74:22]
  wire  trans_0_clock; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_95; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 79:25]
  wire [1:0] trans_0_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_0_io_pipe_phv_in_next_config_id; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_95; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_0_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_0_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 79:25]
  wire [1:0] trans_0_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_0_io_pipe_phv_out_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_0_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 79:25]
  wire  trans_0_io_next_proc_exist; // @[ipsa.scala 79:25]
  wire [1:0] trans_0_io_next_proc_id; // @[ipsa.scala 79:25]
  wire  trans_1_clock; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_95; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 79:25]
  wire [1:0] trans_1_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_1_io_pipe_phv_in_next_config_id; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_95; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_1_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_1_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 79:25]
  wire [1:0] trans_1_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_1_io_pipe_phv_out_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_1_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 79:25]
  wire  trans_1_io_next_proc_exist; // @[ipsa.scala 79:25]
  wire [1:0] trans_1_io_next_proc_id; // @[ipsa.scala 79:25]
  wire  trans_2_clock; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_95; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 79:25]
  wire [1:0] trans_2_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_2_io_pipe_phv_in_next_config_id; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_95; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_2_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_2_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 79:25]
  wire [1:0] trans_2_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_2_io_pipe_phv_out_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_2_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 79:25]
  wire  trans_2_io_next_proc_exist; // @[ipsa.scala 79:25]
  wire [1:0] trans_2_io_next_proc_id; // @[ipsa.scala 79:25]
  wire  trans_3_clock; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_95; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 79:25]
  wire [1:0] trans_3_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_3_io_pipe_phv_in_next_config_id; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_0; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_1; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_2; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_3; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_4; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_5; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_6; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_7; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_8; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_9; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_10; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_11; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_12; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_13; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_14; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_16; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_17; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_18; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_19; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_20; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_21; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_22; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_23; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_24; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_25; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_26; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_27; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_28; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_29; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_30; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_31; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_32; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_33; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_34; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_35; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_36; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_37; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_38; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_39; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_40; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_41; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_42; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_43; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_44; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_45; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_46; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_47; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_48; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_49; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_50; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_51; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_52; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_53; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_54; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_55; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_56; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_57; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_58; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_59; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_60; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_61; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_62; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_63; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_64; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_65; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_66; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_67; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_68; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_69; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_70; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_71; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_72; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_73; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_74; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_75; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_76; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_77; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_78; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_79; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_80; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_81; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_82; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_83; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_84; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_85; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_86; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_87; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_88; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_89; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_90; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_91; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_92; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_93; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_94; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_95; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_0; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_1; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_2; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_3; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_4; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_5; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_6; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_7; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_8; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_9; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_10; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_11; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_12; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_13; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_14; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_15; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 79:25]
  wire [7:0] trans_3_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 79:25]
  wire [15:0] trans_3_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 79:25]
  wire [1:0] trans_3_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 79:25]
  wire  trans_3_io_pipe_phv_out_next_config_id; // @[ipsa.scala 79:25]
  wire  trans_3_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 79:25]
  wire  trans_3_io_next_proc_exist; // @[ipsa.scala 79:25]
  wire [1:0] trans_3_io_next_proc_id; // @[ipsa.scala 79:25]
  reg [1:0] first_proc_id; // @[ipsa.scala 43:28]
  reg [1:0] last_proc_id; // @[ipsa.scala 44:28]
  reg [1:0] next_proc_id_0; // @[ipsa.scala 45:28]
  reg [1:0] next_proc_id_1; // @[ipsa.scala 45:28]
  reg [1:0] next_proc_id_2; // @[ipsa.scala 45:28]
  reg [1:0] next_proc_id_3; // @[ipsa.scala 45:28]
  wire  _GEN_6 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_is_valid_processor : 2'h0 == first_proc_id; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 89:51]
  wire  _GEN_7 = 2'h0 == next_proc_id_0 & trans_0_io_pipe_phv_out_next_config_id; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [1:0] _GEN_8 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_next_processor_id :
    init_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_9 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_parse_transition_field :
    init_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_10 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_parse_current_offset :
    init_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_11 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_parse_current_state :
    init_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_12 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_0 : init_io_pipe_phv_out_header_0; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_13 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_1 : init_io_pipe_phv_out_header_1; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_14 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_2 : init_io_pipe_phv_out_header_2; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_15 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_3 : init_io_pipe_phv_out_header_3; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_16 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_4 : init_io_pipe_phv_out_header_4; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_17 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_5 : init_io_pipe_phv_out_header_5; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_18 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_6 : init_io_pipe_phv_out_header_6; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_19 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_7 : init_io_pipe_phv_out_header_7; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_20 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_8 : init_io_pipe_phv_out_header_8; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_21 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_9 : init_io_pipe_phv_out_header_9; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_22 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_10 : init_io_pipe_phv_out_header_10; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_23 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_11 : init_io_pipe_phv_out_header_11; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_24 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_12 : init_io_pipe_phv_out_header_12; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_25 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_13 : init_io_pipe_phv_out_header_13; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_26 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_14 : init_io_pipe_phv_out_header_14; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_27 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_15 : init_io_pipe_phv_out_header_15; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_28 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_0 : init_io_pipe_phv_out_data_0; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_29 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_1 : init_io_pipe_phv_out_data_1; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_30 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_2 : init_io_pipe_phv_out_data_2; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_31 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_3 : init_io_pipe_phv_out_data_3; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_32 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_4 : init_io_pipe_phv_out_data_4; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_33 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_5 : init_io_pipe_phv_out_data_5; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_34 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_6 : init_io_pipe_phv_out_data_6; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_35 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_7 : init_io_pipe_phv_out_data_7; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_36 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_8 : init_io_pipe_phv_out_data_8; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_37 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_9 : init_io_pipe_phv_out_data_9; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_38 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_10 : init_io_pipe_phv_out_data_10; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_39 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_11 : init_io_pipe_phv_out_data_11; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_40 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_12 : init_io_pipe_phv_out_data_12; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_41 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_13 : init_io_pipe_phv_out_data_13; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_42 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_14 : init_io_pipe_phv_out_data_14; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_43 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_15 : init_io_pipe_phv_out_data_15; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_44 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_16 : init_io_pipe_phv_out_data_16; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_45 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_17 : init_io_pipe_phv_out_data_17; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_46 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_18 : init_io_pipe_phv_out_data_18; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_47 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_19 : init_io_pipe_phv_out_data_19; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_48 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_20 : init_io_pipe_phv_out_data_20; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_49 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_21 : init_io_pipe_phv_out_data_21; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_50 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_22 : init_io_pipe_phv_out_data_22; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_51 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_23 : init_io_pipe_phv_out_data_23; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_52 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_24 : init_io_pipe_phv_out_data_24; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_53 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_25 : init_io_pipe_phv_out_data_25; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_54 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_26 : init_io_pipe_phv_out_data_26; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_55 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_27 : init_io_pipe_phv_out_data_27; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_56 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_28 : init_io_pipe_phv_out_data_28; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_57 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_29 : init_io_pipe_phv_out_data_29; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_58 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_30 : init_io_pipe_phv_out_data_30; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_59 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_31 : init_io_pipe_phv_out_data_31; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_60 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_32 : init_io_pipe_phv_out_data_32; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_61 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_33 : init_io_pipe_phv_out_data_33; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_62 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_34 : init_io_pipe_phv_out_data_34; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_63 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_35 : init_io_pipe_phv_out_data_35; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_64 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_36 : init_io_pipe_phv_out_data_36; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_65 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_37 : init_io_pipe_phv_out_data_37; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_66 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_38 : init_io_pipe_phv_out_data_38; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_67 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_39 : init_io_pipe_phv_out_data_39; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_68 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_40 : init_io_pipe_phv_out_data_40; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_69 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_41 : init_io_pipe_phv_out_data_41; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_70 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_42 : init_io_pipe_phv_out_data_42; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_71 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_43 : init_io_pipe_phv_out_data_43; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_72 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_44 : init_io_pipe_phv_out_data_44; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_73 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_45 : init_io_pipe_phv_out_data_45; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_74 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_46 : init_io_pipe_phv_out_data_46; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_75 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_47 : init_io_pipe_phv_out_data_47; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_76 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_48 : init_io_pipe_phv_out_data_48; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_77 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_49 : init_io_pipe_phv_out_data_49; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_78 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_50 : init_io_pipe_phv_out_data_50; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_79 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_51 : init_io_pipe_phv_out_data_51; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_80 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_52 : init_io_pipe_phv_out_data_52; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_81 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_53 : init_io_pipe_phv_out_data_53; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_82 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_54 : init_io_pipe_phv_out_data_54; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_83 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_55 : init_io_pipe_phv_out_data_55; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_84 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_56 : init_io_pipe_phv_out_data_56; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_85 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_57 : init_io_pipe_phv_out_data_57; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_86 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_58 : init_io_pipe_phv_out_data_58; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_87 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_59 : init_io_pipe_phv_out_data_59; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_88 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_60 : init_io_pipe_phv_out_data_60; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_89 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_61 : init_io_pipe_phv_out_data_61; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_90 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_62 : init_io_pipe_phv_out_data_62; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_91 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_63 : init_io_pipe_phv_out_data_63; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_92 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_64 : init_io_pipe_phv_out_data_64; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_93 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_65 : init_io_pipe_phv_out_data_65; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_94 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_66 : init_io_pipe_phv_out_data_66; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_95 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_67 : init_io_pipe_phv_out_data_67; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_96 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_68 : init_io_pipe_phv_out_data_68; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_97 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_69 : init_io_pipe_phv_out_data_69; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_98 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_70 : init_io_pipe_phv_out_data_70; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_99 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_71 : init_io_pipe_phv_out_data_71; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_100 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_72 : init_io_pipe_phv_out_data_72; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_101 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_73 : init_io_pipe_phv_out_data_73; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_102 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_74 : init_io_pipe_phv_out_data_74; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_103 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_75 : init_io_pipe_phv_out_data_75; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_104 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_76 : init_io_pipe_phv_out_data_76; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_105 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_77 : init_io_pipe_phv_out_data_77; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_106 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_78 : init_io_pipe_phv_out_data_78; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_107 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_79 : init_io_pipe_phv_out_data_79; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_108 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_80 : init_io_pipe_phv_out_data_80; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_109 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_81 : init_io_pipe_phv_out_data_81; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_110 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_82 : init_io_pipe_phv_out_data_82; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_111 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_83 : init_io_pipe_phv_out_data_83; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_112 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_84 : init_io_pipe_phv_out_data_84; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_113 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_85 : init_io_pipe_phv_out_data_85; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_114 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_86 : init_io_pipe_phv_out_data_86; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_115 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_87 : init_io_pipe_phv_out_data_87; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_116 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_88 : init_io_pipe_phv_out_data_88; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_117 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_89 : init_io_pipe_phv_out_data_89; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_118 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_90 : init_io_pipe_phv_out_data_90; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_119 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_91 : init_io_pipe_phv_out_data_91; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_120 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_92 : init_io_pipe_phv_out_data_92; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_121 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_93 : init_io_pipe_phv_out_data_93; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_122 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_94 : init_io_pipe_phv_out_data_94; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_123 = 2'h0 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_95 : init_io_pipe_phv_out_data_95; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire  _GEN_124 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_is_valid_processor : 2'h1 == first_proc_id; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 89:51]
  wire  _GEN_125 = 2'h1 == next_proc_id_0 & trans_0_io_pipe_phv_out_next_config_id; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [1:0] _GEN_126 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_next_processor_id :
    init_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_127 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_parse_transition_field :
    init_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_128 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_parse_current_offset :
    init_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_129 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_parse_current_state :
    init_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_130 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_0 : init_io_pipe_phv_out_header_0; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_131 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_1 : init_io_pipe_phv_out_header_1; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_132 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_2 : init_io_pipe_phv_out_header_2; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_133 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_3 : init_io_pipe_phv_out_header_3; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_134 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_4 : init_io_pipe_phv_out_header_4; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_135 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_5 : init_io_pipe_phv_out_header_5; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_136 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_6 : init_io_pipe_phv_out_header_6; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_137 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_7 : init_io_pipe_phv_out_header_7; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_138 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_8 : init_io_pipe_phv_out_header_8; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_139 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_9 : init_io_pipe_phv_out_header_9; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_140 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_10 : init_io_pipe_phv_out_header_10; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_141 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_11 : init_io_pipe_phv_out_header_11; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_142 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_12 : init_io_pipe_phv_out_header_12; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_143 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_13 : init_io_pipe_phv_out_header_13; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_144 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_14 : init_io_pipe_phv_out_header_14; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_145 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_15 : init_io_pipe_phv_out_header_15; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_146 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_0 : init_io_pipe_phv_out_data_0; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_147 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_1 : init_io_pipe_phv_out_data_1; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_148 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_2 : init_io_pipe_phv_out_data_2; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_149 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_3 : init_io_pipe_phv_out_data_3; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_150 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_4 : init_io_pipe_phv_out_data_4; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_151 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_5 : init_io_pipe_phv_out_data_5; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_152 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_6 : init_io_pipe_phv_out_data_6; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_153 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_7 : init_io_pipe_phv_out_data_7; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_154 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_8 : init_io_pipe_phv_out_data_8; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_155 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_9 : init_io_pipe_phv_out_data_9; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_156 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_10 : init_io_pipe_phv_out_data_10; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_157 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_11 : init_io_pipe_phv_out_data_11; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_158 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_12 : init_io_pipe_phv_out_data_12; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_159 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_13 : init_io_pipe_phv_out_data_13; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_160 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_14 : init_io_pipe_phv_out_data_14; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_161 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_15 : init_io_pipe_phv_out_data_15; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_162 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_16 : init_io_pipe_phv_out_data_16; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_163 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_17 : init_io_pipe_phv_out_data_17; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_164 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_18 : init_io_pipe_phv_out_data_18; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_165 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_19 : init_io_pipe_phv_out_data_19; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_166 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_20 : init_io_pipe_phv_out_data_20; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_167 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_21 : init_io_pipe_phv_out_data_21; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_168 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_22 : init_io_pipe_phv_out_data_22; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_169 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_23 : init_io_pipe_phv_out_data_23; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_170 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_24 : init_io_pipe_phv_out_data_24; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_171 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_25 : init_io_pipe_phv_out_data_25; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_172 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_26 : init_io_pipe_phv_out_data_26; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_173 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_27 : init_io_pipe_phv_out_data_27; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_174 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_28 : init_io_pipe_phv_out_data_28; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_175 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_29 : init_io_pipe_phv_out_data_29; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_176 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_30 : init_io_pipe_phv_out_data_30; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_177 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_31 : init_io_pipe_phv_out_data_31; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_178 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_32 : init_io_pipe_phv_out_data_32; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_179 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_33 : init_io_pipe_phv_out_data_33; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_180 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_34 : init_io_pipe_phv_out_data_34; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_181 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_35 : init_io_pipe_phv_out_data_35; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_182 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_36 : init_io_pipe_phv_out_data_36; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_183 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_37 : init_io_pipe_phv_out_data_37; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_184 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_38 : init_io_pipe_phv_out_data_38; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_185 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_39 : init_io_pipe_phv_out_data_39; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_186 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_40 : init_io_pipe_phv_out_data_40; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_187 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_41 : init_io_pipe_phv_out_data_41; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_188 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_42 : init_io_pipe_phv_out_data_42; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_189 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_43 : init_io_pipe_phv_out_data_43; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_190 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_44 : init_io_pipe_phv_out_data_44; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_191 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_45 : init_io_pipe_phv_out_data_45; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_192 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_46 : init_io_pipe_phv_out_data_46; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_193 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_47 : init_io_pipe_phv_out_data_47; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_194 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_48 : init_io_pipe_phv_out_data_48; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_195 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_49 : init_io_pipe_phv_out_data_49; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_196 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_50 : init_io_pipe_phv_out_data_50; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_197 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_51 : init_io_pipe_phv_out_data_51; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_198 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_52 : init_io_pipe_phv_out_data_52; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_199 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_53 : init_io_pipe_phv_out_data_53; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_200 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_54 : init_io_pipe_phv_out_data_54; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_201 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_55 : init_io_pipe_phv_out_data_55; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_202 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_56 : init_io_pipe_phv_out_data_56; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_203 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_57 : init_io_pipe_phv_out_data_57; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_204 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_58 : init_io_pipe_phv_out_data_58; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_205 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_59 : init_io_pipe_phv_out_data_59; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_206 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_60 : init_io_pipe_phv_out_data_60; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_207 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_61 : init_io_pipe_phv_out_data_61; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_208 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_62 : init_io_pipe_phv_out_data_62; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_209 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_63 : init_io_pipe_phv_out_data_63; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_210 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_64 : init_io_pipe_phv_out_data_64; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_211 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_65 : init_io_pipe_phv_out_data_65; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_212 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_66 : init_io_pipe_phv_out_data_66; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_213 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_67 : init_io_pipe_phv_out_data_67; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_214 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_68 : init_io_pipe_phv_out_data_68; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_215 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_69 : init_io_pipe_phv_out_data_69; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_216 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_70 : init_io_pipe_phv_out_data_70; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_217 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_71 : init_io_pipe_phv_out_data_71; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_218 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_72 : init_io_pipe_phv_out_data_72; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_219 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_73 : init_io_pipe_phv_out_data_73; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_220 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_74 : init_io_pipe_phv_out_data_74; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_221 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_75 : init_io_pipe_phv_out_data_75; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_222 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_76 : init_io_pipe_phv_out_data_76; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_223 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_77 : init_io_pipe_phv_out_data_77; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_224 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_78 : init_io_pipe_phv_out_data_78; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_225 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_79 : init_io_pipe_phv_out_data_79; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_226 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_80 : init_io_pipe_phv_out_data_80; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_227 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_81 : init_io_pipe_phv_out_data_81; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_228 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_82 : init_io_pipe_phv_out_data_82; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_229 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_83 : init_io_pipe_phv_out_data_83; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_230 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_84 : init_io_pipe_phv_out_data_84; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_231 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_85 : init_io_pipe_phv_out_data_85; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_232 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_86 : init_io_pipe_phv_out_data_86; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_233 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_87 : init_io_pipe_phv_out_data_87; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_234 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_88 : init_io_pipe_phv_out_data_88; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_235 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_89 : init_io_pipe_phv_out_data_89; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_236 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_90 : init_io_pipe_phv_out_data_90; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_237 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_91 : init_io_pipe_phv_out_data_91; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_238 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_92 : init_io_pipe_phv_out_data_92; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_239 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_93 : init_io_pipe_phv_out_data_93; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_240 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_94 : init_io_pipe_phv_out_data_94; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_241 = 2'h1 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_95 : init_io_pipe_phv_out_data_95; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire  _GEN_242 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_is_valid_processor : 2'h2 == first_proc_id; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 89:51]
  wire  _GEN_243 = 2'h2 == next_proc_id_0 & trans_0_io_pipe_phv_out_next_config_id; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [1:0] _GEN_244 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_next_processor_id :
    init_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_245 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_parse_transition_field :
    init_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_246 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_parse_current_offset :
    init_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_247 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_parse_current_state :
    init_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_248 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_0 : init_io_pipe_phv_out_header_0; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_249 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_1 : init_io_pipe_phv_out_header_1; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_250 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_2 : init_io_pipe_phv_out_header_2; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_251 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_3 : init_io_pipe_phv_out_header_3; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_252 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_4 : init_io_pipe_phv_out_header_4; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_253 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_5 : init_io_pipe_phv_out_header_5; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_254 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_6 : init_io_pipe_phv_out_header_6; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_255 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_7 : init_io_pipe_phv_out_header_7; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_256 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_8 : init_io_pipe_phv_out_header_8; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_257 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_9 : init_io_pipe_phv_out_header_9; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_258 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_10 : init_io_pipe_phv_out_header_10; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_259 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_11 : init_io_pipe_phv_out_header_11; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_260 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_12 : init_io_pipe_phv_out_header_12; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_261 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_13 : init_io_pipe_phv_out_header_13; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_262 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_14 : init_io_pipe_phv_out_header_14; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_263 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_15 : init_io_pipe_phv_out_header_15; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_264 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_0 : init_io_pipe_phv_out_data_0; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_265 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_1 : init_io_pipe_phv_out_data_1; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_266 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_2 : init_io_pipe_phv_out_data_2; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_267 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_3 : init_io_pipe_phv_out_data_3; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_268 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_4 : init_io_pipe_phv_out_data_4; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_269 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_5 : init_io_pipe_phv_out_data_5; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_270 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_6 : init_io_pipe_phv_out_data_6; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_271 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_7 : init_io_pipe_phv_out_data_7; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_272 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_8 : init_io_pipe_phv_out_data_8; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_273 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_9 : init_io_pipe_phv_out_data_9; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_274 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_10 : init_io_pipe_phv_out_data_10; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_275 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_11 : init_io_pipe_phv_out_data_11; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_276 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_12 : init_io_pipe_phv_out_data_12; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_277 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_13 : init_io_pipe_phv_out_data_13; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_278 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_14 : init_io_pipe_phv_out_data_14; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_279 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_15 : init_io_pipe_phv_out_data_15; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_280 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_16 : init_io_pipe_phv_out_data_16; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_281 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_17 : init_io_pipe_phv_out_data_17; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_282 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_18 : init_io_pipe_phv_out_data_18; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_283 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_19 : init_io_pipe_phv_out_data_19; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_284 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_20 : init_io_pipe_phv_out_data_20; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_285 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_21 : init_io_pipe_phv_out_data_21; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_286 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_22 : init_io_pipe_phv_out_data_22; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_287 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_23 : init_io_pipe_phv_out_data_23; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_288 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_24 : init_io_pipe_phv_out_data_24; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_289 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_25 : init_io_pipe_phv_out_data_25; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_290 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_26 : init_io_pipe_phv_out_data_26; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_291 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_27 : init_io_pipe_phv_out_data_27; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_292 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_28 : init_io_pipe_phv_out_data_28; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_293 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_29 : init_io_pipe_phv_out_data_29; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_294 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_30 : init_io_pipe_phv_out_data_30; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_295 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_31 : init_io_pipe_phv_out_data_31; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_296 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_32 : init_io_pipe_phv_out_data_32; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_297 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_33 : init_io_pipe_phv_out_data_33; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_298 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_34 : init_io_pipe_phv_out_data_34; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_299 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_35 : init_io_pipe_phv_out_data_35; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_300 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_36 : init_io_pipe_phv_out_data_36; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_301 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_37 : init_io_pipe_phv_out_data_37; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_302 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_38 : init_io_pipe_phv_out_data_38; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_303 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_39 : init_io_pipe_phv_out_data_39; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_304 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_40 : init_io_pipe_phv_out_data_40; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_305 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_41 : init_io_pipe_phv_out_data_41; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_306 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_42 : init_io_pipe_phv_out_data_42; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_307 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_43 : init_io_pipe_phv_out_data_43; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_308 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_44 : init_io_pipe_phv_out_data_44; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_309 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_45 : init_io_pipe_phv_out_data_45; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_310 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_46 : init_io_pipe_phv_out_data_46; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_311 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_47 : init_io_pipe_phv_out_data_47; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_312 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_48 : init_io_pipe_phv_out_data_48; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_313 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_49 : init_io_pipe_phv_out_data_49; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_314 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_50 : init_io_pipe_phv_out_data_50; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_315 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_51 : init_io_pipe_phv_out_data_51; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_316 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_52 : init_io_pipe_phv_out_data_52; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_317 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_53 : init_io_pipe_phv_out_data_53; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_318 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_54 : init_io_pipe_phv_out_data_54; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_319 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_55 : init_io_pipe_phv_out_data_55; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_320 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_56 : init_io_pipe_phv_out_data_56; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_321 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_57 : init_io_pipe_phv_out_data_57; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_322 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_58 : init_io_pipe_phv_out_data_58; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_323 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_59 : init_io_pipe_phv_out_data_59; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_324 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_60 : init_io_pipe_phv_out_data_60; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_325 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_61 : init_io_pipe_phv_out_data_61; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_326 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_62 : init_io_pipe_phv_out_data_62; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_327 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_63 : init_io_pipe_phv_out_data_63; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_328 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_64 : init_io_pipe_phv_out_data_64; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_329 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_65 : init_io_pipe_phv_out_data_65; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_330 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_66 : init_io_pipe_phv_out_data_66; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_331 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_67 : init_io_pipe_phv_out_data_67; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_332 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_68 : init_io_pipe_phv_out_data_68; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_333 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_69 : init_io_pipe_phv_out_data_69; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_334 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_70 : init_io_pipe_phv_out_data_70; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_335 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_71 : init_io_pipe_phv_out_data_71; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_336 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_72 : init_io_pipe_phv_out_data_72; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_337 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_73 : init_io_pipe_phv_out_data_73; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_338 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_74 : init_io_pipe_phv_out_data_74; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_339 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_75 : init_io_pipe_phv_out_data_75; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_340 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_76 : init_io_pipe_phv_out_data_76; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_341 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_77 : init_io_pipe_phv_out_data_77; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_342 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_78 : init_io_pipe_phv_out_data_78; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_343 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_79 : init_io_pipe_phv_out_data_79; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_344 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_80 : init_io_pipe_phv_out_data_80; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_345 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_81 : init_io_pipe_phv_out_data_81; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_346 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_82 : init_io_pipe_phv_out_data_82; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_347 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_83 : init_io_pipe_phv_out_data_83; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_348 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_84 : init_io_pipe_phv_out_data_84; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_349 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_85 : init_io_pipe_phv_out_data_85; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_350 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_86 : init_io_pipe_phv_out_data_86; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_351 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_87 : init_io_pipe_phv_out_data_87; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_352 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_88 : init_io_pipe_phv_out_data_88; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_353 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_89 : init_io_pipe_phv_out_data_89; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_354 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_90 : init_io_pipe_phv_out_data_90; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_355 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_91 : init_io_pipe_phv_out_data_91; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_356 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_92 : init_io_pipe_phv_out_data_92; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_357 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_93 : init_io_pipe_phv_out_data_93; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_358 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_94 : init_io_pipe_phv_out_data_94; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_359 = 2'h2 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_95 : init_io_pipe_phv_out_data_95; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire  _GEN_360 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_is_valid_processor : 2'h3 == first_proc_id; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 89:51]
  wire  _GEN_361 = 2'h3 == next_proc_id_0 & trans_0_io_pipe_phv_out_next_config_id; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [1:0] _GEN_362 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_next_processor_id :
    init_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_363 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_parse_transition_field :
    init_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_364 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_parse_current_offset :
    init_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_365 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_parse_current_state :
    init_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_366 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_0 : init_io_pipe_phv_out_header_0; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_367 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_1 : init_io_pipe_phv_out_header_1; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_368 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_2 : init_io_pipe_phv_out_header_2; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_369 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_3 : init_io_pipe_phv_out_header_3; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_370 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_4 : init_io_pipe_phv_out_header_4; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_371 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_5 : init_io_pipe_phv_out_header_5; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_372 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_6 : init_io_pipe_phv_out_header_6; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_373 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_7 : init_io_pipe_phv_out_header_7; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_374 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_8 : init_io_pipe_phv_out_header_8; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_375 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_9 : init_io_pipe_phv_out_header_9; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_376 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_10 : init_io_pipe_phv_out_header_10; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_377 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_11 : init_io_pipe_phv_out_header_11; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_378 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_12 : init_io_pipe_phv_out_header_12; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_379 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_13 : init_io_pipe_phv_out_header_13; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_380 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_14 : init_io_pipe_phv_out_header_14; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [15:0] _GEN_381 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_header_15 : init_io_pipe_phv_out_header_15; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_382 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_0 : init_io_pipe_phv_out_data_0; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_383 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_1 : init_io_pipe_phv_out_data_1; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_384 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_2 : init_io_pipe_phv_out_data_2; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_385 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_3 : init_io_pipe_phv_out_data_3; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_386 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_4 : init_io_pipe_phv_out_data_4; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_387 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_5 : init_io_pipe_phv_out_data_5; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_388 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_6 : init_io_pipe_phv_out_data_6; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_389 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_7 : init_io_pipe_phv_out_data_7; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_390 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_8 : init_io_pipe_phv_out_data_8; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_391 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_9 : init_io_pipe_phv_out_data_9; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_392 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_10 : init_io_pipe_phv_out_data_10; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_393 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_11 : init_io_pipe_phv_out_data_11; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_394 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_12 : init_io_pipe_phv_out_data_12; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_395 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_13 : init_io_pipe_phv_out_data_13; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_396 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_14 : init_io_pipe_phv_out_data_14; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_397 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_15 : init_io_pipe_phv_out_data_15; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_398 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_16 : init_io_pipe_phv_out_data_16; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_399 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_17 : init_io_pipe_phv_out_data_17; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_400 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_18 : init_io_pipe_phv_out_data_18; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_401 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_19 : init_io_pipe_phv_out_data_19; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_402 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_20 : init_io_pipe_phv_out_data_20; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_403 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_21 : init_io_pipe_phv_out_data_21; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_404 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_22 : init_io_pipe_phv_out_data_22; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_405 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_23 : init_io_pipe_phv_out_data_23; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_406 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_24 : init_io_pipe_phv_out_data_24; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_407 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_25 : init_io_pipe_phv_out_data_25; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_408 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_26 : init_io_pipe_phv_out_data_26; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_409 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_27 : init_io_pipe_phv_out_data_27; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_410 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_28 : init_io_pipe_phv_out_data_28; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_411 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_29 : init_io_pipe_phv_out_data_29; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_412 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_30 : init_io_pipe_phv_out_data_30; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_413 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_31 : init_io_pipe_phv_out_data_31; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_414 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_32 : init_io_pipe_phv_out_data_32; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_415 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_33 : init_io_pipe_phv_out_data_33; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_416 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_34 : init_io_pipe_phv_out_data_34; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_417 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_35 : init_io_pipe_phv_out_data_35; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_418 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_36 : init_io_pipe_phv_out_data_36; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_419 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_37 : init_io_pipe_phv_out_data_37; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_420 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_38 : init_io_pipe_phv_out_data_38; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_421 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_39 : init_io_pipe_phv_out_data_39; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_422 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_40 : init_io_pipe_phv_out_data_40; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_423 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_41 : init_io_pipe_phv_out_data_41; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_424 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_42 : init_io_pipe_phv_out_data_42; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_425 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_43 : init_io_pipe_phv_out_data_43; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_426 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_44 : init_io_pipe_phv_out_data_44; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_427 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_45 : init_io_pipe_phv_out_data_45; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_428 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_46 : init_io_pipe_phv_out_data_46; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_429 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_47 : init_io_pipe_phv_out_data_47; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_430 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_48 : init_io_pipe_phv_out_data_48; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_431 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_49 : init_io_pipe_phv_out_data_49; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_432 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_50 : init_io_pipe_phv_out_data_50; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_433 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_51 : init_io_pipe_phv_out_data_51; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_434 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_52 : init_io_pipe_phv_out_data_52; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_435 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_53 : init_io_pipe_phv_out_data_53; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_436 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_54 : init_io_pipe_phv_out_data_54; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_437 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_55 : init_io_pipe_phv_out_data_55; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_438 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_56 : init_io_pipe_phv_out_data_56; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_439 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_57 : init_io_pipe_phv_out_data_57; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_440 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_58 : init_io_pipe_phv_out_data_58; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_441 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_59 : init_io_pipe_phv_out_data_59; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_442 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_60 : init_io_pipe_phv_out_data_60; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_443 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_61 : init_io_pipe_phv_out_data_61; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_444 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_62 : init_io_pipe_phv_out_data_62; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_445 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_63 : init_io_pipe_phv_out_data_63; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_446 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_64 : init_io_pipe_phv_out_data_64; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_447 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_65 : init_io_pipe_phv_out_data_65; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_448 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_66 : init_io_pipe_phv_out_data_66; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_449 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_67 : init_io_pipe_phv_out_data_67; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_450 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_68 : init_io_pipe_phv_out_data_68; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_451 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_69 : init_io_pipe_phv_out_data_69; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_452 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_70 : init_io_pipe_phv_out_data_70; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_453 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_71 : init_io_pipe_phv_out_data_71; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_454 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_72 : init_io_pipe_phv_out_data_72; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_455 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_73 : init_io_pipe_phv_out_data_73; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_456 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_74 : init_io_pipe_phv_out_data_74; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_457 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_75 : init_io_pipe_phv_out_data_75; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_458 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_76 : init_io_pipe_phv_out_data_76; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_459 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_77 : init_io_pipe_phv_out_data_77; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_460 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_78 : init_io_pipe_phv_out_data_78; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_461 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_79 : init_io_pipe_phv_out_data_79; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_462 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_80 : init_io_pipe_phv_out_data_80; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_463 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_81 : init_io_pipe_phv_out_data_81; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_464 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_82 : init_io_pipe_phv_out_data_82; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_465 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_83 : init_io_pipe_phv_out_data_83; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_466 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_84 : init_io_pipe_phv_out_data_84; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_467 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_85 : init_io_pipe_phv_out_data_85; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_468 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_86 : init_io_pipe_phv_out_data_86; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_469 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_87 : init_io_pipe_phv_out_data_87; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_470 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_88 : init_io_pipe_phv_out_data_88; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_471 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_89 : init_io_pipe_phv_out_data_89; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_472 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_90 : init_io_pipe_phv_out_data_90; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_473 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_91 : init_io_pipe_phv_out_data_91; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_474 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_92 : init_io_pipe_phv_out_data_92; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_475 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_93 : init_io_pipe_phv_out_data_93; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_476 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_94 : init_io_pipe_phv_out_data_94; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire [7:0] _GEN_477 = 2'h3 == next_proc_id_0 ? trans_0_io_pipe_phv_out_data_95 : init_io_pipe_phv_out_data_95; // @[ipsa.scala 96:76 ipsa.scala 97:44 ipsa.scala 88:32]
  wire  _GEN_478 = 2'h0 != last_proc_id ? _GEN_6 : 2'h0 == first_proc_id; // @[ipsa.scala 94:65 ipsa.scala 89:51]
  wire  _GEN_479 = 2'h0 != last_proc_id & _GEN_7; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [1:0] _GEN_480 = 2'h0 != last_proc_id ? _GEN_8 : init_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_481 = 2'h0 != last_proc_id ? _GEN_9 : init_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_482 = 2'h0 != last_proc_id ? _GEN_10 : init_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_483 = 2'h0 != last_proc_id ? _GEN_11 : init_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_484 = 2'h0 != last_proc_id ? _GEN_12 : init_io_pipe_phv_out_header_0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_485 = 2'h0 != last_proc_id ? _GEN_13 : init_io_pipe_phv_out_header_1; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_486 = 2'h0 != last_proc_id ? _GEN_14 : init_io_pipe_phv_out_header_2; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_487 = 2'h0 != last_proc_id ? _GEN_15 : init_io_pipe_phv_out_header_3; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_488 = 2'h0 != last_proc_id ? _GEN_16 : init_io_pipe_phv_out_header_4; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_489 = 2'h0 != last_proc_id ? _GEN_17 : init_io_pipe_phv_out_header_5; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_490 = 2'h0 != last_proc_id ? _GEN_18 : init_io_pipe_phv_out_header_6; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_491 = 2'h0 != last_proc_id ? _GEN_19 : init_io_pipe_phv_out_header_7; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_492 = 2'h0 != last_proc_id ? _GEN_20 : init_io_pipe_phv_out_header_8; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_493 = 2'h0 != last_proc_id ? _GEN_21 : init_io_pipe_phv_out_header_9; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_494 = 2'h0 != last_proc_id ? _GEN_22 : init_io_pipe_phv_out_header_10; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_495 = 2'h0 != last_proc_id ? _GEN_23 : init_io_pipe_phv_out_header_11; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_496 = 2'h0 != last_proc_id ? _GEN_24 : init_io_pipe_phv_out_header_12; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_497 = 2'h0 != last_proc_id ? _GEN_25 : init_io_pipe_phv_out_header_13; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_498 = 2'h0 != last_proc_id ? _GEN_26 : init_io_pipe_phv_out_header_14; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_499 = 2'h0 != last_proc_id ? _GEN_27 : init_io_pipe_phv_out_header_15; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_500 = 2'h0 != last_proc_id ? _GEN_28 : init_io_pipe_phv_out_data_0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_501 = 2'h0 != last_proc_id ? _GEN_29 : init_io_pipe_phv_out_data_1; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_502 = 2'h0 != last_proc_id ? _GEN_30 : init_io_pipe_phv_out_data_2; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_503 = 2'h0 != last_proc_id ? _GEN_31 : init_io_pipe_phv_out_data_3; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_504 = 2'h0 != last_proc_id ? _GEN_32 : init_io_pipe_phv_out_data_4; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_505 = 2'h0 != last_proc_id ? _GEN_33 : init_io_pipe_phv_out_data_5; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_506 = 2'h0 != last_proc_id ? _GEN_34 : init_io_pipe_phv_out_data_6; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_507 = 2'h0 != last_proc_id ? _GEN_35 : init_io_pipe_phv_out_data_7; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_508 = 2'h0 != last_proc_id ? _GEN_36 : init_io_pipe_phv_out_data_8; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_509 = 2'h0 != last_proc_id ? _GEN_37 : init_io_pipe_phv_out_data_9; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_510 = 2'h0 != last_proc_id ? _GEN_38 : init_io_pipe_phv_out_data_10; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_511 = 2'h0 != last_proc_id ? _GEN_39 : init_io_pipe_phv_out_data_11; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_512 = 2'h0 != last_proc_id ? _GEN_40 : init_io_pipe_phv_out_data_12; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_513 = 2'h0 != last_proc_id ? _GEN_41 : init_io_pipe_phv_out_data_13; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_514 = 2'h0 != last_proc_id ? _GEN_42 : init_io_pipe_phv_out_data_14; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_515 = 2'h0 != last_proc_id ? _GEN_43 : init_io_pipe_phv_out_data_15; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_516 = 2'h0 != last_proc_id ? _GEN_44 : init_io_pipe_phv_out_data_16; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_517 = 2'h0 != last_proc_id ? _GEN_45 : init_io_pipe_phv_out_data_17; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_518 = 2'h0 != last_proc_id ? _GEN_46 : init_io_pipe_phv_out_data_18; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_519 = 2'h0 != last_proc_id ? _GEN_47 : init_io_pipe_phv_out_data_19; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_520 = 2'h0 != last_proc_id ? _GEN_48 : init_io_pipe_phv_out_data_20; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_521 = 2'h0 != last_proc_id ? _GEN_49 : init_io_pipe_phv_out_data_21; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_522 = 2'h0 != last_proc_id ? _GEN_50 : init_io_pipe_phv_out_data_22; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_523 = 2'h0 != last_proc_id ? _GEN_51 : init_io_pipe_phv_out_data_23; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_524 = 2'h0 != last_proc_id ? _GEN_52 : init_io_pipe_phv_out_data_24; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_525 = 2'h0 != last_proc_id ? _GEN_53 : init_io_pipe_phv_out_data_25; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_526 = 2'h0 != last_proc_id ? _GEN_54 : init_io_pipe_phv_out_data_26; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_527 = 2'h0 != last_proc_id ? _GEN_55 : init_io_pipe_phv_out_data_27; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_528 = 2'h0 != last_proc_id ? _GEN_56 : init_io_pipe_phv_out_data_28; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_529 = 2'h0 != last_proc_id ? _GEN_57 : init_io_pipe_phv_out_data_29; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_530 = 2'h0 != last_proc_id ? _GEN_58 : init_io_pipe_phv_out_data_30; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_531 = 2'h0 != last_proc_id ? _GEN_59 : init_io_pipe_phv_out_data_31; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_532 = 2'h0 != last_proc_id ? _GEN_60 : init_io_pipe_phv_out_data_32; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_533 = 2'h0 != last_proc_id ? _GEN_61 : init_io_pipe_phv_out_data_33; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_534 = 2'h0 != last_proc_id ? _GEN_62 : init_io_pipe_phv_out_data_34; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_535 = 2'h0 != last_proc_id ? _GEN_63 : init_io_pipe_phv_out_data_35; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_536 = 2'h0 != last_proc_id ? _GEN_64 : init_io_pipe_phv_out_data_36; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_537 = 2'h0 != last_proc_id ? _GEN_65 : init_io_pipe_phv_out_data_37; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_538 = 2'h0 != last_proc_id ? _GEN_66 : init_io_pipe_phv_out_data_38; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_539 = 2'h0 != last_proc_id ? _GEN_67 : init_io_pipe_phv_out_data_39; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_540 = 2'h0 != last_proc_id ? _GEN_68 : init_io_pipe_phv_out_data_40; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_541 = 2'h0 != last_proc_id ? _GEN_69 : init_io_pipe_phv_out_data_41; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_542 = 2'h0 != last_proc_id ? _GEN_70 : init_io_pipe_phv_out_data_42; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_543 = 2'h0 != last_proc_id ? _GEN_71 : init_io_pipe_phv_out_data_43; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_544 = 2'h0 != last_proc_id ? _GEN_72 : init_io_pipe_phv_out_data_44; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_545 = 2'h0 != last_proc_id ? _GEN_73 : init_io_pipe_phv_out_data_45; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_546 = 2'h0 != last_proc_id ? _GEN_74 : init_io_pipe_phv_out_data_46; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_547 = 2'h0 != last_proc_id ? _GEN_75 : init_io_pipe_phv_out_data_47; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_548 = 2'h0 != last_proc_id ? _GEN_76 : init_io_pipe_phv_out_data_48; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_549 = 2'h0 != last_proc_id ? _GEN_77 : init_io_pipe_phv_out_data_49; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_550 = 2'h0 != last_proc_id ? _GEN_78 : init_io_pipe_phv_out_data_50; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_551 = 2'h0 != last_proc_id ? _GEN_79 : init_io_pipe_phv_out_data_51; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_552 = 2'h0 != last_proc_id ? _GEN_80 : init_io_pipe_phv_out_data_52; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_553 = 2'h0 != last_proc_id ? _GEN_81 : init_io_pipe_phv_out_data_53; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_554 = 2'h0 != last_proc_id ? _GEN_82 : init_io_pipe_phv_out_data_54; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_555 = 2'h0 != last_proc_id ? _GEN_83 : init_io_pipe_phv_out_data_55; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_556 = 2'h0 != last_proc_id ? _GEN_84 : init_io_pipe_phv_out_data_56; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_557 = 2'h0 != last_proc_id ? _GEN_85 : init_io_pipe_phv_out_data_57; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_558 = 2'h0 != last_proc_id ? _GEN_86 : init_io_pipe_phv_out_data_58; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_559 = 2'h0 != last_proc_id ? _GEN_87 : init_io_pipe_phv_out_data_59; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_560 = 2'h0 != last_proc_id ? _GEN_88 : init_io_pipe_phv_out_data_60; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_561 = 2'h0 != last_proc_id ? _GEN_89 : init_io_pipe_phv_out_data_61; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_562 = 2'h0 != last_proc_id ? _GEN_90 : init_io_pipe_phv_out_data_62; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_563 = 2'h0 != last_proc_id ? _GEN_91 : init_io_pipe_phv_out_data_63; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_564 = 2'h0 != last_proc_id ? _GEN_92 : init_io_pipe_phv_out_data_64; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_565 = 2'h0 != last_proc_id ? _GEN_93 : init_io_pipe_phv_out_data_65; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_566 = 2'h0 != last_proc_id ? _GEN_94 : init_io_pipe_phv_out_data_66; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_567 = 2'h0 != last_proc_id ? _GEN_95 : init_io_pipe_phv_out_data_67; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_568 = 2'h0 != last_proc_id ? _GEN_96 : init_io_pipe_phv_out_data_68; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_569 = 2'h0 != last_proc_id ? _GEN_97 : init_io_pipe_phv_out_data_69; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_570 = 2'h0 != last_proc_id ? _GEN_98 : init_io_pipe_phv_out_data_70; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_571 = 2'h0 != last_proc_id ? _GEN_99 : init_io_pipe_phv_out_data_71; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_572 = 2'h0 != last_proc_id ? _GEN_100 : init_io_pipe_phv_out_data_72; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_573 = 2'h0 != last_proc_id ? _GEN_101 : init_io_pipe_phv_out_data_73; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_574 = 2'h0 != last_proc_id ? _GEN_102 : init_io_pipe_phv_out_data_74; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_575 = 2'h0 != last_proc_id ? _GEN_103 : init_io_pipe_phv_out_data_75; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_576 = 2'h0 != last_proc_id ? _GEN_104 : init_io_pipe_phv_out_data_76; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_577 = 2'h0 != last_proc_id ? _GEN_105 : init_io_pipe_phv_out_data_77; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_578 = 2'h0 != last_proc_id ? _GEN_106 : init_io_pipe_phv_out_data_78; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_579 = 2'h0 != last_proc_id ? _GEN_107 : init_io_pipe_phv_out_data_79; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_580 = 2'h0 != last_proc_id ? _GEN_108 : init_io_pipe_phv_out_data_80; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_581 = 2'h0 != last_proc_id ? _GEN_109 : init_io_pipe_phv_out_data_81; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_582 = 2'h0 != last_proc_id ? _GEN_110 : init_io_pipe_phv_out_data_82; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_583 = 2'h0 != last_proc_id ? _GEN_111 : init_io_pipe_phv_out_data_83; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_584 = 2'h0 != last_proc_id ? _GEN_112 : init_io_pipe_phv_out_data_84; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_585 = 2'h0 != last_proc_id ? _GEN_113 : init_io_pipe_phv_out_data_85; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_586 = 2'h0 != last_proc_id ? _GEN_114 : init_io_pipe_phv_out_data_86; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_587 = 2'h0 != last_proc_id ? _GEN_115 : init_io_pipe_phv_out_data_87; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_588 = 2'h0 != last_proc_id ? _GEN_116 : init_io_pipe_phv_out_data_88; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_589 = 2'h0 != last_proc_id ? _GEN_117 : init_io_pipe_phv_out_data_89; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_590 = 2'h0 != last_proc_id ? _GEN_118 : init_io_pipe_phv_out_data_90; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_591 = 2'h0 != last_proc_id ? _GEN_119 : init_io_pipe_phv_out_data_91; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_592 = 2'h0 != last_proc_id ? _GEN_120 : init_io_pipe_phv_out_data_92; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_593 = 2'h0 != last_proc_id ? _GEN_121 : init_io_pipe_phv_out_data_93; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_594 = 2'h0 != last_proc_id ? _GEN_122 : init_io_pipe_phv_out_data_94; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_595 = 2'h0 != last_proc_id ? _GEN_123 : init_io_pipe_phv_out_data_95; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire  _GEN_596 = 2'h0 != last_proc_id ? _GEN_124 : 2'h1 == first_proc_id; // @[ipsa.scala 94:65 ipsa.scala 89:51]
  wire  _GEN_597 = 2'h0 != last_proc_id & _GEN_125; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [1:0] _GEN_598 = 2'h0 != last_proc_id ? _GEN_126 : init_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_599 = 2'h0 != last_proc_id ? _GEN_127 : init_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_600 = 2'h0 != last_proc_id ? _GEN_128 : init_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_601 = 2'h0 != last_proc_id ? _GEN_129 : init_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_602 = 2'h0 != last_proc_id ? _GEN_130 : init_io_pipe_phv_out_header_0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_603 = 2'h0 != last_proc_id ? _GEN_131 : init_io_pipe_phv_out_header_1; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_604 = 2'h0 != last_proc_id ? _GEN_132 : init_io_pipe_phv_out_header_2; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_605 = 2'h0 != last_proc_id ? _GEN_133 : init_io_pipe_phv_out_header_3; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_606 = 2'h0 != last_proc_id ? _GEN_134 : init_io_pipe_phv_out_header_4; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_607 = 2'h0 != last_proc_id ? _GEN_135 : init_io_pipe_phv_out_header_5; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_608 = 2'h0 != last_proc_id ? _GEN_136 : init_io_pipe_phv_out_header_6; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_609 = 2'h0 != last_proc_id ? _GEN_137 : init_io_pipe_phv_out_header_7; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_610 = 2'h0 != last_proc_id ? _GEN_138 : init_io_pipe_phv_out_header_8; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_611 = 2'h0 != last_proc_id ? _GEN_139 : init_io_pipe_phv_out_header_9; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_612 = 2'h0 != last_proc_id ? _GEN_140 : init_io_pipe_phv_out_header_10; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_613 = 2'h0 != last_proc_id ? _GEN_141 : init_io_pipe_phv_out_header_11; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_614 = 2'h0 != last_proc_id ? _GEN_142 : init_io_pipe_phv_out_header_12; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_615 = 2'h0 != last_proc_id ? _GEN_143 : init_io_pipe_phv_out_header_13; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_616 = 2'h0 != last_proc_id ? _GEN_144 : init_io_pipe_phv_out_header_14; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_617 = 2'h0 != last_proc_id ? _GEN_145 : init_io_pipe_phv_out_header_15; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_618 = 2'h0 != last_proc_id ? _GEN_146 : init_io_pipe_phv_out_data_0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_619 = 2'h0 != last_proc_id ? _GEN_147 : init_io_pipe_phv_out_data_1; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_620 = 2'h0 != last_proc_id ? _GEN_148 : init_io_pipe_phv_out_data_2; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_621 = 2'h0 != last_proc_id ? _GEN_149 : init_io_pipe_phv_out_data_3; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_622 = 2'h0 != last_proc_id ? _GEN_150 : init_io_pipe_phv_out_data_4; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_623 = 2'h0 != last_proc_id ? _GEN_151 : init_io_pipe_phv_out_data_5; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_624 = 2'h0 != last_proc_id ? _GEN_152 : init_io_pipe_phv_out_data_6; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_625 = 2'h0 != last_proc_id ? _GEN_153 : init_io_pipe_phv_out_data_7; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_626 = 2'h0 != last_proc_id ? _GEN_154 : init_io_pipe_phv_out_data_8; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_627 = 2'h0 != last_proc_id ? _GEN_155 : init_io_pipe_phv_out_data_9; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_628 = 2'h0 != last_proc_id ? _GEN_156 : init_io_pipe_phv_out_data_10; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_629 = 2'h0 != last_proc_id ? _GEN_157 : init_io_pipe_phv_out_data_11; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_630 = 2'h0 != last_proc_id ? _GEN_158 : init_io_pipe_phv_out_data_12; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_631 = 2'h0 != last_proc_id ? _GEN_159 : init_io_pipe_phv_out_data_13; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_632 = 2'h0 != last_proc_id ? _GEN_160 : init_io_pipe_phv_out_data_14; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_633 = 2'h0 != last_proc_id ? _GEN_161 : init_io_pipe_phv_out_data_15; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_634 = 2'h0 != last_proc_id ? _GEN_162 : init_io_pipe_phv_out_data_16; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_635 = 2'h0 != last_proc_id ? _GEN_163 : init_io_pipe_phv_out_data_17; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_636 = 2'h0 != last_proc_id ? _GEN_164 : init_io_pipe_phv_out_data_18; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_637 = 2'h0 != last_proc_id ? _GEN_165 : init_io_pipe_phv_out_data_19; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_638 = 2'h0 != last_proc_id ? _GEN_166 : init_io_pipe_phv_out_data_20; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_639 = 2'h0 != last_proc_id ? _GEN_167 : init_io_pipe_phv_out_data_21; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_640 = 2'h0 != last_proc_id ? _GEN_168 : init_io_pipe_phv_out_data_22; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_641 = 2'h0 != last_proc_id ? _GEN_169 : init_io_pipe_phv_out_data_23; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_642 = 2'h0 != last_proc_id ? _GEN_170 : init_io_pipe_phv_out_data_24; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_643 = 2'h0 != last_proc_id ? _GEN_171 : init_io_pipe_phv_out_data_25; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_644 = 2'h0 != last_proc_id ? _GEN_172 : init_io_pipe_phv_out_data_26; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_645 = 2'h0 != last_proc_id ? _GEN_173 : init_io_pipe_phv_out_data_27; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_646 = 2'h0 != last_proc_id ? _GEN_174 : init_io_pipe_phv_out_data_28; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_647 = 2'h0 != last_proc_id ? _GEN_175 : init_io_pipe_phv_out_data_29; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_648 = 2'h0 != last_proc_id ? _GEN_176 : init_io_pipe_phv_out_data_30; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_649 = 2'h0 != last_proc_id ? _GEN_177 : init_io_pipe_phv_out_data_31; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_650 = 2'h0 != last_proc_id ? _GEN_178 : init_io_pipe_phv_out_data_32; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_651 = 2'h0 != last_proc_id ? _GEN_179 : init_io_pipe_phv_out_data_33; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_652 = 2'h0 != last_proc_id ? _GEN_180 : init_io_pipe_phv_out_data_34; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_653 = 2'h0 != last_proc_id ? _GEN_181 : init_io_pipe_phv_out_data_35; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_654 = 2'h0 != last_proc_id ? _GEN_182 : init_io_pipe_phv_out_data_36; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_655 = 2'h0 != last_proc_id ? _GEN_183 : init_io_pipe_phv_out_data_37; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_656 = 2'h0 != last_proc_id ? _GEN_184 : init_io_pipe_phv_out_data_38; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_657 = 2'h0 != last_proc_id ? _GEN_185 : init_io_pipe_phv_out_data_39; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_658 = 2'h0 != last_proc_id ? _GEN_186 : init_io_pipe_phv_out_data_40; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_659 = 2'h0 != last_proc_id ? _GEN_187 : init_io_pipe_phv_out_data_41; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_660 = 2'h0 != last_proc_id ? _GEN_188 : init_io_pipe_phv_out_data_42; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_661 = 2'h0 != last_proc_id ? _GEN_189 : init_io_pipe_phv_out_data_43; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_662 = 2'h0 != last_proc_id ? _GEN_190 : init_io_pipe_phv_out_data_44; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_663 = 2'h0 != last_proc_id ? _GEN_191 : init_io_pipe_phv_out_data_45; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_664 = 2'h0 != last_proc_id ? _GEN_192 : init_io_pipe_phv_out_data_46; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_665 = 2'h0 != last_proc_id ? _GEN_193 : init_io_pipe_phv_out_data_47; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_666 = 2'h0 != last_proc_id ? _GEN_194 : init_io_pipe_phv_out_data_48; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_667 = 2'h0 != last_proc_id ? _GEN_195 : init_io_pipe_phv_out_data_49; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_668 = 2'h0 != last_proc_id ? _GEN_196 : init_io_pipe_phv_out_data_50; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_669 = 2'h0 != last_proc_id ? _GEN_197 : init_io_pipe_phv_out_data_51; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_670 = 2'h0 != last_proc_id ? _GEN_198 : init_io_pipe_phv_out_data_52; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_671 = 2'h0 != last_proc_id ? _GEN_199 : init_io_pipe_phv_out_data_53; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_672 = 2'h0 != last_proc_id ? _GEN_200 : init_io_pipe_phv_out_data_54; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_673 = 2'h0 != last_proc_id ? _GEN_201 : init_io_pipe_phv_out_data_55; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_674 = 2'h0 != last_proc_id ? _GEN_202 : init_io_pipe_phv_out_data_56; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_675 = 2'h0 != last_proc_id ? _GEN_203 : init_io_pipe_phv_out_data_57; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_676 = 2'h0 != last_proc_id ? _GEN_204 : init_io_pipe_phv_out_data_58; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_677 = 2'h0 != last_proc_id ? _GEN_205 : init_io_pipe_phv_out_data_59; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_678 = 2'h0 != last_proc_id ? _GEN_206 : init_io_pipe_phv_out_data_60; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_679 = 2'h0 != last_proc_id ? _GEN_207 : init_io_pipe_phv_out_data_61; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_680 = 2'h0 != last_proc_id ? _GEN_208 : init_io_pipe_phv_out_data_62; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_681 = 2'h0 != last_proc_id ? _GEN_209 : init_io_pipe_phv_out_data_63; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_682 = 2'h0 != last_proc_id ? _GEN_210 : init_io_pipe_phv_out_data_64; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_683 = 2'h0 != last_proc_id ? _GEN_211 : init_io_pipe_phv_out_data_65; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_684 = 2'h0 != last_proc_id ? _GEN_212 : init_io_pipe_phv_out_data_66; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_685 = 2'h0 != last_proc_id ? _GEN_213 : init_io_pipe_phv_out_data_67; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_686 = 2'h0 != last_proc_id ? _GEN_214 : init_io_pipe_phv_out_data_68; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_687 = 2'h0 != last_proc_id ? _GEN_215 : init_io_pipe_phv_out_data_69; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_688 = 2'h0 != last_proc_id ? _GEN_216 : init_io_pipe_phv_out_data_70; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_689 = 2'h0 != last_proc_id ? _GEN_217 : init_io_pipe_phv_out_data_71; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_690 = 2'h0 != last_proc_id ? _GEN_218 : init_io_pipe_phv_out_data_72; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_691 = 2'h0 != last_proc_id ? _GEN_219 : init_io_pipe_phv_out_data_73; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_692 = 2'h0 != last_proc_id ? _GEN_220 : init_io_pipe_phv_out_data_74; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_693 = 2'h0 != last_proc_id ? _GEN_221 : init_io_pipe_phv_out_data_75; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_694 = 2'h0 != last_proc_id ? _GEN_222 : init_io_pipe_phv_out_data_76; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_695 = 2'h0 != last_proc_id ? _GEN_223 : init_io_pipe_phv_out_data_77; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_696 = 2'h0 != last_proc_id ? _GEN_224 : init_io_pipe_phv_out_data_78; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_697 = 2'h0 != last_proc_id ? _GEN_225 : init_io_pipe_phv_out_data_79; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_698 = 2'h0 != last_proc_id ? _GEN_226 : init_io_pipe_phv_out_data_80; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_699 = 2'h0 != last_proc_id ? _GEN_227 : init_io_pipe_phv_out_data_81; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_700 = 2'h0 != last_proc_id ? _GEN_228 : init_io_pipe_phv_out_data_82; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_701 = 2'h0 != last_proc_id ? _GEN_229 : init_io_pipe_phv_out_data_83; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_702 = 2'h0 != last_proc_id ? _GEN_230 : init_io_pipe_phv_out_data_84; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_703 = 2'h0 != last_proc_id ? _GEN_231 : init_io_pipe_phv_out_data_85; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_704 = 2'h0 != last_proc_id ? _GEN_232 : init_io_pipe_phv_out_data_86; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_705 = 2'h0 != last_proc_id ? _GEN_233 : init_io_pipe_phv_out_data_87; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_706 = 2'h0 != last_proc_id ? _GEN_234 : init_io_pipe_phv_out_data_88; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_707 = 2'h0 != last_proc_id ? _GEN_235 : init_io_pipe_phv_out_data_89; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_708 = 2'h0 != last_proc_id ? _GEN_236 : init_io_pipe_phv_out_data_90; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_709 = 2'h0 != last_proc_id ? _GEN_237 : init_io_pipe_phv_out_data_91; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_710 = 2'h0 != last_proc_id ? _GEN_238 : init_io_pipe_phv_out_data_92; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_711 = 2'h0 != last_proc_id ? _GEN_239 : init_io_pipe_phv_out_data_93; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_712 = 2'h0 != last_proc_id ? _GEN_240 : init_io_pipe_phv_out_data_94; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_713 = 2'h0 != last_proc_id ? _GEN_241 : init_io_pipe_phv_out_data_95; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire  _GEN_714 = 2'h0 != last_proc_id ? _GEN_242 : 2'h2 == first_proc_id; // @[ipsa.scala 94:65 ipsa.scala 89:51]
  wire  _GEN_715 = 2'h0 != last_proc_id & _GEN_243; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [1:0] _GEN_716 = 2'h0 != last_proc_id ? _GEN_244 : init_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_717 = 2'h0 != last_proc_id ? _GEN_245 : init_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_718 = 2'h0 != last_proc_id ? _GEN_246 : init_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_719 = 2'h0 != last_proc_id ? _GEN_247 : init_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_720 = 2'h0 != last_proc_id ? _GEN_248 : init_io_pipe_phv_out_header_0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_721 = 2'h0 != last_proc_id ? _GEN_249 : init_io_pipe_phv_out_header_1; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_722 = 2'h0 != last_proc_id ? _GEN_250 : init_io_pipe_phv_out_header_2; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_723 = 2'h0 != last_proc_id ? _GEN_251 : init_io_pipe_phv_out_header_3; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_724 = 2'h0 != last_proc_id ? _GEN_252 : init_io_pipe_phv_out_header_4; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_725 = 2'h0 != last_proc_id ? _GEN_253 : init_io_pipe_phv_out_header_5; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_726 = 2'h0 != last_proc_id ? _GEN_254 : init_io_pipe_phv_out_header_6; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_727 = 2'h0 != last_proc_id ? _GEN_255 : init_io_pipe_phv_out_header_7; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_728 = 2'h0 != last_proc_id ? _GEN_256 : init_io_pipe_phv_out_header_8; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_729 = 2'h0 != last_proc_id ? _GEN_257 : init_io_pipe_phv_out_header_9; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_730 = 2'h0 != last_proc_id ? _GEN_258 : init_io_pipe_phv_out_header_10; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_731 = 2'h0 != last_proc_id ? _GEN_259 : init_io_pipe_phv_out_header_11; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_732 = 2'h0 != last_proc_id ? _GEN_260 : init_io_pipe_phv_out_header_12; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_733 = 2'h0 != last_proc_id ? _GEN_261 : init_io_pipe_phv_out_header_13; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_734 = 2'h0 != last_proc_id ? _GEN_262 : init_io_pipe_phv_out_header_14; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_735 = 2'h0 != last_proc_id ? _GEN_263 : init_io_pipe_phv_out_header_15; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_736 = 2'h0 != last_proc_id ? _GEN_264 : init_io_pipe_phv_out_data_0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_737 = 2'h0 != last_proc_id ? _GEN_265 : init_io_pipe_phv_out_data_1; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_738 = 2'h0 != last_proc_id ? _GEN_266 : init_io_pipe_phv_out_data_2; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_739 = 2'h0 != last_proc_id ? _GEN_267 : init_io_pipe_phv_out_data_3; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_740 = 2'h0 != last_proc_id ? _GEN_268 : init_io_pipe_phv_out_data_4; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_741 = 2'h0 != last_proc_id ? _GEN_269 : init_io_pipe_phv_out_data_5; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_742 = 2'h0 != last_proc_id ? _GEN_270 : init_io_pipe_phv_out_data_6; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_743 = 2'h0 != last_proc_id ? _GEN_271 : init_io_pipe_phv_out_data_7; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_744 = 2'h0 != last_proc_id ? _GEN_272 : init_io_pipe_phv_out_data_8; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_745 = 2'h0 != last_proc_id ? _GEN_273 : init_io_pipe_phv_out_data_9; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_746 = 2'h0 != last_proc_id ? _GEN_274 : init_io_pipe_phv_out_data_10; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_747 = 2'h0 != last_proc_id ? _GEN_275 : init_io_pipe_phv_out_data_11; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_748 = 2'h0 != last_proc_id ? _GEN_276 : init_io_pipe_phv_out_data_12; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_749 = 2'h0 != last_proc_id ? _GEN_277 : init_io_pipe_phv_out_data_13; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_750 = 2'h0 != last_proc_id ? _GEN_278 : init_io_pipe_phv_out_data_14; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_751 = 2'h0 != last_proc_id ? _GEN_279 : init_io_pipe_phv_out_data_15; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_752 = 2'h0 != last_proc_id ? _GEN_280 : init_io_pipe_phv_out_data_16; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_753 = 2'h0 != last_proc_id ? _GEN_281 : init_io_pipe_phv_out_data_17; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_754 = 2'h0 != last_proc_id ? _GEN_282 : init_io_pipe_phv_out_data_18; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_755 = 2'h0 != last_proc_id ? _GEN_283 : init_io_pipe_phv_out_data_19; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_756 = 2'h0 != last_proc_id ? _GEN_284 : init_io_pipe_phv_out_data_20; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_757 = 2'h0 != last_proc_id ? _GEN_285 : init_io_pipe_phv_out_data_21; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_758 = 2'h0 != last_proc_id ? _GEN_286 : init_io_pipe_phv_out_data_22; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_759 = 2'h0 != last_proc_id ? _GEN_287 : init_io_pipe_phv_out_data_23; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_760 = 2'h0 != last_proc_id ? _GEN_288 : init_io_pipe_phv_out_data_24; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_761 = 2'h0 != last_proc_id ? _GEN_289 : init_io_pipe_phv_out_data_25; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_762 = 2'h0 != last_proc_id ? _GEN_290 : init_io_pipe_phv_out_data_26; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_763 = 2'h0 != last_proc_id ? _GEN_291 : init_io_pipe_phv_out_data_27; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_764 = 2'h0 != last_proc_id ? _GEN_292 : init_io_pipe_phv_out_data_28; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_765 = 2'h0 != last_proc_id ? _GEN_293 : init_io_pipe_phv_out_data_29; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_766 = 2'h0 != last_proc_id ? _GEN_294 : init_io_pipe_phv_out_data_30; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_767 = 2'h0 != last_proc_id ? _GEN_295 : init_io_pipe_phv_out_data_31; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_768 = 2'h0 != last_proc_id ? _GEN_296 : init_io_pipe_phv_out_data_32; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_769 = 2'h0 != last_proc_id ? _GEN_297 : init_io_pipe_phv_out_data_33; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_770 = 2'h0 != last_proc_id ? _GEN_298 : init_io_pipe_phv_out_data_34; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_771 = 2'h0 != last_proc_id ? _GEN_299 : init_io_pipe_phv_out_data_35; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_772 = 2'h0 != last_proc_id ? _GEN_300 : init_io_pipe_phv_out_data_36; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_773 = 2'h0 != last_proc_id ? _GEN_301 : init_io_pipe_phv_out_data_37; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_774 = 2'h0 != last_proc_id ? _GEN_302 : init_io_pipe_phv_out_data_38; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_775 = 2'h0 != last_proc_id ? _GEN_303 : init_io_pipe_phv_out_data_39; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_776 = 2'h0 != last_proc_id ? _GEN_304 : init_io_pipe_phv_out_data_40; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_777 = 2'h0 != last_proc_id ? _GEN_305 : init_io_pipe_phv_out_data_41; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_778 = 2'h0 != last_proc_id ? _GEN_306 : init_io_pipe_phv_out_data_42; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_779 = 2'h0 != last_proc_id ? _GEN_307 : init_io_pipe_phv_out_data_43; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_780 = 2'h0 != last_proc_id ? _GEN_308 : init_io_pipe_phv_out_data_44; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_781 = 2'h0 != last_proc_id ? _GEN_309 : init_io_pipe_phv_out_data_45; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_782 = 2'h0 != last_proc_id ? _GEN_310 : init_io_pipe_phv_out_data_46; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_783 = 2'h0 != last_proc_id ? _GEN_311 : init_io_pipe_phv_out_data_47; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_784 = 2'h0 != last_proc_id ? _GEN_312 : init_io_pipe_phv_out_data_48; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_785 = 2'h0 != last_proc_id ? _GEN_313 : init_io_pipe_phv_out_data_49; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_786 = 2'h0 != last_proc_id ? _GEN_314 : init_io_pipe_phv_out_data_50; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_787 = 2'h0 != last_proc_id ? _GEN_315 : init_io_pipe_phv_out_data_51; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_788 = 2'h0 != last_proc_id ? _GEN_316 : init_io_pipe_phv_out_data_52; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_789 = 2'h0 != last_proc_id ? _GEN_317 : init_io_pipe_phv_out_data_53; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_790 = 2'h0 != last_proc_id ? _GEN_318 : init_io_pipe_phv_out_data_54; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_791 = 2'h0 != last_proc_id ? _GEN_319 : init_io_pipe_phv_out_data_55; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_792 = 2'h0 != last_proc_id ? _GEN_320 : init_io_pipe_phv_out_data_56; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_793 = 2'h0 != last_proc_id ? _GEN_321 : init_io_pipe_phv_out_data_57; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_794 = 2'h0 != last_proc_id ? _GEN_322 : init_io_pipe_phv_out_data_58; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_795 = 2'h0 != last_proc_id ? _GEN_323 : init_io_pipe_phv_out_data_59; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_796 = 2'h0 != last_proc_id ? _GEN_324 : init_io_pipe_phv_out_data_60; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_797 = 2'h0 != last_proc_id ? _GEN_325 : init_io_pipe_phv_out_data_61; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_798 = 2'h0 != last_proc_id ? _GEN_326 : init_io_pipe_phv_out_data_62; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_799 = 2'h0 != last_proc_id ? _GEN_327 : init_io_pipe_phv_out_data_63; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_800 = 2'h0 != last_proc_id ? _GEN_328 : init_io_pipe_phv_out_data_64; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_801 = 2'h0 != last_proc_id ? _GEN_329 : init_io_pipe_phv_out_data_65; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_802 = 2'h0 != last_proc_id ? _GEN_330 : init_io_pipe_phv_out_data_66; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_803 = 2'h0 != last_proc_id ? _GEN_331 : init_io_pipe_phv_out_data_67; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_804 = 2'h0 != last_proc_id ? _GEN_332 : init_io_pipe_phv_out_data_68; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_805 = 2'h0 != last_proc_id ? _GEN_333 : init_io_pipe_phv_out_data_69; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_806 = 2'h0 != last_proc_id ? _GEN_334 : init_io_pipe_phv_out_data_70; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_807 = 2'h0 != last_proc_id ? _GEN_335 : init_io_pipe_phv_out_data_71; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_808 = 2'h0 != last_proc_id ? _GEN_336 : init_io_pipe_phv_out_data_72; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_809 = 2'h0 != last_proc_id ? _GEN_337 : init_io_pipe_phv_out_data_73; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_810 = 2'h0 != last_proc_id ? _GEN_338 : init_io_pipe_phv_out_data_74; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_811 = 2'h0 != last_proc_id ? _GEN_339 : init_io_pipe_phv_out_data_75; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_812 = 2'h0 != last_proc_id ? _GEN_340 : init_io_pipe_phv_out_data_76; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_813 = 2'h0 != last_proc_id ? _GEN_341 : init_io_pipe_phv_out_data_77; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_814 = 2'h0 != last_proc_id ? _GEN_342 : init_io_pipe_phv_out_data_78; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_815 = 2'h0 != last_proc_id ? _GEN_343 : init_io_pipe_phv_out_data_79; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_816 = 2'h0 != last_proc_id ? _GEN_344 : init_io_pipe_phv_out_data_80; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_817 = 2'h0 != last_proc_id ? _GEN_345 : init_io_pipe_phv_out_data_81; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_818 = 2'h0 != last_proc_id ? _GEN_346 : init_io_pipe_phv_out_data_82; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_819 = 2'h0 != last_proc_id ? _GEN_347 : init_io_pipe_phv_out_data_83; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_820 = 2'h0 != last_proc_id ? _GEN_348 : init_io_pipe_phv_out_data_84; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_821 = 2'h0 != last_proc_id ? _GEN_349 : init_io_pipe_phv_out_data_85; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_822 = 2'h0 != last_proc_id ? _GEN_350 : init_io_pipe_phv_out_data_86; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_823 = 2'h0 != last_proc_id ? _GEN_351 : init_io_pipe_phv_out_data_87; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_824 = 2'h0 != last_proc_id ? _GEN_352 : init_io_pipe_phv_out_data_88; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_825 = 2'h0 != last_proc_id ? _GEN_353 : init_io_pipe_phv_out_data_89; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_826 = 2'h0 != last_proc_id ? _GEN_354 : init_io_pipe_phv_out_data_90; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_827 = 2'h0 != last_proc_id ? _GEN_355 : init_io_pipe_phv_out_data_91; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_828 = 2'h0 != last_proc_id ? _GEN_356 : init_io_pipe_phv_out_data_92; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_829 = 2'h0 != last_proc_id ? _GEN_357 : init_io_pipe_phv_out_data_93; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_830 = 2'h0 != last_proc_id ? _GEN_358 : init_io_pipe_phv_out_data_94; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_831 = 2'h0 != last_proc_id ? _GEN_359 : init_io_pipe_phv_out_data_95; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire  _GEN_832 = 2'h0 != last_proc_id ? _GEN_360 : 2'h3 == first_proc_id; // @[ipsa.scala 94:65 ipsa.scala 89:51]
  wire  _GEN_833 = 2'h0 != last_proc_id & _GEN_361; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [1:0] _GEN_834 = 2'h0 != last_proc_id ? _GEN_362 : init_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_835 = 2'h0 != last_proc_id ? _GEN_363 : init_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_836 = 2'h0 != last_proc_id ? _GEN_364 : init_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_837 = 2'h0 != last_proc_id ? _GEN_365 : init_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_838 = 2'h0 != last_proc_id ? _GEN_366 : init_io_pipe_phv_out_header_0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_839 = 2'h0 != last_proc_id ? _GEN_367 : init_io_pipe_phv_out_header_1; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_840 = 2'h0 != last_proc_id ? _GEN_368 : init_io_pipe_phv_out_header_2; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_841 = 2'h0 != last_proc_id ? _GEN_369 : init_io_pipe_phv_out_header_3; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_842 = 2'h0 != last_proc_id ? _GEN_370 : init_io_pipe_phv_out_header_4; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_843 = 2'h0 != last_proc_id ? _GEN_371 : init_io_pipe_phv_out_header_5; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_844 = 2'h0 != last_proc_id ? _GEN_372 : init_io_pipe_phv_out_header_6; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_845 = 2'h0 != last_proc_id ? _GEN_373 : init_io_pipe_phv_out_header_7; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_846 = 2'h0 != last_proc_id ? _GEN_374 : init_io_pipe_phv_out_header_8; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_847 = 2'h0 != last_proc_id ? _GEN_375 : init_io_pipe_phv_out_header_9; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_848 = 2'h0 != last_proc_id ? _GEN_376 : init_io_pipe_phv_out_header_10; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_849 = 2'h0 != last_proc_id ? _GEN_377 : init_io_pipe_phv_out_header_11; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_850 = 2'h0 != last_proc_id ? _GEN_378 : init_io_pipe_phv_out_header_12; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_851 = 2'h0 != last_proc_id ? _GEN_379 : init_io_pipe_phv_out_header_13; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_852 = 2'h0 != last_proc_id ? _GEN_380 : init_io_pipe_phv_out_header_14; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [15:0] _GEN_853 = 2'h0 != last_proc_id ? _GEN_381 : init_io_pipe_phv_out_header_15; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_854 = 2'h0 != last_proc_id ? _GEN_382 : init_io_pipe_phv_out_data_0; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_855 = 2'h0 != last_proc_id ? _GEN_383 : init_io_pipe_phv_out_data_1; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_856 = 2'h0 != last_proc_id ? _GEN_384 : init_io_pipe_phv_out_data_2; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_857 = 2'h0 != last_proc_id ? _GEN_385 : init_io_pipe_phv_out_data_3; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_858 = 2'h0 != last_proc_id ? _GEN_386 : init_io_pipe_phv_out_data_4; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_859 = 2'h0 != last_proc_id ? _GEN_387 : init_io_pipe_phv_out_data_5; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_860 = 2'h0 != last_proc_id ? _GEN_388 : init_io_pipe_phv_out_data_6; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_861 = 2'h0 != last_proc_id ? _GEN_389 : init_io_pipe_phv_out_data_7; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_862 = 2'h0 != last_proc_id ? _GEN_390 : init_io_pipe_phv_out_data_8; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_863 = 2'h0 != last_proc_id ? _GEN_391 : init_io_pipe_phv_out_data_9; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_864 = 2'h0 != last_proc_id ? _GEN_392 : init_io_pipe_phv_out_data_10; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_865 = 2'h0 != last_proc_id ? _GEN_393 : init_io_pipe_phv_out_data_11; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_866 = 2'h0 != last_proc_id ? _GEN_394 : init_io_pipe_phv_out_data_12; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_867 = 2'h0 != last_proc_id ? _GEN_395 : init_io_pipe_phv_out_data_13; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_868 = 2'h0 != last_proc_id ? _GEN_396 : init_io_pipe_phv_out_data_14; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_869 = 2'h0 != last_proc_id ? _GEN_397 : init_io_pipe_phv_out_data_15; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_870 = 2'h0 != last_proc_id ? _GEN_398 : init_io_pipe_phv_out_data_16; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_871 = 2'h0 != last_proc_id ? _GEN_399 : init_io_pipe_phv_out_data_17; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_872 = 2'h0 != last_proc_id ? _GEN_400 : init_io_pipe_phv_out_data_18; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_873 = 2'h0 != last_proc_id ? _GEN_401 : init_io_pipe_phv_out_data_19; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_874 = 2'h0 != last_proc_id ? _GEN_402 : init_io_pipe_phv_out_data_20; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_875 = 2'h0 != last_proc_id ? _GEN_403 : init_io_pipe_phv_out_data_21; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_876 = 2'h0 != last_proc_id ? _GEN_404 : init_io_pipe_phv_out_data_22; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_877 = 2'h0 != last_proc_id ? _GEN_405 : init_io_pipe_phv_out_data_23; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_878 = 2'h0 != last_proc_id ? _GEN_406 : init_io_pipe_phv_out_data_24; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_879 = 2'h0 != last_proc_id ? _GEN_407 : init_io_pipe_phv_out_data_25; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_880 = 2'h0 != last_proc_id ? _GEN_408 : init_io_pipe_phv_out_data_26; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_881 = 2'h0 != last_proc_id ? _GEN_409 : init_io_pipe_phv_out_data_27; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_882 = 2'h0 != last_proc_id ? _GEN_410 : init_io_pipe_phv_out_data_28; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_883 = 2'h0 != last_proc_id ? _GEN_411 : init_io_pipe_phv_out_data_29; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_884 = 2'h0 != last_proc_id ? _GEN_412 : init_io_pipe_phv_out_data_30; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_885 = 2'h0 != last_proc_id ? _GEN_413 : init_io_pipe_phv_out_data_31; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_886 = 2'h0 != last_proc_id ? _GEN_414 : init_io_pipe_phv_out_data_32; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_887 = 2'h0 != last_proc_id ? _GEN_415 : init_io_pipe_phv_out_data_33; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_888 = 2'h0 != last_proc_id ? _GEN_416 : init_io_pipe_phv_out_data_34; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_889 = 2'h0 != last_proc_id ? _GEN_417 : init_io_pipe_phv_out_data_35; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_890 = 2'h0 != last_proc_id ? _GEN_418 : init_io_pipe_phv_out_data_36; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_891 = 2'h0 != last_proc_id ? _GEN_419 : init_io_pipe_phv_out_data_37; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_892 = 2'h0 != last_proc_id ? _GEN_420 : init_io_pipe_phv_out_data_38; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_893 = 2'h0 != last_proc_id ? _GEN_421 : init_io_pipe_phv_out_data_39; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_894 = 2'h0 != last_proc_id ? _GEN_422 : init_io_pipe_phv_out_data_40; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_895 = 2'h0 != last_proc_id ? _GEN_423 : init_io_pipe_phv_out_data_41; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_896 = 2'h0 != last_proc_id ? _GEN_424 : init_io_pipe_phv_out_data_42; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_897 = 2'h0 != last_proc_id ? _GEN_425 : init_io_pipe_phv_out_data_43; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_898 = 2'h0 != last_proc_id ? _GEN_426 : init_io_pipe_phv_out_data_44; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_899 = 2'h0 != last_proc_id ? _GEN_427 : init_io_pipe_phv_out_data_45; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_900 = 2'h0 != last_proc_id ? _GEN_428 : init_io_pipe_phv_out_data_46; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_901 = 2'h0 != last_proc_id ? _GEN_429 : init_io_pipe_phv_out_data_47; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_902 = 2'h0 != last_proc_id ? _GEN_430 : init_io_pipe_phv_out_data_48; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_903 = 2'h0 != last_proc_id ? _GEN_431 : init_io_pipe_phv_out_data_49; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_904 = 2'h0 != last_proc_id ? _GEN_432 : init_io_pipe_phv_out_data_50; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_905 = 2'h0 != last_proc_id ? _GEN_433 : init_io_pipe_phv_out_data_51; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_906 = 2'h0 != last_proc_id ? _GEN_434 : init_io_pipe_phv_out_data_52; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_907 = 2'h0 != last_proc_id ? _GEN_435 : init_io_pipe_phv_out_data_53; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_908 = 2'h0 != last_proc_id ? _GEN_436 : init_io_pipe_phv_out_data_54; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_909 = 2'h0 != last_proc_id ? _GEN_437 : init_io_pipe_phv_out_data_55; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_910 = 2'h0 != last_proc_id ? _GEN_438 : init_io_pipe_phv_out_data_56; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_911 = 2'h0 != last_proc_id ? _GEN_439 : init_io_pipe_phv_out_data_57; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_912 = 2'h0 != last_proc_id ? _GEN_440 : init_io_pipe_phv_out_data_58; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_913 = 2'h0 != last_proc_id ? _GEN_441 : init_io_pipe_phv_out_data_59; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_914 = 2'h0 != last_proc_id ? _GEN_442 : init_io_pipe_phv_out_data_60; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_915 = 2'h0 != last_proc_id ? _GEN_443 : init_io_pipe_phv_out_data_61; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_916 = 2'h0 != last_proc_id ? _GEN_444 : init_io_pipe_phv_out_data_62; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_917 = 2'h0 != last_proc_id ? _GEN_445 : init_io_pipe_phv_out_data_63; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_918 = 2'h0 != last_proc_id ? _GEN_446 : init_io_pipe_phv_out_data_64; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_919 = 2'h0 != last_proc_id ? _GEN_447 : init_io_pipe_phv_out_data_65; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_920 = 2'h0 != last_proc_id ? _GEN_448 : init_io_pipe_phv_out_data_66; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_921 = 2'h0 != last_proc_id ? _GEN_449 : init_io_pipe_phv_out_data_67; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_922 = 2'h0 != last_proc_id ? _GEN_450 : init_io_pipe_phv_out_data_68; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_923 = 2'h0 != last_proc_id ? _GEN_451 : init_io_pipe_phv_out_data_69; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_924 = 2'h0 != last_proc_id ? _GEN_452 : init_io_pipe_phv_out_data_70; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_925 = 2'h0 != last_proc_id ? _GEN_453 : init_io_pipe_phv_out_data_71; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_926 = 2'h0 != last_proc_id ? _GEN_454 : init_io_pipe_phv_out_data_72; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_927 = 2'h0 != last_proc_id ? _GEN_455 : init_io_pipe_phv_out_data_73; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_928 = 2'h0 != last_proc_id ? _GEN_456 : init_io_pipe_phv_out_data_74; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_929 = 2'h0 != last_proc_id ? _GEN_457 : init_io_pipe_phv_out_data_75; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_930 = 2'h0 != last_proc_id ? _GEN_458 : init_io_pipe_phv_out_data_76; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_931 = 2'h0 != last_proc_id ? _GEN_459 : init_io_pipe_phv_out_data_77; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_932 = 2'h0 != last_proc_id ? _GEN_460 : init_io_pipe_phv_out_data_78; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_933 = 2'h0 != last_proc_id ? _GEN_461 : init_io_pipe_phv_out_data_79; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_934 = 2'h0 != last_proc_id ? _GEN_462 : init_io_pipe_phv_out_data_80; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_935 = 2'h0 != last_proc_id ? _GEN_463 : init_io_pipe_phv_out_data_81; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_936 = 2'h0 != last_proc_id ? _GEN_464 : init_io_pipe_phv_out_data_82; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_937 = 2'h0 != last_proc_id ? _GEN_465 : init_io_pipe_phv_out_data_83; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_938 = 2'h0 != last_proc_id ? _GEN_466 : init_io_pipe_phv_out_data_84; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_939 = 2'h0 != last_proc_id ? _GEN_467 : init_io_pipe_phv_out_data_85; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_940 = 2'h0 != last_proc_id ? _GEN_468 : init_io_pipe_phv_out_data_86; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_941 = 2'h0 != last_proc_id ? _GEN_469 : init_io_pipe_phv_out_data_87; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_942 = 2'h0 != last_proc_id ? _GEN_470 : init_io_pipe_phv_out_data_88; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_943 = 2'h0 != last_proc_id ? _GEN_471 : init_io_pipe_phv_out_data_89; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_944 = 2'h0 != last_proc_id ? _GEN_472 : init_io_pipe_phv_out_data_90; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_945 = 2'h0 != last_proc_id ? _GEN_473 : init_io_pipe_phv_out_data_91; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_946 = 2'h0 != last_proc_id ? _GEN_474 : init_io_pipe_phv_out_data_92; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_947 = 2'h0 != last_proc_id ? _GEN_475 : init_io_pipe_phv_out_data_93; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_948 = 2'h0 != last_proc_id ? _GEN_476 : init_io_pipe_phv_out_data_94; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire [7:0] _GEN_949 = 2'h0 != last_proc_id ? _GEN_477 : init_io_pipe_phv_out_data_95; // @[ipsa.scala 94:65 ipsa.scala 88:32]
  wire  _GEN_950 = 2'h0 != last_proc_id ? io_pipe_phv_in_is_valid_processor : trans_0_io_pipe_phv_out_is_valid_processor
    ; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire  _GEN_951 = 2'h0 != last_proc_id ? io_pipe_phv_in_next_config_id : trans_0_io_pipe_phv_out_next_config_id; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [1:0] _GEN_952 = 2'h0 != last_proc_id ? io_pipe_phv_in_next_processor_id :
    trans_0_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [15:0] _GEN_953 = 2'h0 != last_proc_id ? io_pipe_phv_in_parse_transition_field :
    trans_0_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_954 = 2'h0 != last_proc_id ? io_pipe_phv_in_parse_current_offset :
    trans_0_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_955 = 2'h0 != last_proc_id ? io_pipe_phv_in_parse_current_state :
    trans_0_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [15:0] _GEN_956 = 2'h0 != last_proc_id ? io_pipe_phv_in_header_0 : trans_0_io_pipe_phv_out_header_0; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [15:0] _GEN_957 = 2'h0 != last_proc_id ? io_pipe_phv_in_header_1 : trans_0_io_pipe_phv_out_header_1; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [15:0] _GEN_958 = 2'h0 != last_proc_id ? io_pipe_phv_in_header_2 : trans_0_io_pipe_phv_out_header_2; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [15:0] _GEN_959 = 2'h0 != last_proc_id ? io_pipe_phv_in_header_3 : trans_0_io_pipe_phv_out_header_3; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [15:0] _GEN_960 = 2'h0 != last_proc_id ? io_pipe_phv_in_header_4 : trans_0_io_pipe_phv_out_header_4; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [15:0] _GEN_961 = 2'h0 != last_proc_id ? io_pipe_phv_in_header_5 : trans_0_io_pipe_phv_out_header_5; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [15:0] _GEN_962 = 2'h0 != last_proc_id ? io_pipe_phv_in_header_6 : trans_0_io_pipe_phv_out_header_6; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [15:0] _GEN_963 = 2'h0 != last_proc_id ? io_pipe_phv_in_header_7 : trans_0_io_pipe_phv_out_header_7; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [15:0] _GEN_964 = 2'h0 != last_proc_id ? io_pipe_phv_in_header_8 : trans_0_io_pipe_phv_out_header_8; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [15:0] _GEN_965 = 2'h0 != last_proc_id ? io_pipe_phv_in_header_9 : trans_0_io_pipe_phv_out_header_9; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [15:0] _GEN_966 = 2'h0 != last_proc_id ? io_pipe_phv_in_header_10 : trans_0_io_pipe_phv_out_header_10; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [15:0] _GEN_967 = 2'h0 != last_proc_id ? io_pipe_phv_in_header_11 : trans_0_io_pipe_phv_out_header_11; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [15:0] _GEN_968 = 2'h0 != last_proc_id ? io_pipe_phv_in_header_12 : trans_0_io_pipe_phv_out_header_12; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [15:0] _GEN_969 = 2'h0 != last_proc_id ? io_pipe_phv_in_header_13 : trans_0_io_pipe_phv_out_header_13; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [15:0] _GEN_970 = 2'h0 != last_proc_id ? io_pipe_phv_in_header_14 : trans_0_io_pipe_phv_out_header_14; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [15:0] _GEN_971 = 2'h0 != last_proc_id ? io_pipe_phv_in_header_15 : trans_0_io_pipe_phv_out_header_15; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_972 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_0 : trans_0_io_pipe_phv_out_data_0; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_973 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_1 : trans_0_io_pipe_phv_out_data_1; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_974 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_2 : trans_0_io_pipe_phv_out_data_2; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_975 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_3 : trans_0_io_pipe_phv_out_data_3; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_976 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_4 : trans_0_io_pipe_phv_out_data_4; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_977 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_5 : trans_0_io_pipe_phv_out_data_5; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_978 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_6 : trans_0_io_pipe_phv_out_data_6; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_979 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_7 : trans_0_io_pipe_phv_out_data_7; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_980 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_8 : trans_0_io_pipe_phv_out_data_8; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_981 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_9 : trans_0_io_pipe_phv_out_data_9; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_982 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_10 : trans_0_io_pipe_phv_out_data_10; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_983 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_11 : trans_0_io_pipe_phv_out_data_11; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_984 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_12 : trans_0_io_pipe_phv_out_data_12; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_985 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_13 : trans_0_io_pipe_phv_out_data_13; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_986 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_14 : trans_0_io_pipe_phv_out_data_14; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_987 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_15 : trans_0_io_pipe_phv_out_data_15; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_988 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_16 : trans_0_io_pipe_phv_out_data_16; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_989 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_17 : trans_0_io_pipe_phv_out_data_17; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_990 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_18 : trans_0_io_pipe_phv_out_data_18; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_991 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_19 : trans_0_io_pipe_phv_out_data_19; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_992 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_20 : trans_0_io_pipe_phv_out_data_20; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_993 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_21 : trans_0_io_pipe_phv_out_data_21; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_994 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_22 : trans_0_io_pipe_phv_out_data_22; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_995 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_23 : trans_0_io_pipe_phv_out_data_23; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_996 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_24 : trans_0_io_pipe_phv_out_data_24; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_997 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_25 : trans_0_io_pipe_phv_out_data_25; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_998 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_26 : trans_0_io_pipe_phv_out_data_26; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_999 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_27 : trans_0_io_pipe_phv_out_data_27; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1000 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_28 : trans_0_io_pipe_phv_out_data_28; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1001 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_29 : trans_0_io_pipe_phv_out_data_29; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1002 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_30 : trans_0_io_pipe_phv_out_data_30; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1003 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_31 : trans_0_io_pipe_phv_out_data_31; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1004 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_32 : trans_0_io_pipe_phv_out_data_32; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1005 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_33 : trans_0_io_pipe_phv_out_data_33; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1006 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_34 : trans_0_io_pipe_phv_out_data_34; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1007 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_35 : trans_0_io_pipe_phv_out_data_35; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1008 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_36 : trans_0_io_pipe_phv_out_data_36; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1009 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_37 : trans_0_io_pipe_phv_out_data_37; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1010 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_38 : trans_0_io_pipe_phv_out_data_38; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1011 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_39 : trans_0_io_pipe_phv_out_data_39; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1012 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_40 : trans_0_io_pipe_phv_out_data_40; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1013 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_41 : trans_0_io_pipe_phv_out_data_41; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1014 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_42 : trans_0_io_pipe_phv_out_data_42; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1015 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_43 : trans_0_io_pipe_phv_out_data_43; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1016 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_44 : trans_0_io_pipe_phv_out_data_44; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1017 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_45 : trans_0_io_pipe_phv_out_data_45; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1018 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_46 : trans_0_io_pipe_phv_out_data_46; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1019 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_47 : trans_0_io_pipe_phv_out_data_47; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1020 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_48 : trans_0_io_pipe_phv_out_data_48; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1021 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_49 : trans_0_io_pipe_phv_out_data_49; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1022 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_50 : trans_0_io_pipe_phv_out_data_50; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1023 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_51 : trans_0_io_pipe_phv_out_data_51; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1024 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_52 : trans_0_io_pipe_phv_out_data_52; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1025 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_53 : trans_0_io_pipe_phv_out_data_53; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1026 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_54 : trans_0_io_pipe_phv_out_data_54; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1027 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_55 : trans_0_io_pipe_phv_out_data_55; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1028 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_56 : trans_0_io_pipe_phv_out_data_56; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1029 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_57 : trans_0_io_pipe_phv_out_data_57; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1030 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_58 : trans_0_io_pipe_phv_out_data_58; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1031 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_59 : trans_0_io_pipe_phv_out_data_59; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1032 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_60 : trans_0_io_pipe_phv_out_data_60; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1033 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_61 : trans_0_io_pipe_phv_out_data_61; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1034 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_62 : trans_0_io_pipe_phv_out_data_62; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1035 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_63 : trans_0_io_pipe_phv_out_data_63; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1036 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_64 : trans_0_io_pipe_phv_out_data_64; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1037 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_65 : trans_0_io_pipe_phv_out_data_65; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1038 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_66 : trans_0_io_pipe_phv_out_data_66; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1039 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_67 : trans_0_io_pipe_phv_out_data_67; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1040 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_68 : trans_0_io_pipe_phv_out_data_68; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1041 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_69 : trans_0_io_pipe_phv_out_data_69; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1042 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_70 : trans_0_io_pipe_phv_out_data_70; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1043 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_71 : trans_0_io_pipe_phv_out_data_71; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1044 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_72 : trans_0_io_pipe_phv_out_data_72; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1045 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_73 : trans_0_io_pipe_phv_out_data_73; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1046 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_74 : trans_0_io_pipe_phv_out_data_74; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1047 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_75 : trans_0_io_pipe_phv_out_data_75; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1048 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_76 : trans_0_io_pipe_phv_out_data_76; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1049 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_77 : trans_0_io_pipe_phv_out_data_77; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1050 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_78 : trans_0_io_pipe_phv_out_data_78; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1051 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_79 : trans_0_io_pipe_phv_out_data_79; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1052 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_80 : trans_0_io_pipe_phv_out_data_80; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1053 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_81 : trans_0_io_pipe_phv_out_data_81; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1054 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_82 : trans_0_io_pipe_phv_out_data_82; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1055 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_83 : trans_0_io_pipe_phv_out_data_83; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1056 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_84 : trans_0_io_pipe_phv_out_data_84; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1057 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_85 : trans_0_io_pipe_phv_out_data_85; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1058 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_86 : trans_0_io_pipe_phv_out_data_86; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1059 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_87 : trans_0_io_pipe_phv_out_data_87; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1060 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_88 : trans_0_io_pipe_phv_out_data_88; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1061 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_89 : trans_0_io_pipe_phv_out_data_89; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1062 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_90 : trans_0_io_pipe_phv_out_data_90; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1063 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_91 : trans_0_io_pipe_phv_out_data_91; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1064 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_92 : trans_0_io_pipe_phv_out_data_92; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1065 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_93 : trans_0_io_pipe_phv_out_data_93; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1066 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_94 : trans_0_io_pipe_phv_out_data_94; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire [7:0] _GEN_1067 = 2'h0 != last_proc_id ? io_pipe_phv_in_data_95 : trans_0_io_pipe_phv_out_data_95; // @[ipsa.scala 94:65 ipsa.scala 86:21 ipsa.scala 101:29]
  wire  _GEN_1068 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_is_valid_processor : _GEN_478; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire  _GEN_1069 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_next_config_id : _GEN_479; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [1:0] _GEN_1070 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_next_processor_id : _GEN_480; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1071 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_parse_transition_field : _GEN_481; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1072 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_parse_current_offset : _GEN_482; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1073 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_parse_current_state : _GEN_483; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1074 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_0 : _GEN_484; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1075 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_1 : _GEN_485; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1076 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_2 : _GEN_486; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1077 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_3 : _GEN_487; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1078 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_4 : _GEN_488; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1079 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_5 : _GEN_489; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1080 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_6 : _GEN_490; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1081 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_7 : _GEN_491; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1082 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_8 : _GEN_492; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1083 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_9 : _GEN_493; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1084 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_10 : _GEN_494; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1085 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_11 : _GEN_495; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1086 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_12 : _GEN_496; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1087 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_13 : _GEN_497; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1088 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_14 : _GEN_498; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1089 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_15 : _GEN_499; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1090 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_0 : _GEN_500; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1091 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_1 : _GEN_501; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1092 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_2 : _GEN_502; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1093 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_3 : _GEN_503; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1094 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_4 : _GEN_504; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1095 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_5 : _GEN_505; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1096 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_6 : _GEN_506; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1097 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_7 : _GEN_507; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1098 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_8 : _GEN_508; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1099 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_9 : _GEN_509; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1100 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_10 : _GEN_510; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1101 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_11 : _GEN_511; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1102 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_12 : _GEN_512; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1103 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_13 : _GEN_513; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1104 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_14 : _GEN_514; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1105 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_15 : _GEN_515; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1106 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_16 : _GEN_516; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1107 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_17 : _GEN_517; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1108 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_18 : _GEN_518; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1109 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_19 : _GEN_519; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1110 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_20 : _GEN_520; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1111 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_21 : _GEN_521; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1112 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_22 : _GEN_522; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1113 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_23 : _GEN_523; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1114 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_24 : _GEN_524; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1115 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_25 : _GEN_525; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1116 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_26 : _GEN_526; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1117 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_27 : _GEN_527; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1118 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_28 : _GEN_528; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1119 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_29 : _GEN_529; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1120 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_30 : _GEN_530; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1121 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_31 : _GEN_531; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1122 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_32 : _GEN_532; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1123 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_33 : _GEN_533; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1124 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_34 : _GEN_534; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1125 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_35 : _GEN_535; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1126 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_36 : _GEN_536; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1127 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_37 : _GEN_537; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1128 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_38 : _GEN_538; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1129 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_39 : _GEN_539; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1130 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_40 : _GEN_540; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1131 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_41 : _GEN_541; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1132 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_42 : _GEN_542; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1133 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_43 : _GEN_543; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1134 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_44 : _GEN_544; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1135 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_45 : _GEN_545; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1136 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_46 : _GEN_546; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1137 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_47 : _GEN_547; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1138 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_48 : _GEN_548; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1139 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_49 : _GEN_549; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1140 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_50 : _GEN_550; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1141 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_51 : _GEN_551; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1142 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_52 : _GEN_552; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1143 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_53 : _GEN_553; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1144 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_54 : _GEN_554; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1145 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_55 : _GEN_555; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1146 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_56 : _GEN_556; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1147 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_57 : _GEN_557; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1148 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_58 : _GEN_558; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1149 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_59 : _GEN_559; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1150 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_60 : _GEN_560; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1151 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_61 : _GEN_561; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1152 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_62 : _GEN_562; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1153 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_63 : _GEN_563; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1154 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_64 : _GEN_564; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1155 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_65 : _GEN_565; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1156 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_66 : _GEN_566; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1157 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_67 : _GEN_567; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1158 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_68 : _GEN_568; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1159 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_69 : _GEN_569; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1160 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_70 : _GEN_570; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1161 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_71 : _GEN_571; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1162 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_72 : _GEN_572; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1163 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_73 : _GEN_573; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1164 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_74 : _GEN_574; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1165 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_75 : _GEN_575; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1166 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_76 : _GEN_576; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1167 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_77 : _GEN_577; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1168 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_78 : _GEN_578; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1169 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_79 : _GEN_579; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1170 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_80 : _GEN_580; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1171 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_81 : _GEN_581; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1172 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_82 : _GEN_582; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1173 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_83 : _GEN_583; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1174 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_84 : _GEN_584; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1175 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_85 : _GEN_585; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1176 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_86 : _GEN_586; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1177 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_87 : _GEN_587; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1178 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_88 : _GEN_588; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1179 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_89 : _GEN_589; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1180 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_90 : _GEN_590; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1181 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_91 : _GEN_591; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1182 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_92 : _GEN_592; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1183 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_93 : _GEN_593; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1184 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_94 : _GEN_594; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1185 = 2'h0 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_95 : _GEN_595; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire  _GEN_1186 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_is_valid_processor : _GEN_596; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire  _GEN_1187 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_next_config_id : _GEN_597; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [1:0] _GEN_1188 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_next_processor_id : _GEN_598; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1189 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_parse_transition_field : _GEN_599; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1190 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_parse_current_offset : _GEN_600; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1191 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_parse_current_state : _GEN_601; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1192 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_0 : _GEN_602; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1193 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_1 : _GEN_603; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1194 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_2 : _GEN_604; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1195 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_3 : _GEN_605; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1196 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_4 : _GEN_606; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1197 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_5 : _GEN_607; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1198 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_6 : _GEN_608; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1199 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_7 : _GEN_609; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1200 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_8 : _GEN_610; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1201 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_9 : _GEN_611; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1202 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_10 : _GEN_612; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1203 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_11 : _GEN_613; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1204 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_12 : _GEN_614; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1205 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_13 : _GEN_615; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1206 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_14 : _GEN_616; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1207 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_15 : _GEN_617; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1208 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_0 : _GEN_618; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1209 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_1 : _GEN_619; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1210 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_2 : _GEN_620; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1211 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_3 : _GEN_621; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1212 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_4 : _GEN_622; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1213 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_5 : _GEN_623; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1214 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_6 : _GEN_624; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1215 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_7 : _GEN_625; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1216 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_8 : _GEN_626; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1217 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_9 : _GEN_627; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1218 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_10 : _GEN_628; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1219 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_11 : _GEN_629; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1220 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_12 : _GEN_630; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1221 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_13 : _GEN_631; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1222 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_14 : _GEN_632; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1223 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_15 : _GEN_633; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1224 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_16 : _GEN_634; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1225 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_17 : _GEN_635; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1226 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_18 : _GEN_636; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1227 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_19 : _GEN_637; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1228 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_20 : _GEN_638; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1229 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_21 : _GEN_639; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1230 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_22 : _GEN_640; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1231 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_23 : _GEN_641; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1232 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_24 : _GEN_642; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1233 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_25 : _GEN_643; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1234 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_26 : _GEN_644; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1235 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_27 : _GEN_645; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1236 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_28 : _GEN_646; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1237 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_29 : _GEN_647; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1238 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_30 : _GEN_648; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1239 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_31 : _GEN_649; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1240 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_32 : _GEN_650; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1241 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_33 : _GEN_651; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1242 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_34 : _GEN_652; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1243 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_35 : _GEN_653; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1244 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_36 : _GEN_654; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1245 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_37 : _GEN_655; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1246 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_38 : _GEN_656; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1247 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_39 : _GEN_657; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1248 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_40 : _GEN_658; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1249 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_41 : _GEN_659; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1250 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_42 : _GEN_660; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1251 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_43 : _GEN_661; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1252 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_44 : _GEN_662; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1253 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_45 : _GEN_663; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1254 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_46 : _GEN_664; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1255 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_47 : _GEN_665; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1256 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_48 : _GEN_666; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1257 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_49 : _GEN_667; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1258 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_50 : _GEN_668; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1259 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_51 : _GEN_669; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1260 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_52 : _GEN_670; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1261 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_53 : _GEN_671; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1262 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_54 : _GEN_672; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1263 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_55 : _GEN_673; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1264 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_56 : _GEN_674; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1265 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_57 : _GEN_675; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1266 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_58 : _GEN_676; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1267 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_59 : _GEN_677; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1268 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_60 : _GEN_678; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1269 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_61 : _GEN_679; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1270 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_62 : _GEN_680; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1271 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_63 : _GEN_681; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1272 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_64 : _GEN_682; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1273 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_65 : _GEN_683; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1274 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_66 : _GEN_684; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1275 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_67 : _GEN_685; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1276 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_68 : _GEN_686; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1277 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_69 : _GEN_687; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1278 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_70 : _GEN_688; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1279 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_71 : _GEN_689; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1280 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_72 : _GEN_690; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1281 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_73 : _GEN_691; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1282 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_74 : _GEN_692; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1283 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_75 : _GEN_693; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1284 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_76 : _GEN_694; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1285 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_77 : _GEN_695; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1286 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_78 : _GEN_696; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1287 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_79 : _GEN_697; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1288 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_80 : _GEN_698; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1289 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_81 : _GEN_699; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1290 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_82 : _GEN_700; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1291 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_83 : _GEN_701; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1292 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_84 : _GEN_702; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1293 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_85 : _GEN_703; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1294 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_86 : _GEN_704; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1295 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_87 : _GEN_705; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1296 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_88 : _GEN_706; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1297 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_89 : _GEN_707; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1298 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_90 : _GEN_708; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1299 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_91 : _GEN_709; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1300 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_92 : _GEN_710; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1301 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_93 : _GEN_711; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1302 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_94 : _GEN_712; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1303 = 2'h1 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_95 : _GEN_713; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire  _GEN_1304 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_is_valid_processor : _GEN_714; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire  _GEN_1305 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_next_config_id : _GEN_715; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [1:0] _GEN_1306 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_next_processor_id : _GEN_716; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1307 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_parse_transition_field : _GEN_717; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1308 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_parse_current_offset : _GEN_718; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1309 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_parse_current_state : _GEN_719; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1310 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_0 : _GEN_720; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1311 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_1 : _GEN_721; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1312 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_2 : _GEN_722; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1313 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_3 : _GEN_723; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1314 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_4 : _GEN_724; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1315 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_5 : _GEN_725; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1316 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_6 : _GEN_726; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1317 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_7 : _GEN_727; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1318 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_8 : _GEN_728; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1319 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_9 : _GEN_729; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1320 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_10 : _GEN_730; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1321 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_11 : _GEN_731; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1322 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_12 : _GEN_732; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1323 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_13 : _GEN_733; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1324 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_14 : _GEN_734; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1325 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_15 : _GEN_735; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1326 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_0 : _GEN_736; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1327 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_1 : _GEN_737; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1328 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_2 : _GEN_738; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1329 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_3 : _GEN_739; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1330 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_4 : _GEN_740; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1331 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_5 : _GEN_741; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1332 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_6 : _GEN_742; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1333 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_7 : _GEN_743; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1334 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_8 : _GEN_744; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1335 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_9 : _GEN_745; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1336 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_10 : _GEN_746; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1337 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_11 : _GEN_747; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1338 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_12 : _GEN_748; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1339 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_13 : _GEN_749; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1340 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_14 : _GEN_750; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1341 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_15 : _GEN_751; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1342 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_16 : _GEN_752; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1343 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_17 : _GEN_753; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1344 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_18 : _GEN_754; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1345 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_19 : _GEN_755; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1346 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_20 : _GEN_756; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1347 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_21 : _GEN_757; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1348 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_22 : _GEN_758; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1349 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_23 : _GEN_759; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1350 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_24 : _GEN_760; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1351 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_25 : _GEN_761; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1352 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_26 : _GEN_762; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1353 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_27 : _GEN_763; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1354 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_28 : _GEN_764; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1355 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_29 : _GEN_765; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1356 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_30 : _GEN_766; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1357 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_31 : _GEN_767; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1358 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_32 : _GEN_768; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1359 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_33 : _GEN_769; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1360 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_34 : _GEN_770; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1361 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_35 : _GEN_771; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1362 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_36 : _GEN_772; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1363 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_37 : _GEN_773; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1364 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_38 : _GEN_774; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1365 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_39 : _GEN_775; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1366 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_40 : _GEN_776; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1367 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_41 : _GEN_777; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1368 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_42 : _GEN_778; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1369 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_43 : _GEN_779; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1370 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_44 : _GEN_780; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1371 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_45 : _GEN_781; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1372 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_46 : _GEN_782; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1373 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_47 : _GEN_783; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1374 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_48 : _GEN_784; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1375 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_49 : _GEN_785; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1376 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_50 : _GEN_786; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1377 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_51 : _GEN_787; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1378 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_52 : _GEN_788; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1379 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_53 : _GEN_789; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1380 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_54 : _GEN_790; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1381 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_55 : _GEN_791; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1382 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_56 : _GEN_792; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1383 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_57 : _GEN_793; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1384 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_58 : _GEN_794; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1385 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_59 : _GEN_795; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1386 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_60 : _GEN_796; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1387 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_61 : _GEN_797; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1388 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_62 : _GEN_798; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1389 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_63 : _GEN_799; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1390 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_64 : _GEN_800; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1391 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_65 : _GEN_801; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1392 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_66 : _GEN_802; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1393 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_67 : _GEN_803; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1394 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_68 : _GEN_804; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1395 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_69 : _GEN_805; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1396 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_70 : _GEN_806; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1397 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_71 : _GEN_807; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1398 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_72 : _GEN_808; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1399 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_73 : _GEN_809; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1400 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_74 : _GEN_810; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1401 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_75 : _GEN_811; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1402 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_76 : _GEN_812; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1403 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_77 : _GEN_813; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1404 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_78 : _GEN_814; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1405 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_79 : _GEN_815; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1406 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_80 : _GEN_816; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1407 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_81 : _GEN_817; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1408 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_82 : _GEN_818; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1409 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_83 : _GEN_819; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1410 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_84 : _GEN_820; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1411 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_85 : _GEN_821; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1412 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_86 : _GEN_822; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1413 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_87 : _GEN_823; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1414 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_88 : _GEN_824; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1415 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_89 : _GEN_825; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1416 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_90 : _GEN_826; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1417 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_91 : _GEN_827; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1418 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_92 : _GEN_828; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1419 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_93 : _GEN_829; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1420 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_94 : _GEN_830; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1421 = 2'h2 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_95 : _GEN_831; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire  _GEN_1422 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_is_valid_processor : _GEN_832; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire  _GEN_1423 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_next_config_id : _GEN_833; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [1:0] _GEN_1424 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_next_processor_id : _GEN_834; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1425 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_parse_transition_field : _GEN_835; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1426 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_parse_current_offset : _GEN_836; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1427 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_parse_current_state : _GEN_837; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1428 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_0 : _GEN_838; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1429 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_1 : _GEN_839; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1430 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_2 : _GEN_840; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1431 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_3 : _GEN_841; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1432 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_4 : _GEN_842; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1433 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_5 : _GEN_843; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1434 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_6 : _GEN_844; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1435 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_7 : _GEN_845; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1436 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_8 : _GEN_846; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1437 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_9 : _GEN_847; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1438 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_10 : _GEN_848; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1439 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_11 : _GEN_849; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1440 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_12 : _GEN_850; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1441 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_13 : _GEN_851; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1442 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_14 : _GEN_852; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_1443 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_header_15 : _GEN_853; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1444 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_0 : _GEN_854; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1445 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_1 : _GEN_855; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1446 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_2 : _GEN_856; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1447 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_3 : _GEN_857; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1448 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_4 : _GEN_858; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1449 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_5 : _GEN_859; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1450 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_6 : _GEN_860; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1451 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_7 : _GEN_861; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1452 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_8 : _GEN_862; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1453 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_9 : _GEN_863; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1454 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_10 : _GEN_864; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1455 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_11 : _GEN_865; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1456 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_12 : _GEN_866; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1457 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_13 : _GEN_867; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1458 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_14 : _GEN_868; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1459 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_15 : _GEN_869; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1460 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_16 : _GEN_870; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1461 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_17 : _GEN_871; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1462 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_18 : _GEN_872; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1463 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_19 : _GEN_873; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1464 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_20 : _GEN_874; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1465 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_21 : _GEN_875; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1466 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_22 : _GEN_876; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1467 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_23 : _GEN_877; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1468 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_24 : _GEN_878; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1469 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_25 : _GEN_879; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1470 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_26 : _GEN_880; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1471 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_27 : _GEN_881; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1472 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_28 : _GEN_882; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1473 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_29 : _GEN_883; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1474 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_30 : _GEN_884; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1475 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_31 : _GEN_885; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1476 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_32 : _GEN_886; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1477 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_33 : _GEN_887; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1478 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_34 : _GEN_888; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1479 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_35 : _GEN_889; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1480 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_36 : _GEN_890; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1481 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_37 : _GEN_891; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1482 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_38 : _GEN_892; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1483 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_39 : _GEN_893; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1484 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_40 : _GEN_894; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1485 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_41 : _GEN_895; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1486 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_42 : _GEN_896; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1487 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_43 : _GEN_897; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1488 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_44 : _GEN_898; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1489 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_45 : _GEN_899; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1490 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_46 : _GEN_900; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1491 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_47 : _GEN_901; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1492 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_48 : _GEN_902; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1493 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_49 : _GEN_903; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1494 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_50 : _GEN_904; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1495 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_51 : _GEN_905; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1496 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_52 : _GEN_906; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1497 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_53 : _GEN_907; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1498 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_54 : _GEN_908; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1499 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_55 : _GEN_909; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1500 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_56 : _GEN_910; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1501 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_57 : _GEN_911; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1502 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_58 : _GEN_912; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1503 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_59 : _GEN_913; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1504 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_60 : _GEN_914; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1505 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_61 : _GEN_915; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1506 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_62 : _GEN_916; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1507 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_63 : _GEN_917; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1508 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_64 : _GEN_918; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1509 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_65 : _GEN_919; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1510 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_66 : _GEN_920; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1511 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_67 : _GEN_921; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1512 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_68 : _GEN_922; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1513 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_69 : _GEN_923; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1514 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_70 : _GEN_924; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1515 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_71 : _GEN_925; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1516 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_72 : _GEN_926; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1517 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_73 : _GEN_927; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1518 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_74 : _GEN_928; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1519 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_75 : _GEN_929; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1520 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_76 : _GEN_930; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1521 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_77 : _GEN_931; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1522 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_78 : _GEN_932; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1523 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_79 : _GEN_933; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1524 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_80 : _GEN_934; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1525 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_81 : _GEN_935; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1526 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_82 : _GEN_936; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1527 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_83 : _GEN_937; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1528 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_84 : _GEN_938; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1529 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_85 : _GEN_939; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1530 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_86 : _GEN_940; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1531 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_87 : _GEN_941; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1532 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_88 : _GEN_942; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1533 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_89 : _GEN_943; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1534 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_90 : _GEN_944; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1535 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_91 : _GEN_945; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1536 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_92 : _GEN_946; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1537 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_93 : _GEN_947; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1538 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_94 : _GEN_948; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_1539 = 2'h3 == next_proc_id_1 ? trans_1_io_pipe_phv_out_data_95 : _GEN_949; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire  _GEN_1540 = 2'h1 != last_proc_id ? _GEN_1068 : _GEN_478; // @[ipsa.scala 94:65]
  wire  _GEN_1541 = 2'h1 != last_proc_id ? _GEN_1069 : _GEN_479; // @[ipsa.scala 94:65]
  wire [1:0] _GEN_1542 = 2'h1 != last_proc_id ? _GEN_1070 : _GEN_480; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1543 = 2'h1 != last_proc_id ? _GEN_1071 : _GEN_481; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1544 = 2'h1 != last_proc_id ? _GEN_1072 : _GEN_482; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1545 = 2'h1 != last_proc_id ? _GEN_1073 : _GEN_483; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1546 = 2'h1 != last_proc_id ? _GEN_1074 : _GEN_484; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1547 = 2'h1 != last_proc_id ? _GEN_1075 : _GEN_485; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1548 = 2'h1 != last_proc_id ? _GEN_1076 : _GEN_486; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1549 = 2'h1 != last_proc_id ? _GEN_1077 : _GEN_487; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1550 = 2'h1 != last_proc_id ? _GEN_1078 : _GEN_488; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1551 = 2'h1 != last_proc_id ? _GEN_1079 : _GEN_489; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1552 = 2'h1 != last_proc_id ? _GEN_1080 : _GEN_490; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1553 = 2'h1 != last_proc_id ? _GEN_1081 : _GEN_491; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1554 = 2'h1 != last_proc_id ? _GEN_1082 : _GEN_492; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1555 = 2'h1 != last_proc_id ? _GEN_1083 : _GEN_493; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1556 = 2'h1 != last_proc_id ? _GEN_1084 : _GEN_494; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1557 = 2'h1 != last_proc_id ? _GEN_1085 : _GEN_495; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1558 = 2'h1 != last_proc_id ? _GEN_1086 : _GEN_496; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1559 = 2'h1 != last_proc_id ? _GEN_1087 : _GEN_497; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1560 = 2'h1 != last_proc_id ? _GEN_1088 : _GEN_498; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1561 = 2'h1 != last_proc_id ? _GEN_1089 : _GEN_499; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1562 = 2'h1 != last_proc_id ? _GEN_1090 : _GEN_500; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1563 = 2'h1 != last_proc_id ? _GEN_1091 : _GEN_501; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1564 = 2'h1 != last_proc_id ? _GEN_1092 : _GEN_502; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1565 = 2'h1 != last_proc_id ? _GEN_1093 : _GEN_503; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1566 = 2'h1 != last_proc_id ? _GEN_1094 : _GEN_504; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1567 = 2'h1 != last_proc_id ? _GEN_1095 : _GEN_505; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1568 = 2'h1 != last_proc_id ? _GEN_1096 : _GEN_506; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1569 = 2'h1 != last_proc_id ? _GEN_1097 : _GEN_507; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1570 = 2'h1 != last_proc_id ? _GEN_1098 : _GEN_508; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1571 = 2'h1 != last_proc_id ? _GEN_1099 : _GEN_509; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1572 = 2'h1 != last_proc_id ? _GEN_1100 : _GEN_510; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1573 = 2'h1 != last_proc_id ? _GEN_1101 : _GEN_511; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1574 = 2'h1 != last_proc_id ? _GEN_1102 : _GEN_512; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1575 = 2'h1 != last_proc_id ? _GEN_1103 : _GEN_513; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1576 = 2'h1 != last_proc_id ? _GEN_1104 : _GEN_514; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1577 = 2'h1 != last_proc_id ? _GEN_1105 : _GEN_515; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1578 = 2'h1 != last_proc_id ? _GEN_1106 : _GEN_516; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1579 = 2'h1 != last_proc_id ? _GEN_1107 : _GEN_517; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1580 = 2'h1 != last_proc_id ? _GEN_1108 : _GEN_518; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1581 = 2'h1 != last_proc_id ? _GEN_1109 : _GEN_519; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1582 = 2'h1 != last_proc_id ? _GEN_1110 : _GEN_520; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1583 = 2'h1 != last_proc_id ? _GEN_1111 : _GEN_521; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1584 = 2'h1 != last_proc_id ? _GEN_1112 : _GEN_522; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1585 = 2'h1 != last_proc_id ? _GEN_1113 : _GEN_523; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1586 = 2'h1 != last_proc_id ? _GEN_1114 : _GEN_524; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1587 = 2'h1 != last_proc_id ? _GEN_1115 : _GEN_525; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1588 = 2'h1 != last_proc_id ? _GEN_1116 : _GEN_526; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1589 = 2'h1 != last_proc_id ? _GEN_1117 : _GEN_527; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1590 = 2'h1 != last_proc_id ? _GEN_1118 : _GEN_528; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1591 = 2'h1 != last_proc_id ? _GEN_1119 : _GEN_529; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1592 = 2'h1 != last_proc_id ? _GEN_1120 : _GEN_530; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1593 = 2'h1 != last_proc_id ? _GEN_1121 : _GEN_531; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1594 = 2'h1 != last_proc_id ? _GEN_1122 : _GEN_532; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1595 = 2'h1 != last_proc_id ? _GEN_1123 : _GEN_533; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1596 = 2'h1 != last_proc_id ? _GEN_1124 : _GEN_534; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1597 = 2'h1 != last_proc_id ? _GEN_1125 : _GEN_535; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1598 = 2'h1 != last_proc_id ? _GEN_1126 : _GEN_536; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1599 = 2'h1 != last_proc_id ? _GEN_1127 : _GEN_537; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1600 = 2'h1 != last_proc_id ? _GEN_1128 : _GEN_538; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1601 = 2'h1 != last_proc_id ? _GEN_1129 : _GEN_539; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1602 = 2'h1 != last_proc_id ? _GEN_1130 : _GEN_540; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1603 = 2'h1 != last_proc_id ? _GEN_1131 : _GEN_541; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1604 = 2'h1 != last_proc_id ? _GEN_1132 : _GEN_542; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1605 = 2'h1 != last_proc_id ? _GEN_1133 : _GEN_543; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1606 = 2'h1 != last_proc_id ? _GEN_1134 : _GEN_544; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1607 = 2'h1 != last_proc_id ? _GEN_1135 : _GEN_545; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1608 = 2'h1 != last_proc_id ? _GEN_1136 : _GEN_546; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1609 = 2'h1 != last_proc_id ? _GEN_1137 : _GEN_547; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1610 = 2'h1 != last_proc_id ? _GEN_1138 : _GEN_548; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1611 = 2'h1 != last_proc_id ? _GEN_1139 : _GEN_549; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1612 = 2'h1 != last_proc_id ? _GEN_1140 : _GEN_550; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1613 = 2'h1 != last_proc_id ? _GEN_1141 : _GEN_551; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1614 = 2'h1 != last_proc_id ? _GEN_1142 : _GEN_552; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1615 = 2'h1 != last_proc_id ? _GEN_1143 : _GEN_553; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1616 = 2'h1 != last_proc_id ? _GEN_1144 : _GEN_554; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1617 = 2'h1 != last_proc_id ? _GEN_1145 : _GEN_555; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1618 = 2'h1 != last_proc_id ? _GEN_1146 : _GEN_556; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1619 = 2'h1 != last_proc_id ? _GEN_1147 : _GEN_557; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1620 = 2'h1 != last_proc_id ? _GEN_1148 : _GEN_558; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1621 = 2'h1 != last_proc_id ? _GEN_1149 : _GEN_559; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1622 = 2'h1 != last_proc_id ? _GEN_1150 : _GEN_560; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1623 = 2'h1 != last_proc_id ? _GEN_1151 : _GEN_561; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1624 = 2'h1 != last_proc_id ? _GEN_1152 : _GEN_562; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1625 = 2'h1 != last_proc_id ? _GEN_1153 : _GEN_563; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1626 = 2'h1 != last_proc_id ? _GEN_1154 : _GEN_564; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1627 = 2'h1 != last_proc_id ? _GEN_1155 : _GEN_565; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1628 = 2'h1 != last_proc_id ? _GEN_1156 : _GEN_566; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1629 = 2'h1 != last_proc_id ? _GEN_1157 : _GEN_567; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1630 = 2'h1 != last_proc_id ? _GEN_1158 : _GEN_568; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1631 = 2'h1 != last_proc_id ? _GEN_1159 : _GEN_569; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1632 = 2'h1 != last_proc_id ? _GEN_1160 : _GEN_570; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1633 = 2'h1 != last_proc_id ? _GEN_1161 : _GEN_571; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1634 = 2'h1 != last_proc_id ? _GEN_1162 : _GEN_572; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1635 = 2'h1 != last_proc_id ? _GEN_1163 : _GEN_573; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1636 = 2'h1 != last_proc_id ? _GEN_1164 : _GEN_574; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1637 = 2'h1 != last_proc_id ? _GEN_1165 : _GEN_575; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1638 = 2'h1 != last_proc_id ? _GEN_1166 : _GEN_576; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1639 = 2'h1 != last_proc_id ? _GEN_1167 : _GEN_577; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1640 = 2'h1 != last_proc_id ? _GEN_1168 : _GEN_578; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1641 = 2'h1 != last_proc_id ? _GEN_1169 : _GEN_579; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1642 = 2'h1 != last_proc_id ? _GEN_1170 : _GEN_580; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1643 = 2'h1 != last_proc_id ? _GEN_1171 : _GEN_581; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1644 = 2'h1 != last_proc_id ? _GEN_1172 : _GEN_582; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1645 = 2'h1 != last_proc_id ? _GEN_1173 : _GEN_583; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1646 = 2'h1 != last_proc_id ? _GEN_1174 : _GEN_584; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1647 = 2'h1 != last_proc_id ? _GEN_1175 : _GEN_585; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1648 = 2'h1 != last_proc_id ? _GEN_1176 : _GEN_586; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1649 = 2'h1 != last_proc_id ? _GEN_1177 : _GEN_587; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1650 = 2'h1 != last_proc_id ? _GEN_1178 : _GEN_588; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1651 = 2'h1 != last_proc_id ? _GEN_1179 : _GEN_589; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1652 = 2'h1 != last_proc_id ? _GEN_1180 : _GEN_590; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1653 = 2'h1 != last_proc_id ? _GEN_1181 : _GEN_591; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1654 = 2'h1 != last_proc_id ? _GEN_1182 : _GEN_592; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1655 = 2'h1 != last_proc_id ? _GEN_1183 : _GEN_593; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1656 = 2'h1 != last_proc_id ? _GEN_1184 : _GEN_594; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1657 = 2'h1 != last_proc_id ? _GEN_1185 : _GEN_595; // @[ipsa.scala 94:65]
  wire  _GEN_1658 = 2'h1 != last_proc_id ? _GEN_1186 : _GEN_596; // @[ipsa.scala 94:65]
  wire  _GEN_1659 = 2'h1 != last_proc_id ? _GEN_1187 : _GEN_597; // @[ipsa.scala 94:65]
  wire [1:0] _GEN_1660 = 2'h1 != last_proc_id ? _GEN_1188 : _GEN_598; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1661 = 2'h1 != last_proc_id ? _GEN_1189 : _GEN_599; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1662 = 2'h1 != last_proc_id ? _GEN_1190 : _GEN_600; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1663 = 2'h1 != last_proc_id ? _GEN_1191 : _GEN_601; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1664 = 2'h1 != last_proc_id ? _GEN_1192 : _GEN_602; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1665 = 2'h1 != last_proc_id ? _GEN_1193 : _GEN_603; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1666 = 2'h1 != last_proc_id ? _GEN_1194 : _GEN_604; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1667 = 2'h1 != last_proc_id ? _GEN_1195 : _GEN_605; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1668 = 2'h1 != last_proc_id ? _GEN_1196 : _GEN_606; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1669 = 2'h1 != last_proc_id ? _GEN_1197 : _GEN_607; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1670 = 2'h1 != last_proc_id ? _GEN_1198 : _GEN_608; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1671 = 2'h1 != last_proc_id ? _GEN_1199 : _GEN_609; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1672 = 2'h1 != last_proc_id ? _GEN_1200 : _GEN_610; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1673 = 2'h1 != last_proc_id ? _GEN_1201 : _GEN_611; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1674 = 2'h1 != last_proc_id ? _GEN_1202 : _GEN_612; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1675 = 2'h1 != last_proc_id ? _GEN_1203 : _GEN_613; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1676 = 2'h1 != last_proc_id ? _GEN_1204 : _GEN_614; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1677 = 2'h1 != last_proc_id ? _GEN_1205 : _GEN_615; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1678 = 2'h1 != last_proc_id ? _GEN_1206 : _GEN_616; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1679 = 2'h1 != last_proc_id ? _GEN_1207 : _GEN_617; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1680 = 2'h1 != last_proc_id ? _GEN_1208 : _GEN_618; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1681 = 2'h1 != last_proc_id ? _GEN_1209 : _GEN_619; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1682 = 2'h1 != last_proc_id ? _GEN_1210 : _GEN_620; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1683 = 2'h1 != last_proc_id ? _GEN_1211 : _GEN_621; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1684 = 2'h1 != last_proc_id ? _GEN_1212 : _GEN_622; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1685 = 2'h1 != last_proc_id ? _GEN_1213 : _GEN_623; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1686 = 2'h1 != last_proc_id ? _GEN_1214 : _GEN_624; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1687 = 2'h1 != last_proc_id ? _GEN_1215 : _GEN_625; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1688 = 2'h1 != last_proc_id ? _GEN_1216 : _GEN_626; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1689 = 2'h1 != last_proc_id ? _GEN_1217 : _GEN_627; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1690 = 2'h1 != last_proc_id ? _GEN_1218 : _GEN_628; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1691 = 2'h1 != last_proc_id ? _GEN_1219 : _GEN_629; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1692 = 2'h1 != last_proc_id ? _GEN_1220 : _GEN_630; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1693 = 2'h1 != last_proc_id ? _GEN_1221 : _GEN_631; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1694 = 2'h1 != last_proc_id ? _GEN_1222 : _GEN_632; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1695 = 2'h1 != last_proc_id ? _GEN_1223 : _GEN_633; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1696 = 2'h1 != last_proc_id ? _GEN_1224 : _GEN_634; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1697 = 2'h1 != last_proc_id ? _GEN_1225 : _GEN_635; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1698 = 2'h1 != last_proc_id ? _GEN_1226 : _GEN_636; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1699 = 2'h1 != last_proc_id ? _GEN_1227 : _GEN_637; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1700 = 2'h1 != last_proc_id ? _GEN_1228 : _GEN_638; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1701 = 2'h1 != last_proc_id ? _GEN_1229 : _GEN_639; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1702 = 2'h1 != last_proc_id ? _GEN_1230 : _GEN_640; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1703 = 2'h1 != last_proc_id ? _GEN_1231 : _GEN_641; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1704 = 2'h1 != last_proc_id ? _GEN_1232 : _GEN_642; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1705 = 2'h1 != last_proc_id ? _GEN_1233 : _GEN_643; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1706 = 2'h1 != last_proc_id ? _GEN_1234 : _GEN_644; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1707 = 2'h1 != last_proc_id ? _GEN_1235 : _GEN_645; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1708 = 2'h1 != last_proc_id ? _GEN_1236 : _GEN_646; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1709 = 2'h1 != last_proc_id ? _GEN_1237 : _GEN_647; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1710 = 2'h1 != last_proc_id ? _GEN_1238 : _GEN_648; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1711 = 2'h1 != last_proc_id ? _GEN_1239 : _GEN_649; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1712 = 2'h1 != last_proc_id ? _GEN_1240 : _GEN_650; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1713 = 2'h1 != last_proc_id ? _GEN_1241 : _GEN_651; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1714 = 2'h1 != last_proc_id ? _GEN_1242 : _GEN_652; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1715 = 2'h1 != last_proc_id ? _GEN_1243 : _GEN_653; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1716 = 2'h1 != last_proc_id ? _GEN_1244 : _GEN_654; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1717 = 2'h1 != last_proc_id ? _GEN_1245 : _GEN_655; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1718 = 2'h1 != last_proc_id ? _GEN_1246 : _GEN_656; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1719 = 2'h1 != last_proc_id ? _GEN_1247 : _GEN_657; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1720 = 2'h1 != last_proc_id ? _GEN_1248 : _GEN_658; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1721 = 2'h1 != last_proc_id ? _GEN_1249 : _GEN_659; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1722 = 2'h1 != last_proc_id ? _GEN_1250 : _GEN_660; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1723 = 2'h1 != last_proc_id ? _GEN_1251 : _GEN_661; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1724 = 2'h1 != last_proc_id ? _GEN_1252 : _GEN_662; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1725 = 2'h1 != last_proc_id ? _GEN_1253 : _GEN_663; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1726 = 2'h1 != last_proc_id ? _GEN_1254 : _GEN_664; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1727 = 2'h1 != last_proc_id ? _GEN_1255 : _GEN_665; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1728 = 2'h1 != last_proc_id ? _GEN_1256 : _GEN_666; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1729 = 2'h1 != last_proc_id ? _GEN_1257 : _GEN_667; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1730 = 2'h1 != last_proc_id ? _GEN_1258 : _GEN_668; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1731 = 2'h1 != last_proc_id ? _GEN_1259 : _GEN_669; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1732 = 2'h1 != last_proc_id ? _GEN_1260 : _GEN_670; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1733 = 2'h1 != last_proc_id ? _GEN_1261 : _GEN_671; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1734 = 2'h1 != last_proc_id ? _GEN_1262 : _GEN_672; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1735 = 2'h1 != last_proc_id ? _GEN_1263 : _GEN_673; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1736 = 2'h1 != last_proc_id ? _GEN_1264 : _GEN_674; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1737 = 2'h1 != last_proc_id ? _GEN_1265 : _GEN_675; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1738 = 2'h1 != last_proc_id ? _GEN_1266 : _GEN_676; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1739 = 2'h1 != last_proc_id ? _GEN_1267 : _GEN_677; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1740 = 2'h1 != last_proc_id ? _GEN_1268 : _GEN_678; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1741 = 2'h1 != last_proc_id ? _GEN_1269 : _GEN_679; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1742 = 2'h1 != last_proc_id ? _GEN_1270 : _GEN_680; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1743 = 2'h1 != last_proc_id ? _GEN_1271 : _GEN_681; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1744 = 2'h1 != last_proc_id ? _GEN_1272 : _GEN_682; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1745 = 2'h1 != last_proc_id ? _GEN_1273 : _GEN_683; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1746 = 2'h1 != last_proc_id ? _GEN_1274 : _GEN_684; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1747 = 2'h1 != last_proc_id ? _GEN_1275 : _GEN_685; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1748 = 2'h1 != last_proc_id ? _GEN_1276 : _GEN_686; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1749 = 2'h1 != last_proc_id ? _GEN_1277 : _GEN_687; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1750 = 2'h1 != last_proc_id ? _GEN_1278 : _GEN_688; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1751 = 2'h1 != last_proc_id ? _GEN_1279 : _GEN_689; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1752 = 2'h1 != last_proc_id ? _GEN_1280 : _GEN_690; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1753 = 2'h1 != last_proc_id ? _GEN_1281 : _GEN_691; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1754 = 2'h1 != last_proc_id ? _GEN_1282 : _GEN_692; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1755 = 2'h1 != last_proc_id ? _GEN_1283 : _GEN_693; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1756 = 2'h1 != last_proc_id ? _GEN_1284 : _GEN_694; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1757 = 2'h1 != last_proc_id ? _GEN_1285 : _GEN_695; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1758 = 2'h1 != last_proc_id ? _GEN_1286 : _GEN_696; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1759 = 2'h1 != last_proc_id ? _GEN_1287 : _GEN_697; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1760 = 2'h1 != last_proc_id ? _GEN_1288 : _GEN_698; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1761 = 2'h1 != last_proc_id ? _GEN_1289 : _GEN_699; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1762 = 2'h1 != last_proc_id ? _GEN_1290 : _GEN_700; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1763 = 2'h1 != last_proc_id ? _GEN_1291 : _GEN_701; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1764 = 2'h1 != last_proc_id ? _GEN_1292 : _GEN_702; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1765 = 2'h1 != last_proc_id ? _GEN_1293 : _GEN_703; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1766 = 2'h1 != last_proc_id ? _GEN_1294 : _GEN_704; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1767 = 2'h1 != last_proc_id ? _GEN_1295 : _GEN_705; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1768 = 2'h1 != last_proc_id ? _GEN_1296 : _GEN_706; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1769 = 2'h1 != last_proc_id ? _GEN_1297 : _GEN_707; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1770 = 2'h1 != last_proc_id ? _GEN_1298 : _GEN_708; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1771 = 2'h1 != last_proc_id ? _GEN_1299 : _GEN_709; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1772 = 2'h1 != last_proc_id ? _GEN_1300 : _GEN_710; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1773 = 2'h1 != last_proc_id ? _GEN_1301 : _GEN_711; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1774 = 2'h1 != last_proc_id ? _GEN_1302 : _GEN_712; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1775 = 2'h1 != last_proc_id ? _GEN_1303 : _GEN_713; // @[ipsa.scala 94:65]
  wire  _GEN_1776 = 2'h1 != last_proc_id ? _GEN_1304 : _GEN_714; // @[ipsa.scala 94:65]
  wire  _GEN_1777 = 2'h1 != last_proc_id ? _GEN_1305 : _GEN_715; // @[ipsa.scala 94:65]
  wire [1:0] _GEN_1778 = 2'h1 != last_proc_id ? _GEN_1306 : _GEN_716; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1779 = 2'h1 != last_proc_id ? _GEN_1307 : _GEN_717; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1780 = 2'h1 != last_proc_id ? _GEN_1308 : _GEN_718; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1781 = 2'h1 != last_proc_id ? _GEN_1309 : _GEN_719; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1782 = 2'h1 != last_proc_id ? _GEN_1310 : _GEN_720; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1783 = 2'h1 != last_proc_id ? _GEN_1311 : _GEN_721; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1784 = 2'h1 != last_proc_id ? _GEN_1312 : _GEN_722; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1785 = 2'h1 != last_proc_id ? _GEN_1313 : _GEN_723; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1786 = 2'h1 != last_proc_id ? _GEN_1314 : _GEN_724; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1787 = 2'h1 != last_proc_id ? _GEN_1315 : _GEN_725; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1788 = 2'h1 != last_proc_id ? _GEN_1316 : _GEN_726; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1789 = 2'h1 != last_proc_id ? _GEN_1317 : _GEN_727; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1790 = 2'h1 != last_proc_id ? _GEN_1318 : _GEN_728; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1791 = 2'h1 != last_proc_id ? _GEN_1319 : _GEN_729; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1792 = 2'h1 != last_proc_id ? _GEN_1320 : _GEN_730; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1793 = 2'h1 != last_proc_id ? _GEN_1321 : _GEN_731; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1794 = 2'h1 != last_proc_id ? _GEN_1322 : _GEN_732; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1795 = 2'h1 != last_proc_id ? _GEN_1323 : _GEN_733; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1796 = 2'h1 != last_proc_id ? _GEN_1324 : _GEN_734; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1797 = 2'h1 != last_proc_id ? _GEN_1325 : _GEN_735; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1798 = 2'h1 != last_proc_id ? _GEN_1326 : _GEN_736; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1799 = 2'h1 != last_proc_id ? _GEN_1327 : _GEN_737; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1800 = 2'h1 != last_proc_id ? _GEN_1328 : _GEN_738; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1801 = 2'h1 != last_proc_id ? _GEN_1329 : _GEN_739; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1802 = 2'h1 != last_proc_id ? _GEN_1330 : _GEN_740; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1803 = 2'h1 != last_proc_id ? _GEN_1331 : _GEN_741; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1804 = 2'h1 != last_proc_id ? _GEN_1332 : _GEN_742; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1805 = 2'h1 != last_proc_id ? _GEN_1333 : _GEN_743; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1806 = 2'h1 != last_proc_id ? _GEN_1334 : _GEN_744; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1807 = 2'h1 != last_proc_id ? _GEN_1335 : _GEN_745; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1808 = 2'h1 != last_proc_id ? _GEN_1336 : _GEN_746; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1809 = 2'h1 != last_proc_id ? _GEN_1337 : _GEN_747; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1810 = 2'h1 != last_proc_id ? _GEN_1338 : _GEN_748; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1811 = 2'h1 != last_proc_id ? _GEN_1339 : _GEN_749; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1812 = 2'h1 != last_proc_id ? _GEN_1340 : _GEN_750; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1813 = 2'h1 != last_proc_id ? _GEN_1341 : _GEN_751; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1814 = 2'h1 != last_proc_id ? _GEN_1342 : _GEN_752; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1815 = 2'h1 != last_proc_id ? _GEN_1343 : _GEN_753; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1816 = 2'h1 != last_proc_id ? _GEN_1344 : _GEN_754; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1817 = 2'h1 != last_proc_id ? _GEN_1345 : _GEN_755; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1818 = 2'h1 != last_proc_id ? _GEN_1346 : _GEN_756; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1819 = 2'h1 != last_proc_id ? _GEN_1347 : _GEN_757; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1820 = 2'h1 != last_proc_id ? _GEN_1348 : _GEN_758; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1821 = 2'h1 != last_proc_id ? _GEN_1349 : _GEN_759; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1822 = 2'h1 != last_proc_id ? _GEN_1350 : _GEN_760; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1823 = 2'h1 != last_proc_id ? _GEN_1351 : _GEN_761; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1824 = 2'h1 != last_proc_id ? _GEN_1352 : _GEN_762; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1825 = 2'h1 != last_proc_id ? _GEN_1353 : _GEN_763; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1826 = 2'h1 != last_proc_id ? _GEN_1354 : _GEN_764; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1827 = 2'h1 != last_proc_id ? _GEN_1355 : _GEN_765; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1828 = 2'h1 != last_proc_id ? _GEN_1356 : _GEN_766; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1829 = 2'h1 != last_proc_id ? _GEN_1357 : _GEN_767; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1830 = 2'h1 != last_proc_id ? _GEN_1358 : _GEN_768; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1831 = 2'h1 != last_proc_id ? _GEN_1359 : _GEN_769; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1832 = 2'h1 != last_proc_id ? _GEN_1360 : _GEN_770; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1833 = 2'h1 != last_proc_id ? _GEN_1361 : _GEN_771; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1834 = 2'h1 != last_proc_id ? _GEN_1362 : _GEN_772; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1835 = 2'h1 != last_proc_id ? _GEN_1363 : _GEN_773; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1836 = 2'h1 != last_proc_id ? _GEN_1364 : _GEN_774; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1837 = 2'h1 != last_proc_id ? _GEN_1365 : _GEN_775; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1838 = 2'h1 != last_proc_id ? _GEN_1366 : _GEN_776; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1839 = 2'h1 != last_proc_id ? _GEN_1367 : _GEN_777; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1840 = 2'h1 != last_proc_id ? _GEN_1368 : _GEN_778; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1841 = 2'h1 != last_proc_id ? _GEN_1369 : _GEN_779; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1842 = 2'h1 != last_proc_id ? _GEN_1370 : _GEN_780; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1843 = 2'h1 != last_proc_id ? _GEN_1371 : _GEN_781; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1844 = 2'h1 != last_proc_id ? _GEN_1372 : _GEN_782; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1845 = 2'h1 != last_proc_id ? _GEN_1373 : _GEN_783; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1846 = 2'h1 != last_proc_id ? _GEN_1374 : _GEN_784; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1847 = 2'h1 != last_proc_id ? _GEN_1375 : _GEN_785; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1848 = 2'h1 != last_proc_id ? _GEN_1376 : _GEN_786; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1849 = 2'h1 != last_proc_id ? _GEN_1377 : _GEN_787; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1850 = 2'h1 != last_proc_id ? _GEN_1378 : _GEN_788; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1851 = 2'h1 != last_proc_id ? _GEN_1379 : _GEN_789; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1852 = 2'h1 != last_proc_id ? _GEN_1380 : _GEN_790; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1853 = 2'h1 != last_proc_id ? _GEN_1381 : _GEN_791; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1854 = 2'h1 != last_proc_id ? _GEN_1382 : _GEN_792; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1855 = 2'h1 != last_proc_id ? _GEN_1383 : _GEN_793; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1856 = 2'h1 != last_proc_id ? _GEN_1384 : _GEN_794; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1857 = 2'h1 != last_proc_id ? _GEN_1385 : _GEN_795; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1858 = 2'h1 != last_proc_id ? _GEN_1386 : _GEN_796; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1859 = 2'h1 != last_proc_id ? _GEN_1387 : _GEN_797; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1860 = 2'h1 != last_proc_id ? _GEN_1388 : _GEN_798; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1861 = 2'h1 != last_proc_id ? _GEN_1389 : _GEN_799; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1862 = 2'h1 != last_proc_id ? _GEN_1390 : _GEN_800; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1863 = 2'h1 != last_proc_id ? _GEN_1391 : _GEN_801; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1864 = 2'h1 != last_proc_id ? _GEN_1392 : _GEN_802; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1865 = 2'h1 != last_proc_id ? _GEN_1393 : _GEN_803; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1866 = 2'h1 != last_proc_id ? _GEN_1394 : _GEN_804; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1867 = 2'h1 != last_proc_id ? _GEN_1395 : _GEN_805; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1868 = 2'h1 != last_proc_id ? _GEN_1396 : _GEN_806; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1869 = 2'h1 != last_proc_id ? _GEN_1397 : _GEN_807; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1870 = 2'h1 != last_proc_id ? _GEN_1398 : _GEN_808; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1871 = 2'h1 != last_proc_id ? _GEN_1399 : _GEN_809; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1872 = 2'h1 != last_proc_id ? _GEN_1400 : _GEN_810; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1873 = 2'h1 != last_proc_id ? _GEN_1401 : _GEN_811; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1874 = 2'h1 != last_proc_id ? _GEN_1402 : _GEN_812; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1875 = 2'h1 != last_proc_id ? _GEN_1403 : _GEN_813; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1876 = 2'h1 != last_proc_id ? _GEN_1404 : _GEN_814; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1877 = 2'h1 != last_proc_id ? _GEN_1405 : _GEN_815; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1878 = 2'h1 != last_proc_id ? _GEN_1406 : _GEN_816; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1879 = 2'h1 != last_proc_id ? _GEN_1407 : _GEN_817; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1880 = 2'h1 != last_proc_id ? _GEN_1408 : _GEN_818; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1881 = 2'h1 != last_proc_id ? _GEN_1409 : _GEN_819; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1882 = 2'h1 != last_proc_id ? _GEN_1410 : _GEN_820; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1883 = 2'h1 != last_proc_id ? _GEN_1411 : _GEN_821; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1884 = 2'h1 != last_proc_id ? _GEN_1412 : _GEN_822; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1885 = 2'h1 != last_proc_id ? _GEN_1413 : _GEN_823; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1886 = 2'h1 != last_proc_id ? _GEN_1414 : _GEN_824; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1887 = 2'h1 != last_proc_id ? _GEN_1415 : _GEN_825; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1888 = 2'h1 != last_proc_id ? _GEN_1416 : _GEN_826; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1889 = 2'h1 != last_proc_id ? _GEN_1417 : _GEN_827; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1890 = 2'h1 != last_proc_id ? _GEN_1418 : _GEN_828; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1891 = 2'h1 != last_proc_id ? _GEN_1419 : _GEN_829; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1892 = 2'h1 != last_proc_id ? _GEN_1420 : _GEN_830; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1893 = 2'h1 != last_proc_id ? _GEN_1421 : _GEN_831; // @[ipsa.scala 94:65]
  wire  _GEN_1894 = 2'h1 != last_proc_id ? _GEN_1422 : _GEN_832; // @[ipsa.scala 94:65]
  wire  _GEN_1895 = 2'h1 != last_proc_id ? _GEN_1423 : _GEN_833; // @[ipsa.scala 94:65]
  wire [1:0] _GEN_1896 = 2'h1 != last_proc_id ? _GEN_1424 : _GEN_834; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1897 = 2'h1 != last_proc_id ? _GEN_1425 : _GEN_835; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1898 = 2'h1 != last_proc_id ? _GEN_1426 : _GEN_836; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1899 = 2'h1 != last_proc_id ? _GEN_1427 : _GEN_837; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1900 = 2'h1 != last_proc_id ? _GEN_1428 : _GEN_838; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1901 = 2'h1 != last_proc_id ? _GEN_1429 : _GEN_839; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1902 = 2'h1 != last_proc_id ? _GEN_1430 : _GEN_840; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1903 = 2'h1 != last_proc_id ? _GEN_1431 : _GEN_841; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1904 = 2'h1 != last_proc_id ? _GEN_1432 : _GEN_842; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1905 = 2'h1 != last_proc_id ? _GEN_1433 : _GEN_843; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1906 = 2'h1 != last_proc_id ? _GEN_1434 : _GEN_844; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1907 = 2'h1 != last_proc_id ? _GEN_1435 : _GEN_845; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1908 = 2'h1 != last_proc_id ? _GEN_1436 : _GEN_846; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1909 = 2'h1 != last_proc_id ? _GEN_1437 : _GEN_847; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1910 = 2'h1 != last_proc_id ? _GEN_1438 : _GEN_848; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1911 = 2'h1 != last_proc_id ? _GEN_1439 : _GEN_849; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1912 = 2'h1 != last_proc_id ? _GEN_1440 : _GEN_850; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1913 = 2'h1 != last_proc_id ? _GEN_1441 : _GEN_851; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1914 = 2'h1 != last_proc_id ? _GEN_1442 : _GEN_852; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_1915 = 2'h1 != last_proc_id ? _GEN_1443 : _GEN_853; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1916 = 2'h1 != last_proc_id ? _GEN_1444 : _GEN_854; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1917 = 2'h1 != last_proc_id ? _GEN_1445 : _GEN_855; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1918 = 2'h1 != last_proc_id ? _GEN_1446 : _GEN_856; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1919 = 2'h1 != last_proc_id ? _GEN_1447 : _GEN_857; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1920 = 2'h1 != last_proc_id ? _GEN_1448 : _GEN_858; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1921 = 2'h1 != last_proc_id ? _GEN_1449 : _GEN_859; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1922 = 2'h1 != last_proc_id ? _GEN_1450 : _GEN_860; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1923 = 2'h1 != last_proc_id ? _GEN_1451 : _GEN_861; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1924 = 2'h1 != last_proc_id ? _GEN_1452 : _GEN_862; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1925 = 2'h1 != last_proc_id ? _GEN_1453 : _GEN_863; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1926 = 2'h1 != last_proc_id ? _GEN_1454 : _GEN_864; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1927 = 2'h1 != last_proc_id ? _GEN_1455 : _GEN_865; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1928 = 2'h1 != last_proc_id ? _GEN_1456 : _GEN_866; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1929 = 2'h1 != last_proc_id ? _GEN_1457 : _GEN_867; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1930 = 2'h1 != last_proc_id ? _GEN_1458 : _GEN_868; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1931 = 2'h1 != last_proc_id ? _GEN_1459 : _GEN_869; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1932 = 2'h1 != last_proc_id ? _GEN_1460 : _GEN_870; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1933 = 2'h1 != last_proc_id ? _GEN_1461 : _GEN_871; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1934 = 2'h1 != last_proc_id ? _GEN_1462 : _GEN_872; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1935 = 2'h1 != last_proc_id ? _GEN_1463 : _GEN_873; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1936 = 2'h1 != last_proc_id ? _GEN_1464 : _GEN_874; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1937 = 2'h1 != last_proc_id ? _GEN_1465 : _GEN_875; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1938 = 2'h1 != last_proc_id ? _GEN_1466 : _GEN_876; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1939 = 2'h1 != last_proc_id ? _GEN_1467 : _GEN_877; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1940 = 2'h1 != last_proc_id ? _GEN_1468 : _GEN_878; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1941 = 2'h1 != last_proc_id ? _GEN_1469 : _GEN_879; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1942 = 2'h1 != last_proc_id ? _GEN_1470 : _GEN_880; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1943 = 2'h1 != last_proc_id ? _GEN_1471 : _GEN_881; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1944 = 2'h1 != last_proc_id ? _GEN_1472 : _GEN_882; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1945 = 2'h1 != last_proc_id ? _GEN_1473 : _GEN_883; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1946 = 2'h1 != last_proc_id ? _GEN_1474 : _GEN_884; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1947 = 2'h1 != last_proc_id ? _GEN_1475 : _GEN_885; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1948 = 2'h1 != last_proc_id ? _GEN_1476 : _GEN_886; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1949 = 2'h1 != last_proc_id ? _GEN_1477 : _GEN_887; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1950 = 2'h1 != last_proc_id ? _GEN_1478 : _GEN_888; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1951 = 2'h1 != last_proc_id ? _GEN_1479 : _GEN_889; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1952 = 2'h1 != last_proc_id ? _GEN_1480 : _GEN_890; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1953 = 2'h1 != last_proc_id ? _GEN_1481 : _GEN_891; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1954 = 2'h1 != last_proc_id ? _GEN_1482 : _GEN_892; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1955 = 2'h1 != last_proc_id ? _GEN_1483 : _GEN_893; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1956 = 2'h1 != last_proc_id ? _GEN_1484 : _GEN_894; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1957 = 2'h1 != last_proc_id ? _GEN_1485 : _GEN_895; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1958 = 2'h1 != last_proc_id ? _GEN_1486 : _GEN_896; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1959 = 2'h1 != last_proc_id ? _GEN_1487 : _GEN_897; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1960 = 2'h1 != last_proc_id ? _GEN_1488 : _GEN_898; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1961 = 2'h1 != last_proc_id ? _GEN_1489 : _GEN_899; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1962 = 2'h1 != last_proc_id ? _GEN_1490 : _GEN_900; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1963 = 2'h1 != last_proc_id ? _GEN_1491 : _GEN_901; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1964 = 2'h1 != last_proc_id ? _GEN_1492 : _GEN_902; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1965 = 2'h1 != last_proc_id ? _GEN_1493 : _GEN_903; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1966 = 2'h1 != last_proc_id ? _GEN_1494 : _GEN_904; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1967 = 2'h1 != last_proc_id ? _GEN_1495 : _GEN_905; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1968 = 2'h1 != last_proc_id ? _GEN_1496 : _GEN_906; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1969 = 2'h1 != last_proc_id ? _GEN_1497 : _GEN_907; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1970 = 2'h1 != last_proc_id ? _GEN_1498 : _GEN_908; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1971 = 2'h1 != last_proc_id ? _GEN_1499 : _GEN_909; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1972 = 2'h1 != last_proc_id ? _GEN_1500 : _GEN_910; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1973 = 2'h1 != last_proc_id ? _GEN_1501 : _GEN_911; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1974 = 2'h1 != last_proc_id ? _GEN_1502 : _GEN_912; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1975 = 2'h1 != last_proc_id ? _GEN_1503 : _GEN_913; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1976 = 2'h1 != last_proc_id ? _GEN_1504 : _GEN_914; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1977 = 2'h1 != last_proc_id ? _GEN_1505 : _GEN_915; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1978 = 2'h1 != last_proc_id ? _GEN_1506 : _GEN_916; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1979 = 2'h1 != last_proc_id ? _GEN_1507 : _GEN_917; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1980 = 2'h1 != last_proc_id ? _GEN_1508 : _GEN_918; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1981 = 2'h1 != last_proc_id ? _GEN_1509 : _GEN_919; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1982 = 2'h1 != last_proc_id ? _GEN_1510 : _GEN_920; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1983 = 2'h1 != last_proc_id ? _GEN_1511 : _GEN_921; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1984 = 2'h1 != last_proc_id ? _GEN_1512 : _GEN_922; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1985 = 2'h1 != last_proc_id ? _GEN_1513 : _GEN_923; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1986 = 2'h1 != last_proc_id ? _GEN_1514 : _GEN_924; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1987 = 2'h1 != last_proc_id ? _GEN_1515 : _GEN_925; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1988 = 2'h1 != last_proc_id ? _GEN_1516 : _GEN_926; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1989 = 2'h1 != last_proc_id ? _GEN_1517 : _GEN_927; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1990 = 2'h1 != last_proc_id ? _GEN_1518 : _GEN_928; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1991 = 2'h1 != last_proc_id ? _GEN_1519 : _GEN_929; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1992 = 2'h1 != last_proc_id ? _GEN_1520 : _GEN_930; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1993 = 2'h1 != last_proc_id ? _GEN_1521 : _GEN_931; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1994 = 2'h1 != last_proc_id ? _GEN_1522 : _GEN_932; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1995 = 2'h1 != last_proc_id ? _GEN_1523 : _GEN_933; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1996 = 2'h1 != last_proc_id ? _GEN_1524 : _GEN_934; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1997 = 2'h1 != last_proc_id ? _GEN_1525 : _GEN_935; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1998 = 2'h1 != last_proc_id ? _GEN_1526 : _GEN_936; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_1999 = 2'h1 != last_proc_id ? _GEN_1527 : _GEN_937; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2000 = 2'h1 != last_proc_id ? _GEN_1528 : _GEN_938; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2001 = 2'h1 != last_proc_id ? _GEN_1529 : _GEN_939; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2002 = 2'h1 != last_proc_id ? _GEN_1530 : _GEN_940; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2003 = 2'h1 != last_proc_id ? _GEN_1531 : _GEN_941; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2004 = 2'h1 != last_proc_id ? _GEN_1532 : _GEN_942; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2005 = 2'h1 != last_proc_id ? _GEN_1533 : _GEN_943; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2006 = 2'h1 != last_proc_id ? _GEN_1534 : _GEN_944; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2007 = 2'h1 != last_proc_id ? _GEN_1535 : _GEN_945; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2008 = 2'h1 != last_proc_id ? _GEN_1536 : _GEN_946; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2009 = 2'h1 != last_proc_id ? _GEN_1537 : _GEN_947; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2010 = 2'h1 != last_proc_id ? _GEN_1538 : _GEN_948; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2011 = 2'h1 != last_proc_id ? _GEN_1539 : _GEN_949; // @[ipsa.scala 94:65]
  wire  _GEN_2012 = 2'h1 != last_proc_id ? _GEN_950 : trans_1_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire  _GEN_2013 = 2'h1 != last_proc_id ? _GEN_951 : trans_1_io_pipe_phv_out_next_config_id; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [1:0] _GEN_2014 = 2'h1 != last_proc_id ? _GEN_952 : trans_1_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_2015 = 2'h1 != last_proc_id ? _GEN_953 : trans_1_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2016 = 2'h1 != last_proc_id ? _GEN_954 : trans_1_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2017 = 2'h1 != last_proc_id ? _GEN_955 : trans_1_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_2018 = 2'h1 != last_proc_id ? _GEN_956 : trans_1_io_pipe_phv_out_header_0; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_2019 = 2'h1 != last_proc_id ? _GEN_957 : trans_1_io_pipe_phv_out_header_1; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_2020 = 2'h1 != last_proc_id ? _GEN_958 : trans_1_io_pipe_phv_out_header_2; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_2021 = 2'h1 != last_proc_id ? _GEN_959 : trans_1_io_pipe_phv_out_header_3; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_2022 = 2'h1 != last_proc_id ? _GEN_960 : trans_1_io_pipe_phv_out_header_4; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_2023 = 2'h1 != last_proc_id ? _GEN_961 : trans_1_io_pipe_phv_out_header_5; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_2024 = 2'h1 != last_proc_id ? _GEN_962 : trans_1_io_pipe_phv_out_header_6; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_2025 = 2'h1 != last_proc_id ? _GEN_963 : trans_1_io_pipe_phv_out_header_7; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_2026 = 2'h1 != last_proc_id ? _GEN_964 : trans_1_io_pipe_phv_out_header_8; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_2027 = 2'h1 != last_proc_id ? _GEN_965 : trans_1_io_pipe_phv_out_header_9; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_2028 = 2'h1 != last_proc_id ? _GEN_966 : trans_1_io_pipe_phv_out_header_10; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_2029 = 2'h1 != last_proc_id ? _GEN_967 : trans_1_io_pipe_phv_out_header_11; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_2030 = 2'h1 != last_proc_id ? _GEN_968 : trans_1_io_pipe_phv_out_header_12; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_2031 = 2'h1 != last_proc_id ? _GEN_969 : trans_1_io_pipe_phv_out_header_13; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_2032 = 2'h1 != last_proc_id ? _GEN_970 : trans_1_io_pipe_phv_out_header_14; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_2033 = 2'h1 != last_proc_id ? _GEN_971 : trans_1_io_pipe_phv_out_header_15; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2034 = 2'h1 != last_proc_id ? _GEN_972 : trans_1_io_pipe_phv_out_data_0; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2035 = 2'h1 != last_proc_id ? _GEN_973 : trans_1_io_pipe_phv_out_data_1; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2036 = 2'h1 != last_proc_id ? _GEN_974 : trans_1_io_pipe_phv_out_data_2; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2037 = 2'h1 != last_proc_id ? _GEN_975 : trans_1_io_pipe_phv_out_data_3; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2038 = 2'h1 != last_proc_id ? _GEN_976 : trans_1_io_pipe_phv_out_data_4; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2039 = 2'h1 != last_proc_id ? _GEN_977 : trans_1_io_pipe_phv_out_data_5; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2040 = 2'h1 != last_proc_id ? _GEN_978 : trans_1_io_pipe_phv_out_data_6; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2041 = 2'h1 != last_proc_id ? _GEN_979 : trans_1_io_pipe_phv_out_data_7; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2042 = 2'h1 != last_proc_id ? _GEN_980 : trans_1_io_pipe_phv_out_data_8; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2043 = 2'h1 != last_proc_id ? _GEN_981 : trans_1_io_pipe_phv_out_data_9; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2044 = 2'h1 != last_proc_id ? _GEN_982 : trans_1_io_pipe_phv_out_data_10; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2045 = 2'h1 != last_proc_id ? _GEN_983 : trans_1_io_pipe_phv_out_data_11; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2046 = 2'h1 != last_proc_id ? _GEN_984 : trans_1_io_pipe_phv_out_data_12; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2047 = 2'h1 != last_proc_id ? _GEN_985 : trans_1_io_pipe_phv_out_data_13; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2048 = 2'h1 != last_proc_id ? _GEN_986 : trans_1_io_pipe_phv_out_data_14; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2049 = 2'h1 != last_proc_id ? _GEN_987 : trans_1_io_pipe_phv_out_data_15; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2050 = 2'h1 != last_proc_id ? _GEN_988 : trans_1_io_pipe_phv_out_data_16; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2051 = 2'h1 != last_proc_id ? _GEN_989 : trans_1_io_pipe_phv_out_data_17; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2052 = 2'h1 != last_proc_id ? _GEN_990 : trans_1_io_pipe_phv_out_data_18; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2053 = 2'h1 != last_proc_id ? _GEN_991 : trans_1_io_pipe_phv_out_data_19; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2054 = 2'h1 != last_proc_id ? _GEN_992 : trans_1_io_pipe_phv_out_data_20; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2055 = 2'h1 != last_proc_id ? _GEN_993 : trans_1_io_pipe_phv_out_data_21; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2056 = 2'h1 != last_proc_id ? _GEN_994 : trans_1_io_pipe_phv_out_data_22; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2057 = 2'h1 != last_proc_id ? _GEN_995 : trans_1_io_pipe_phv_out_data_23; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2058 = 2'h1 != last_proc_id ? _GEN_996 : trans_1_io_pipe_phv_out_data_24; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2059 = 2'h1 != last_proc_id ? _GEN_997 : trans_1_io_pipe_phv_out_data_25; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2060 = 2'h1 != last_proc_id ? _GEN_998 : trans_1_io_pipe_phv_out_data_26; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2061 = 2'h1 != last_proc_id ? _GEN_999 : trans_1_io_pipe_phv_out_data_27; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2062 = 2'h1 != last_proc_id ? _GEN_1000 : trans_1_io_pipe_phv_out_data_28; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2063 = 2'h1 != last_proc_id ? _GEN_1001 : trans_1_io_pipe_phv_out_data_29; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2064 = 2'h1 != last_proc_id ? _GEN_1002 : trans_1_io_pipe_phv_out_data_30; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2065 = 2'h1 != last_proc_id ? _GEN_1003 : trans_1_io_pipe_phv_out_data_31; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2066 = 2'h1 != last_proc_id ? _GEN_1004 : trans_1_io_pipe_phv_out_data_32; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2067 = 2'h1 != last_proc_id ? _GEN_1005 : trans_1_io_pipe_phv_out_data_33; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2068 = 2'h1 != last_proc_id ? _GEN_1006 : trans_1_io_pipe_phv_out_data_34; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2069 = 2'h1 != last_proc_id ? _GEN_1007 : trans_1_io_pipe_phv_out_data_35; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2070 = 2'h1 != last_proc_id ? _GEN_1008 : trans_1_io_pipe_phv_out_data_36; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2071 = 2'h1 != last_proc_id ? _GEN_1009 : trans_1_io_pipe_phv_out_data_37; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2072 = 2'h1 != last_proc_id ? _GEN_1010 : trans_1_io_pipe_phv_out_data_38; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2073 = 2'h1 != last_proc_id ? _GEN_1011 : trans_1_io_pipe_phv_out_data_39; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2074 = 2'h1 != last_proc_id ? _GEN_1012 : trans_1_io_pipe_phv_out_data_40; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2075 = 2'h1 != last_proc_id ? _GEN_1013 : trans_1_io_pipe_phv_out_data_41; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2076 = 2'h1 != last_proc_id ? _GEN_1014 : trans_1_io_pipe_phv_out_data_42; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2077 = 2'h1 != last_proc_id ? _GEN_1015 : trans_1_io_pipe_phv_out_data_43; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2078 = 2'h1 != last_proc_id ? _GEN_1016 : trans_1_io_pipe_phv_out_data_44; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2079 = 2'h1 != last_proc_id ? _GEN_1017 : trans_1_io_pipe_phv_out_data_45; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2080 = 2'h1 != last_proc_id ? _GEN_1018 : trans_1_io_pipe_phv_out_data_46; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2081 = 2'h1 != last_proc_id ? _GEN_1019 : trans_1_io_pipe_phv_out_data_47; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2082 = 2'h1 != last_proc_id ? _GEN_1020 : trans_1_io_pipe_phv_out_data_48; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2083 = 2'h1 != last_proc_id ? _GEN_1021 : trans_1_io_pipe_phv_out_data_49; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2084 = 2'h1 != last_proc_id ? _GEN_1022 : trans_1_io_pipe_phv_out_data_50; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2085 = 2'h1 != last_proc_id ? _GEN_1023 : trans_1_io_pipe_phv_out_data_51; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2086 = 2'h1 != last_proc_id ? _GEN_1024 : trans_1_io_pipe_phv_out_data_52; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2087 = 2'h1 != last_proc_id ? _GEN_1025 : trans_1_io_pipe_phv_out_data_53; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2088 = 2'h1 != last_proc_id ? _GEN_1026 : trans_1_io_pipe_phv_out_data_54; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2089 = 2'h1 != last_proc_id ? _GEN_1027 : trans_1_io_pipe_phv_out_data_55; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2090 = 2'h1 != last_proc_id ? _GEN_1028 : trans_1_io_pipe_phv_out_data_56; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2091 = 2'h1 != last_proc_id ? _GEN_1029 : trans_1_io_pipe_phv_out_data_57; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2092 = 2'h1 != last_proc_id ? _GEN_1030 : trans_1_io_pipe_phv_out_data_58; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2093 = 2'h1 != last_proc_id ? _GEN_1031 : trans_1_io_pipe_phv_out_data_59; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2094 = 2'h1 != last_proc_id ? _GEN_1032 : trans_1_io_pipe_phv_out_data_60; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2095 = 2'h1 != last_proc_id ? _GEN_1033 : trans_1_io_pipe_phv_out_data_61; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2096 = 2'h1 != last_proc_id ? _GEN_1034 : trans_1_io_pipe_phv_out_data_62; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2097 = 2'h1 != last_proc_id ? _GEN_1035 : trans_1_io_pipe_phv_out_data_63; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2098 = 2'h1 != last_proc_id ? _GEN_1036 : trans_1_io_pipe_phv_out_data_64; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2099 = 2'h1 != last_proc_id ? _GEN_1037 : trans_1_io_pipe_phv_out_data_65; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2100 = 2'h1 != last_proc_id ? _GEN_1038 : trans_1_io_pipe_phv_out_data_66; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2101 = 2'h1 != last_proc_id ? _GEN_1039 : trans_1_io_pipe_phv_out_data_67; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2102 = 2'h1 != last_proc_id ? _GEN_1040 : trans_1_io_pipe_phv_out_data_68; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2103 = 2'h1 != last_proc_id ? _GEN_1041 : trans_1_io_pipe_phv_out_data_69; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2104 = 2'h1 != last_proc_id ? _GEN_1042 : trans_1_io_pipe_phv_out_data_70; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2105 = 2'h1 != last_proc_id ? _GEN_1043 : trans_1_io_pipe_phv_out_data_71; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2106 = 2'h1 != last_proc_id ? _GEN_1044 : trans_1_io_pipe_phv_out_data_72; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2107 = 2'h1 != last_proc_id ? _GEN_1045 : trans_1_io_pipe_phv_out_data_73; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2108 = 2'h1 != last_proc_id ? _GEN_1046 : trans_1_io_pipe_phv_out_data_74; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2109 = 2'h1 != last_proc_id ? _GEN_1047 : trans_1_io_pipe_phv_out_data_75; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2110 = 2'h1 != last_proc_id ? _GEN_1048 : trans_1_io_pipe_phv_out_data_76; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2111 = 2'h1 != last_proc_id ? _GEN_1049 : trans_1_io_pipe_phv_out_data_77; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2112 = 2'h1 != last_proc_id ? _GEN_1050 : trans_1_io_pipe_phv_out_data_78; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2113 = 2'h1 != last_proc_id ? _GEN_1051 : trans_1_io_pipe_phv_out_data_79; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2114 = 2'h1 != last_proc_id ? _GEN_1052 : trans_1_io_pipe_phv_out_data_80; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2115 = 2'h1 != last_proc_id ? _GEN_1053 : trans_1_io_pipe_phv_out_data_81; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2116 = 2'h1 != last_proc_id ? _GEN_1054 : trans_1_io_pipe_phv_out_data_82; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2117 = 2'h1 != last_proc_id ? _GEN_1055 : trans_1_io_pipe_phv_out_data_83; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2118 = 2'h1 != last_proc_id ? _GEN_1056 : trans_1_io_pipe_phv_out_data_84; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2119 = 2'h1 != last_proc_id ? _GEN_1057 : trans_1_io_pipe_phv_out_data_85; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2120 = 2'h1 != last_proc_id ? _GEN_1058 : trans_1_io_pipe_phv_out_data_86; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2121 = 2'h1 != last_proc_id ? _GEN_1059 : trans_1_io_pipe_phv_out_data_87; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2122 = 2'h1 != last_proc_id ? _GEN_1060 : trans_1_io_pipe_phv_out_data_88; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2123 = 2'h1 != last_proc_id ? _GEN_1061 : trans_1_io_pipe_phv_out_data_89; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2124 = 2'h1 != last_proc_id ? _GEN_1062 : trans_1_io_pipe_phv_out_data_90; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2125 = 2'h1 != last_proc_id ? _GEN_1063 : trans_1_io_pipe_phv_out_data_91; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2126 = 2'h1 != last_proc_id ? _GEN_1064 : trans_1_io_pipe_phv_out_data_92; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2127 = 2'h1 != last_proc_id ? _GEN_1065 : trans_1_io_pipe_phv_out_data_93; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2128 = 2'h1 != last_proc_id ? _GEN_1066 : trans_1_io_pipe_phv_out_data_94; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_2129 = 2'h1 != last_proc_id ? _GEN_1067 : trans_1_io_pipe_phv_out_data_95; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire  _GEN_2130 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_is_valid_processor : _GEN_1540; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire  _GEN_2131 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_next_config_id : _GEN_1541; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [1:0] _GEN_2132 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_next_processor_id : _GEN_1542; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2133 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_parse_transition_field : _GEN_1543; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2134 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_parse_current_offset : _GEN_1544; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2135 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_parse_current_state : _GEN_1545; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2136 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_0 : _GEN_1546; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2137 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_1 : _GEN_1547; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2138 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_2 : _GEN_1548; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2139 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_3 : _GEN_1549; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2140 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_4 : _GEN_1550; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2141 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_5 : _GEN_1551; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2142 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_6 : _GEN_1552; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2143 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_7 : _GEN_1553; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2144 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_8 : _GEN_1554; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2145 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_9 : _GEN_1555; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2146 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_10 : _GEN_1556; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2147 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_11 : _GEN_1557; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2148 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_12 : _GEN_1558; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2149 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_13 : _GEN_1559; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2150 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_14 : _GEN_1560; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2151 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_15 : _GEN_1561; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2152 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_0 : _GEN_1562; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2153 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_1 : _GEN_1563; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2154 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_2 : _GEN_1564; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2155 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_3 : _GEN_1565; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2156 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_4 : _GEN_1566; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2157 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_5 : _GEN_1567; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2158 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_6 : _GEN_1568; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2159 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_7 : _GEN_1569; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2160 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_8 : _GEN_1570; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2161 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_9 : _GEN_1571; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2162 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_10 : _GEN_1572; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2163 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_11 : _GEN_1573; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2164 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_12 : _GEN_1574; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2165 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_13 : _GEN_1575; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2166 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_14 : _GEN_1576; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2167 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_15 : _GEN_1577; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2168 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_16 : _GEN_1578; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2169 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_17 : _GEN_1579; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2170 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_18 : _GEN_1580; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2171 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_19 : _GEN_1581; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2172 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_20 : _GEN_1582; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2173 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_21 : _GEN_1583; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2174 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_22 : _GEN_1584; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2175 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_23 : _GEN_1585; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2176 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_24 : _GEN_1586; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2177 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_25 : _GEN_1587; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2178 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_26 : _GEN_1588; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2179 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_27 : _GEN_1589; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2180 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_28 : _GEN_1590; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2181 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_29 : _GEN_1591; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2182 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_30 : _GEN_1592; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2183 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_31 : _GEN_1593; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2184 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_32 : _GEN_1594; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2185 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_33 : _GEN_1595; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2186 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_34 : _GEN_1596; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2187 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_35 : _GEN_1597; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2188 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_36 : _GEN_1598; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2189 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_37 : _GEN_1599; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2190 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_38 : _GEN_1600; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2191 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_39 : _GEN_1601; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2192 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_40 : _GEN_1602; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2193 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_41 : _GEN_1603; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2194 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_42 : _GEN_1604; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2195 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_43 : _GEN_1605; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2196 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_44 : _GEN_1606; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2197 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_45 : _GEN_1607; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2198 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_46 : _GEN_1608; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2199 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_47 : _GEN_1609; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2200 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_48 : _GEN_1610; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2201 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_49 : _GEN_1611; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2202 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_50 : _GEN_1612; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2203 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_51 : _GEN_1613; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2204 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_52 : _GEN_1614; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2205 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_53 : _GEN_1615; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2206 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_54 : _GEN_1616; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2207 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_55 : _GEN_1617; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2208 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_56 : _GEN_1618; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2209 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_57 : _GEN_1619; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2210 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_58 : _GEN_1620; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2211 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_59 : _GEN_1621; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2212 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_60 : _GEN_1622; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2213 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_61 : _GEN_1623; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2214 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_62 : _GEN_1624; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2215 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_63 : _GEN_1625; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2216 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_64 : _GEN_1626; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2217 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_65 : _GEN_1627; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2218 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_66 : _GEN_1628; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2219 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_67 : _GEN_1629; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2220 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_68 : _GEN_1630; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2221 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_69 : _GEN_1631; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2222 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_70 : _GEN_1632; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2223 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_71 : _GEN_1633; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2224 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_72 : _GEN_1634; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2225 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_73 : _GEN_1635; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2226 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_74 : _GEN_1636; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2227 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_75 : _GEN_1637; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2228 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_76 : _GEN_1638; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2229 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_77 : _GEN_1639; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2230 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_78 : _GEN_1640; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2231 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_79 : _GEN_1641; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2232 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_80 : _GEN_1642; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2233 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_81 : _GEN_1643; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2234 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_82 : _GEN_1644; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2235 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_83 : _GEN_1645; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2236 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_84 : _GEN_1646; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2237 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_85 : _GEN_1647; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2238 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_86 : _GEN_1648; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2239 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_87 : _GEN_1649; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2240 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_88 : _GEN_1650; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2241 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_89 : _GEN_1651; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2242 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_90 : _GEN_1652; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2243 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_91 : _GEN_1653; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2244 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_92 : _GEN_1654; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2245 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_93 : _GEN_1655; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2246 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_94 : _GEN_1656; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2247 = 2'h0 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_95 : _GEN_1657; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire  _GEN_2248 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_is_valid_processor : _GEN_1658; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire  _GEN_2249 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_next_config_id : _GEN_1659; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [1:0] _GEN_2250 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_next_processor_id : _GEN_1660; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2251 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_parse_transition_field : _GEN_1661; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2252 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_parse_current_offset : _GEN_1662; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2253 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_parse_current_state : _GEN_1663; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2254 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_0 : _GEN_1664; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2255 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_1 : _GEN_1665; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2256 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_2 : _GEN_1666; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2257 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_3 : _GEN_1667; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2258 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_4 : _GEN_1668; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2259 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_5 : _GEN_1669; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2260 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_6 : _GEN_1670; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2261 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_7 : _GEN_1671; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2262 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_8 : _GEN_1672; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2263 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_9 : _GEN_1673; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2264 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_10 : _GEN_1674; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2265 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_11 : _GEN_1675; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2266 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_12 : _GEN_1676; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2267 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_13 : _GEN_1677; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2268 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_14 : _GEN_1678; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2269 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_15 : _GEN_1679; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2270 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_0 : _GEN_1680; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2271 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_1 : _GEN_1681; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2272 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_2 : _GEN_1682; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2273 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_3 : _GEN_1683; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2274 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_4 : _GEN_1684; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2275 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_5 : _GEN_1685; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2276 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_6 : _GEN_1686; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2277 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_7 : _GEN_1687; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2278 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_8 : _GEN_1688; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2279 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_9 : _GEN_1689; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2280 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_10 : _GEN_1690; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2281 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_11 : _GEN_1691; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2282 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_12 : _GEN_1692; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2283 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_13 : _GEN_1693; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2284 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_14 : _GEN_1694; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2285 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_15 : _GEN_1695; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2286 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_16 : _GEN_1696; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2287 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_17 : _GEN_1697; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2288 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_18 : _GEN_1698; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2289 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_19 : _GEN_1699; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2290 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_20 : _GEN_1700; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2291 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_21 : _GEN_1701; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2292 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_22 : _GEN_1702; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2293 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_23 : _GEN_1703; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2294 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_24 : _GEN_1704; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2295 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_25 : _GEN_1705; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2296 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_26 : _GEN_1706; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2297 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_27 : _GEN_1707; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2298 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_28 : _GEN_1708; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2299 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_29 : _GEN_1709; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2300 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_30 : _GEN_1710; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2301 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_31 : _GEN_1711; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2302 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_32 : _GEN_1712; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2303 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_33 : _GEN_1713; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2304 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_34 : _GEN_1714; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2305 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_35 : _GEN_1715; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2306 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_36 : _GEN_1716; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2307 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_37 : _GEN_1717; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2308 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_38 : _GEN_1718; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2309 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_39 : _GEN_1719; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2310 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_40 : _GEN_1720; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2311 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_41 : _GEN_1721; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2312 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_42 : _GEN_1722; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2313 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_43 : _GEN_1723; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2314 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_44 : _GEN_1724; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2315 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_45 : _GEN_1725; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2316 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_46 : _GEN_1726; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2317 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_47 : _GEN_1727; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2318 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_48 : _GEN_1728; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2319 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_49 : _GEN_1729; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2320 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_50 : _GEN_1730; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2321 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_51 : _GEN_1731; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2322 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_52 : _GEN_1732; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2323 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_53 : _GEN_1733; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2324 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_54 : _GEN_1734; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2325 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_55 : _GEN_1735; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2326 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_56 : _GEN_1736; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2327 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_57 : _GEN_1737; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2328 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_58 : _GEN_1738; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2329 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_59 : _GEN_1739; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2330 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_60 : _GEN_1740; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2331 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_61 : _GEN_1741; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2332 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_62 : _GEN_1742; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2333 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_63 : _GEN_1743; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2334 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_64 : _GEN_1744; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2335 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_65 : _GEN_1745; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2336 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_66 : _GEN_1746; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2337 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_67 : _GEN_1747; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2338 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_68 : _GEN_1748; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2339 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_69 : _GEN_1749; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2340 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_70 : _GEN_1750; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2341 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_71 : _GEN_1751; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2342 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_72 : _GEN_1752; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2343 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_73 : _GEN_1753; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2344 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_74 : _GEN_1754; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2345 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_75 : _GEN_1755; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2346 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_76 : _GEN_1756; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2347 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_77 : _GEN_1757; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2348 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_78 : _GEN_1758; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2349 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_79 : _GEN_1759; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2350 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_80 : _GEN_1760; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2351 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_81 : _GEN_1761; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2352 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_82 : _GEN_1762; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2353 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_83 : _GEN_1763; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2354 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_84 : _GEN_1764; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2355 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_85 : _GEN_1765; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2356 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_86 : _GEN_1766; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2357 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_87 : _GEN_1767; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2358 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_88 : _GEN_1768; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2359 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_89 : _GEN_1769; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2360 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_90 : _GEN_1770; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2361 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_91 : _GEN_1771; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2362 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_92 : _GEN_1772; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2363 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_93 : _GEN_1773; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2364 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_94 : _GEN_1774; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2365 = 2'h1 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_95 : _GEN_1775; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire  _GEN_2366 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_is_valid_processor : _GEN_1776; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire  _GEN_2367 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_next_config_id : _GEN_1777; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [1:0] _GEN_2368 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_next_processor_id : _GEN_1778; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2369 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_parse_transition_field : _GEN_1779; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2370 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_parse_current_offset : _GEN_1780; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2371 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_parse_current_state : _GEN_1781; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2372 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_0 : _GEN_1782; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2373 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_1 : _GEN_1783; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2374 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_2 : _GEN_1784; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2375 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_3 : _GEN_1785; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2376 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_4 : _GEN_1786; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2377 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_5 : _GEN_1787; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2378 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_6 : _GEN_1788; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2379 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_7 : _GEN_1789; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2380 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_8 : _GEN_1790; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2381 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_9 : _GEN_1791; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2382 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_10 : _GEN_1792; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2383 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_11 : _GEN_1793; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2384 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_12 : _GEN_1794; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2385 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_13 : _GEN_1795; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2386 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_14 : _GEN_1796; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2387 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_15 : _GEN_1797; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2388 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_0 : _GEN_1798; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2389 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_1 : _GEN_1799; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2390 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_2 : _GEN_1800; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2391 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_3 : _GEN_1801; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2392 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_4 : _GEN_1802; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2393 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_5 : _GEN_1803; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2394 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_6 : _GEN_1804; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2395 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_7 : _GEN_1805; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2396 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_8 : _GEN_1806; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2397 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_9 : _GEN_1807; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2398 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_10 : _GEN_1808; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2399 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_11 : _GEN_1809; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2400 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_12 : _GEN_1810; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2401 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_13 : _GEN_1811; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2402 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_14 : _GEN_1812; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2403 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_15 : _GEN_1813; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2404 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_16 : _GEN_1814; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2405 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_17 : _GEN_1815; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2406 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_18 : _GEN_1816; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2407 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_19 : _GEN_1817; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2408 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_20 : _GEN_1818; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2409 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_21 : _GEN_1819; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2410 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_22 : _GEN_1820; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2411 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_23 : _GEN_1821; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2412 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_24 : _GEN_1822; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2413 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_25 : _GEN_1823; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2414 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_26 : _GEN_1824; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2415 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_27 : _GEN_1825; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2416 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_28 : _GEN_1826; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2417 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_29 : _GEN_1827; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2418 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_30 : _GEN_1828; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2419 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_31 : _GEN_1829; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2420 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_32 : _GEN_1830; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2421 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_33 : _GEN_1831; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2422 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_34 : _GEN_1832; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2423 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_35 : _GEN_1833; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2424 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_36 : _GEN_1834; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2425 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_37 : _GEN_1835; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2426 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_38 : _GEN_1836; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2427 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_39 : _GEN_1837; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2428 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_40 : _GEN_1838; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2429 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_41 : _GEN_1839; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2430 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_42 : _GEN_1840; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2431 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_43 : _GEN_1841; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2432 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_44 : _GEN_1842; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2433 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_45 : _GEN_1843; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2434 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_46 : _GEN_1844; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2435 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_47 : _GEN_1845; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2436 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_48 : _GEN_1846; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2437 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_49 : _GEN_1847; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2438 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_50 : _GEN_1848; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2439 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_51 : _GEN_1849; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2440 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_52 : _GEN_1850; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2441 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_53 : _GEN_1851; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2442 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_54 : _GEN_1852; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2443 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_55 : _GEN_1853; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2444 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_56 : _GEN_1854; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2445 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_57 : _GEN_1855; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2446 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_58 : _GEN_1856; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2447 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_59 : _GEN_1857; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2448 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_60 : _GEN_1858; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2449 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_61 : _GEN_1859; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2450 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_62 : _GEN_1860; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2451 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_63 : _GEN_1861; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2452 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_64 : _GEN_1862; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2453 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_65 : _GEN_1863; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2454 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_66 : _GEN_1864; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2455 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_67 : _GEN_1865; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2456 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_68 : _GEN_1866; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2457 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_69 : _GEN_1867; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2458 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_70 : _GEN_1868; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2459 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_71 : _GEN_1869; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2460 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_72 : _GEN_1870; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2461 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_73 : _GEN_1871; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2462 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_74 : _GEN_1872; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2463 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_75 : _GEN_1873; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2464 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_76 : _GEN_1874; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2465 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_77 : _GEN_1875; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2466 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_78 : _GEN_1876; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2467 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_79 : _GEN_1877; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2468 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_80 : _GEN_1878; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2469 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_81 : _GEN_1879; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2470 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_82 : _GEN_1880; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2471 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_83 : _GEN_1881; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2472 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_84 : _GEN_1882; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2473 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_85 : _GEN_1883; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2474 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_86 : _GEN_1884; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2475 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_87 : _GEN_1885; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2476 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_88 : _GEN_1886; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2477 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_89 : _GEN_1887; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2478 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_90 : _GEN_1888; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2479 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_91 : _GEN_1889; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2480 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_92 : _GEN_1890; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2481 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_93 : _GEN_1891; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2482 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_94 : _GEN_1892; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2483 = 2'h2 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_95 : _GEN_1893; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire  _GEN_2484 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_is_valid_processor : _GEN_1894; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire  _GEN_2485 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_next_config_id : _GEN_1895; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [1:0] _GEN_2486 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_next_processor_id : _GEN_1896; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2487 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_parse_transition_field : _GEN_1897; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2488 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_parse_current_offset : _GEN_1898; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2489 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_parse_current_state : _GEN_1899; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2490 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_0 : _GEN_1900; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2491 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_1 : _GEN_1901; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2492 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_2 : _GEN_1902; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2493 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_3 : _GEN_1903; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2494 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_4 : _GEN_1904; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2495 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_5 : _GEN_1905; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2496 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_6 : _GEN_1906; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2497 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_7 : _GEN_1907; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2498 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_8 : _GEN_1908; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2499 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_9 : _GEN_1909; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2500 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_10 : _GEN_1910; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2501 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_11 : _GEN_1911; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2502 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_12 : _GEN_1912; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2503 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_13 : _GEN_1913; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2504 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_14 : _GEN_1914; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_2505 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_header_15 : _GEN_1915; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2506 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_0 : _GEN_1916; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2507 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_1 : _GEN_1917; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2508 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_2 : _GEN_1918; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2509 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_3 : _GEN_1919; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2510 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_4 : _GEN_1920; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2511 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_5 : _GEN_1921; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2512 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_6 : _GEN_1922; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2513 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_7 : _GEN_1923; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2514 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_8 : _GEN_1924; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2515 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_9 : _GEN_1925; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2516 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_10 : _GEN_1926; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2517 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_11 : _GEN_1927; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2518 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_12 : _GEN_1928; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2519 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_13 : _GEN_1929; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2520 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_14 : _GEN_1930; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2521 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_15 : _GEN_1931; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2522 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_16 : _GEN_1932; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2523 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_17 : _GEN_1933; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2524 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_18 : _GEN_1934; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2525 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_19 : _GEN_1935; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2526 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_20 : _GEN_1936; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2527 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_21 : _GEN_1937; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2528 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_22 : _GEN_1938; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2529 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_23 : _GEN_1939; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2530 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_24 : _GEN_1940; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2531 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_25 : _GEN_1941; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2532 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_26 : _GEN_1942; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2533 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_27 : _GEN_1943; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2534 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_28 : _GEN_1944; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2535 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_29 : _GEN_1945; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2536 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_30 : _GEN_1946; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2537 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_31 : _GEN_1947; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2538 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_32 : _GEN_1948; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2539 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_33 : _GEN_1949; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2540 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_34 : _GEN_1950; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2541 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_35 : _GEN_1951; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2542 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_36 : _GEN_1952; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2543 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_37 : _GEN_1953; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2544 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_38 : _GEN_1954; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2545 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_39 : _GEN_1955; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2546 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_40 : _GEN_1956; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2547 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_41 : _GEN_1957; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2548 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_42 : _GEN_1958; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2549 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_43 : _GEN_1959; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2550 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_44 : _GEN_1960; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2551 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_45 : _GEN_1961; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2552 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_46 : _GEN_1962; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2553 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_47 : _GEN_1963; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2554 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_48 : _GEN_1964; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2555 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_49 : _GEN_1965; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2556 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_50 : _GEN_1966; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2557 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_51 : _GEN_1967; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2558 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_52 : _GEN_1968; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2559 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_53 : _GEN_1969; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2560 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_54 : _GEN_1970; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2561 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_55 : _GEN_1971; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2562 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_56 : _GEN_1972; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2563 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_57 : _GEN_1973; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2564 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_58 : _GEN_1974; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2565 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_59 : _GEN_1975; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2566 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_60 : _GEN_1976; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2567 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_61 : _GEN_1977; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2568 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_62 : _GEN_1978; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2569 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_63 : _GEN_1979; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2570 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_64 : _GEN_1980; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2571 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_65 : _GEN_1981; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2572 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_66 : _GEN_1982; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2573 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_67 : _GEN_1983; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2574 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_68 : _GEN_1984; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2575 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_69 : _GEN_1985; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2576 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_70 : _GEN_1986; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2577 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_71 : _GEN_1987; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2578 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_72 : _GEN_1988; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2579 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_73 : _GEN_1989; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2580 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_74 : _GEN_1990; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2581 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_75 : _GEN_1991; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2582 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_76 : _GEN_1992; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2583 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_77 : _GEN_1993; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2584 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_78 : _GEN_1994; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2585 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_79 : _GEN_1995; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2586 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_80 : _GEN_1996; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2587 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_81 : _GEN_1997; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2588 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_82 : _GEN_1998; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2589 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_83 : _GEN_1999; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2590 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_84 : _GEN_2000; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2591 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_85 : _GEN_2001; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2592 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_86 : _GEN_2002; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2593 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_87 : _GEN_2003; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2594 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_88 : _GEN_2004; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2595 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_89 : _GEN_2005; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2596 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_90 : _GEN_2006; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2597 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_91 : _GEN_2007; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2598 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_92 : _GEN_2008; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2599 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_93 : _GEN_2009; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2600 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_94 : _GEN_2010; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_2601 = 2'h3 == next_proc_id_2 ? trans_2_io_pipe_phv_out_data_95 : _GEN_2011; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire  _GEN_2602 = 2'h2 != last_proc_id ? _GEN_2130 : _GEN_1540; // @[ipsa.scala 94:65]
  wire  _GEN_2603 = 2'h2 != last_proc_id ? _GEN_2131 : _GEN_1541; // @[ipsa.scala 94:65]
  wire [1:0] _GEN_2604 = 2'h2 != last_proc_id ? _GEN_2132 : _GEN_1542; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2605 = 2'h2 != last_proc_id ? _GEN_2133 : _GEN_1543; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2606 = 2'h2 != last_proc_id ? _GEN_2134 : _GEN_1544; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2607 = 2'h2 != last_proc_id ? _GEN_2135 : _GEN_1545; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2608 = 2'h2 != last_proc_id ? _GEN_2136 : _GEN_1546; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2609 = 2'h2 != last_proc_id ? _GEN_2137 : _GEN_1547; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2610 = 2'h2 != last_proc_id ? _GEN_2138 : _GEN_1548; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2611 = 2'h2 != last_proc_id ? _GEN_2139 : _GEN_1549; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2612 = 2'h2 != last_proc_id ? _GEN_2140 : _GEN_1550; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2613 = 2'h2 != last_proc_id ? _GEN_2141 : _GEN_1551; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2614 = 2'h2 != last_proc_id ? _GEN_2142 : _GEN_1552; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2615 = 2'h2 != last_proc_id ? _GEN_2143 : _GEN_1553; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2616 = 2'h2 != last_proc_id ? _GEN_2144 : _GEN_1554; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2617 = 2'h2 != last_proc_id ? _GEN_2145 : _GEN_1555; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2618 = 2'h2 != last_proc_id ? _GEN_2146 : _GEN_1556; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2619 = 2'h2 != last_proc_id ? _GEN_2147 : _GEN_1557; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2620 = 2'h2 != last_proc_id ? _GEN_2148 : _GEN_1558; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2621 = 2'h2 != last_proc_id ? _GEN_2149 : _GEN_1559; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2622 = 2'h2 != last_proc_id ? _GEN_2150 : _GEN_1560; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2623 = 2'h2 != last_proc_id ? _GEN_2151 : _GEN_1561; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2624 = 2'h2 != last_proc_id ? _GEN_2152 : _GEN_1562; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2625 = 2'h2 != last_proc_id ? _GEN_2153 : _GEN_1563; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2626 = 2'h2 != last_proc_id ? _GEN_2154 : _GEN_1564; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2627 = 2'h2 != last_proc_id ? _GEN_2155 : _GEN_1565; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2628 = 2'h2 != last_proc_id ? _GEN_2156 : _GEN_1566; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2629 = 2'h2 != last_proc_id ? _GEN_2157 : _GEN_1567; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2630 = 2'h2 != last_proc_id ? _GEN_2158 : _GEN_1568; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2631 = 2'h2 != last_proc_id ? _GEN_2159 : _GEN_1569; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2632 = 2'h2 != last_proc_id ? _GEN_2160 : _GEN_1570; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2633 = 2'h2 != last_proc_id ? _GEN_2161 : _GEN_1571; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2634 = 2'h2 != last_proc_id ? _GEN_2162 : _GEN_1572; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2635 = 2'h2 != last_proc_id ? _GEN_2163 : _GEN_1573; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2636 = 2'h2 != last_proc_id ? _GEN_2164 : _GEN_1574; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2637 = 2'h2 != last_proc_id ? _GEN_2165 : _GEN_1575; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2638 = 2'h2 != last_proc_id ? _GEN_2166 : _GEN_1576; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2639 = 2'h2 != last_proc_id ? _GEN_2167 : _GEN_1577; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2640 = 2'h2 != last_proc_id ? _GEN_2168 : _GEN_1578; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2641 = 2'h2 != last_proc_id ? _GEN_2169 : _GEN_1579; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2642 = 2'h2 != last_proc_id ? _GEN_2170 : _GEN_1580; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2643 = 2'h2 != last_proc_id ? _GEN_2171 : _GEN_1581; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2644 = 2'h2 != last_proc_id ? _GEN_2172 : _GEN_1582; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2645 = 2'h2 != last_proc_id ? _GEN_2173 : _GEN_1583; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2646 = 2'h2 != last_proc_id ? _GEN_2174 : _GEN_1584; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2647 = 2'h2 != last_proc_id ? _GEN_2175 : _GEN_1585; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2648 = 2'h2 != last_proc_id ? _GEN_2176 : _GEN_1586; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2649 = 2'h2 != last_proc_id ? _GEN_2177 : _GEN_1587; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2650 = 2'h2 != last_proc_id ? _GEN_2178 : _GEN_1588; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2651 = 2'h2 != last_proc_id ? _GEN_2179 : _GEN_1589; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2652 = 2'h2 != last_proc_id ? _GEN_2180 : _GEN_1590; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2653 = 2'h2 != last_proc_id ? _GEN_2181 : _GEN_1591; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2654 = 2'h2 != last_proc_id ? _GEN_2182 : _GEN_1592; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2655 = 2'h2 != last_proc_id ? _GEN_2183 : _GEN_1593; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2656 = 2'h2 != last_proc_id ? _GEN_2184 : _GEN_1594; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2657 = 2'h2 != last_proc_id ? _GEN_2185 : _GEN_1595; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2658 = 2'h2 != last_proc_id ? _GEN_2186 : _GEN_1596; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2659 = 2'h2 != last_proc_id ? _GEN_2187 : _GEN_1597; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2660 = 2'h2 != last_proc_id ? _GEN_2188 : _GEN_1598; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2661 = 2'h2 != last_proc_id ? _GEN_2189 : _GEN_1599; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2662 = 2'h2 != last_proc_id ? _GEN_2190 : _GEN_1600; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2663 = 2'h2 != last_proc_id ? _GEN_2191 : _GEN_1601; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2664 = 2'h2 != last_proc_id ? _GEN_2192 : _GEN_1602; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2665 = 2'h2 != last_proc_id ? _GEN_2193 : _GEN_1603; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2666 = 2'h2 != last_proc_id ? _GEN_2194 : _GEN_1604; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2667 = 2'h2 != last_proc_id ? _GEN_2195 : _GEN_1605; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2668 = 2'h2 != last_proc_id ? _GEN_2196 : _GEN_1606; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2669 = 2'h2 != last_proc_id ? _GEN_2197 : _GEN_1607; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2670 = 2'h2 != last_proc_id ? _GEN_2198 : _GEN_1608; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2671 = 2'h2 != last_proc_id ? _GEN_2199 : _GEN_1609; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2672 = 2'h2 != last_proc_id ? _GEN_2200 : _GEN_1610; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2673 = 2'h2 != last_proc_id ? _GEN_2201 : _GEN_1611; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2674 = 2'h2 != last_proc_id ? _GEN_2202 : _GEN_1612; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2675 = 2'h2 != last_proc_id ? _GEN_2203 : _GEN_1613; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2676 = 2'h2 != last_proc_id ? _GEN_2204 : _GEN_1614; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2677 = 2'h2 != last_proc_id ? _GEN_2205 : _GEN_1615; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2678 = 2'h2 != last_proc_id ? _GEN_2206 : _GEN_1616; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2679 = 2'h2 != last_proc_id ? _GEN_2207 : _GEN_1617; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2680 = 2'h2 != last_proc_id ? _GEN_2208 : _GEN_1618; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2681 = 2'h2 != last_proc_id ? _GEN_2209 : _GEN_1619; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2682 = 2'h2 != last_proc_id ? _GEN_2210 : _GEN_1620; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2683 = 2'h2 != last_proc_id ? _GEN_2211 : _GEN_1621; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2684 = 2'h2 != last_proc_id ? _GEN_2212 : _GEN_1622; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2685 = 2'h2 != last_proc_id ? _GEN_2213 : _GEN_1623; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2686 = 2'h2 != last_proc_id ? _GEN_2214 : _GEN_1624; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2687 = 2'h2 != last_proc_id ? _GEN_2215 : _GEN_1625; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2688 = 2'h2 != last_proc_id ? _GEN_2216 : _GEN_1626; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2689 = 2'h2 != last_proc_id ? _GEN_2217 : _GEN_1627; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2690 = 2'h2 != last_proc_id ? _GEN_2218 : _GEN_1628; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2691 = 2'h2 != last_proc_id ? _GEN_2219 : _GEN_1629; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2692 = 2'h2 != last_proc_id ? _GEN_2220 : _GEN_1630; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2693 = 2'h2 != last_proc_id ? _GEN_2221 : _GEN_1631; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2694 = 2'h2 != last_proc_id ? _GEN_2222 : _GEN_1632; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2695 = 2'h2 != last_proc_id ? _GEN_2223 : _GEN_1633; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2696 = 2'h2 != last_proc_id ? _GEN_2224 : _GEN_1634; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2697 = 2'h2 != last_proc_id ? _GEN_2225 : _GEN_1635; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2698 = 2'h2 != last_proc_id ? _GEN_2226 : _GEN_1636; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2699 = 2'h2 != last_proc_id ? _GEN_2227 : _GEN_1637; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2700 = 2'h2 != last_proc_id ? _GEN_2228 : _GEN_1638; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2701 = 2'h2 != last_proc_id ? _GEN_2229 : _GEN_1639; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2702 = 2'h2 != last_proc_id ? _GEN_2230 : _GEN_1640; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2703 = 2'h2 != last_proc_id ? _GEN_2231 : _GEN_1641; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2704 = 2'h2 != last_proc_id ? _GEN_2232 : _GEN_1642; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2705 = 2'h2 != last_proc_id ? _GEN_2233 : _GEN_1643; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2706 = 2'h2 != last_proc_id ? _GEN_2234 : _GEN_1644; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2707 = 2'h2 != last_proc_id ? _GEN_2235 : _GEN_1645; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2708 = 2'h2 != last_proc_id ? _GEN_2236 : _GEN_1646; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2709 = 2'h2 != last_proc_id ? _GEN_2237 : _GEN_1647; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2710 = 2'h2 != last_proc_id ? _GEN_2238 : _GEN_1648; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2711 = 2'h2 != last_proc_id ? _GEN_2239 : _GEN_1649; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2712 = 2'h2 != last_proc_id ? _GEN_2240 : _GEN_1650; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2713 = 2'h2 != last_proc_id ? _GEN_2241 : _GEN_1651; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2714 = 2'h2 != last_proc_id ? _GEN_2242 : _GEN_1652; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2715 = 2'h2 != last_proc_id ? _GEN_2243 : _GEN_1653; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2716 = 2'h2 != last_proc_id ? _GEN_2244 : _GEN_1654; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2717 = 2'h2 != last_proc_id ? _GEN_2245 : _GEN_1655; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2718 = 2'h2 != last_proc_id ? _GEN_2246 : _GEN_1656; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2719 = 2'h2 != last_proc_id ? _GEN_2247 : _GEN_1657; // @[ipsa.scala 94:65]
  wire  _GEN_2720 = 2'h2 != last_proc_id ? _GEN_2248 : _GEN_1658; // @[ipsa.scala 94:65]
  wire  _GEN_2721 = 2'h2 != last_proc_id ? _GEN_2249 : _GEN_1659; // @[ipsa.scala 94:65]
  wire [1:0] _GEN_2722 = 2'h2 != last_proc_id ? _GEN_2250 : _GEN_1660; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2723 = 2'h2 != last_proc_id ? _GEN_2251 : _GEN_1661; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2724 = 2'h2 != last_proc_id ? _GEN_2252 : _GEN_1662; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2725 = 2'h2 != last_proc_id ? _GEN_2253 : _GEN_1663; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2726 = 2'h2 != last_proc_id ? _GEN_2254 : _GEN_1664; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2727 = 2'h2 != last_proc_id ? _GEN_2255 : _GEN_1665; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2728 = 2'h2 != last_proc_id ? _GEN_2256 : _GEN_1666; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2729 = 2'h2 != last_proc_id ? _GEN_2257 : _GEN_1667; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2730 = 2'h2 != last_proc_id ? _GEN_2258 : _GEN_1668; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2731 = 2'h2 != last_proc_id ? _GEN_2259 : _GEN_1669; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2732 = 2'h2 != last_proc_id ? _GEN_2260 : _GEN_1670; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2733 = 2'h2 != last_proc_id ? _GEN_2261 : _GEN_1671; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2734 = 2'h2 != last_proc_id ? _GEN_2262 : _GEN_1672; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2735 = 2'h2 != last_proc_id ? _GEN_2263 : _GEN_1673; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2736 = 2'h2 != last_proc_id ? _GEN_2264 : _GEN_1674; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2737 = 2'h2 != last_proc_id ? _GEN_2265 : _GEN_1675; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2738 = 2'h2 != last_proc_id ? _GEN_2266 : _GEN_1676; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2739 = 2'h2 != last_proc_id ? _GEN_2267 : _GEN_1677; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2740 = 2'h2 != last_proc_id ? _GEN_2268 : _GEN_1678; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2741 = 2'h2 != last_proc_id ? _GEN_2269 : _GEN_1679; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2742 = 2'h2 != last_proc_id ? _GEN_2270 : _GEN_1680; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2743 = 2'h2 != last_proc_id ? _GEN_2271 : _GEN_1681; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2744 = 2'h2 != last_proc_id ? _GEN_2272 : _GEN_1682; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2745 = 2'h2 != last_proc_id ? _GEN_2273 : _GEN_1683; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2746 = 2'h2 != last_proc_id ? _GEN_2274 : _GEN_1684; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2747 = 2'h2 != last_proc_id ? _GEN_2275 : _GEN_1685; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2748 = 2'h2 != last_proc_id ? _GEN_2276 : _GEN_1686; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2749 = 2'h2 != last_proc_id ? _GEN_2277 : _GEN_1687; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2750 = 2'h2 != last_proc_id ? _GEN_2278 : _GEN_1688; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2751 = 2'h2 != last_proc_id ? _GEN_2279 : _GEN_1689; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2752 = 2'h2 != last_proc_id ? _GEN_2280 : _GEN_1690; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2753 = 2'h2 != last_proc_id ? _GEN_2281 : _GEN_1691; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2754 = 2'h2 != last_proc_id ? _GEN_2282 : _GEN_1692; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2755 = 2'h2 != last_proc_id ? _GEN_2283 : _GEN_1693; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2756 = 2'h2 != last_proc_id ? _GEN_2284 : _GEN_1694; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2757 = 2'h2 != last_proc_id ? _GEN_2285 : _GEN_1695; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2758 = 2'h2 != last_proc_id ? _GEN_2286 : _GEN_1696; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2759 = 2'h2 != last_proc_id ? _GEN_2287 : _GEN_1697; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2760 = 2'h2 != last_proc_id ? _GEN_2288 : _GEN_1698; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2761 = 2'h2 != last_proc_id ? _GEN_2289 : _GEN_1699; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2762 = 2'h2 != last_proc_id ? _GEN_2290 : _GEN_1700; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2763 = 2'h2 != last_proc_id ? _GEN_2291 : _GEN_1701; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2764 = 2'h2 != last_proc_id ? _GEN_2292 : _GEN_1702; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2765 = 2'h2 != last_proc_id ? _GEN_2293 : _GEN_1703; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2766 = 2'h2 != last_proc_id ? _GEN_2294 : _GEN_1704; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2767 = 2'h2 != last_proc_id ? _GEN_2295 : _GEN_1705; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2768 = 2'h2 != last_proc_id ? _GEN_2296 : _GEN_1706; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2769 = 2'h2 != last_proc_id ? _GEN_2297 : _GEN_1707; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2770 = 2'h2 != last_proc_id ? _GEN_2298 : _GEN_1708; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2771 = 2'h2 != last_proc_id ? _GEN_2299 : _GEN_1709; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2772 = 2'h2 != last_proc_id ? _GEN_2300 : _GEN_1710; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2773 = 2'h2 != last_proc_id ? _GEN_2301 : _GEN_1711; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2774 = 2'h2 != last_proc_id ? _GEN_2302 : _GEN_1712; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2775 = 2'h2 != last_proc_id ? _GEN_2303 : _GEN_1713; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2776 = 2'h2 != last_proc_id ? _GEN_2304 : _GEN_1714; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2777 = 2'h2 != last_proc_id ? _GEN_2305 : _GEN_1715; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2778 = 2'h2 != last_proc_id ? _GEN_2306 : _GEN_1716; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2779 = 2'h2 != last_proc_id ? _GEN_2307 : _GEN_1717; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2780 = 2'h2 != last_proc_id ? _GEN_2308 : _GEN_1718; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2781 = 2'h2 != last_proc_id ? _GEN_2309 : _GEN_1719; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2782 = 2'h2 != last_proc_id ? _GEN_2310 : _GEN_1720; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2783 = 2'h2 != last_proc_id ? _GEN_2311 : _GEN_1721; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2784 = 2'h2 != last_proc_id ? _GEN_2312 : _GEN_1722; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2785 = 2'h2 != last_proc_id ? _GEN_2313 : _GEN_1723; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2786 = 2'h2 != last_proc_id ? _GEN_2314 : _GEN_1724; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2787 = 2'h2 != last_proc_id ? _GEN_2315 : _GEN_1725; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2788 = 2'h2 != last_proc_id ? _GEN_2316 : _GEN_1726; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2789 = 2'h2 != last_proc_id ? _GEN_2317 : _GEN_1727; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2790 = 2'h2 != last_proc_id ? _GEN_2318 : _GEN_1728; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2791 = 2'h2 != last_proc_id ? _GEN_2319 : _GEN_1729; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2792 = 2'h2 != last_proc_id ? _GEN_2320 : _GEN_1730; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2793 = 2'h2 != last_proc_id ? _GEN_2321 : _GEN_1731; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2794 = 2'h2 != last_proc_id ? _GEN_2322 : _GEN_1732; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2795 = 2'h2 != last_proc_id ? _GEN_2323 : _GEN_1733; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2796 = 2'h2 != last_proc_id ? _GEN_2324 : _GEN_1734; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2797 = 2'h2 != last_proc_id ? _GEN_2325 : _GEN_1735; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2798 = 2'h2 != last_proc_id ? _GEN_2326 : _GEN_1736; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2799 = 2'h2 != last_proc_id ? _GEN_2327 : _GEN_1737; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2800 = 2'h2 != last_proc_id ? _GEN_2328 : _GEN_1738; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2801 = 2'h2 != last_proc_id ? _GEN_2329 : _GEN_1739; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2802 = 2'h2 != last_proc_id ? _GEN_2330 : _GEN_1740; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2803 = 2'h2 != last_proc_id ? _GEN_2331 : _GEN_1741; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2804 = 2'h2 != last_proc_id ? _GEN_2332 : _GEN_1742; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2805 = 2'h2 != last_proc_id ? _GEN_2333 : _GEN_1743; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2806 = 2'h2 != last_proc_id ? _GEN_2334 : _GEN_1744; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2807 = 2'h2 != last_proc_id ? _GEN_2335 : _GEN_1745; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2808 = 2'h2 != last_proc_id ? _GEN_2336 : _GEN_1746; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2809 = 2'h2 != last_proc_id ? _GEN_2337 : _GEN_1747; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2810 = 2'h2 != last_proc_id ? _GEN_2338 : _GEN_1748; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2811 = 2'h2 != last_proc_id ? _GEN_2339 : _GEN_1749; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2812 = 2'h2 != last_proc_id ? _GEN_2340 : _GEN_1750; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2813 = 2'h2 != last_proc_id ? _GEN_2341 : _GEN_1751; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2814 = 2'h2 != last_proc_id ? _GEN_2342 : _GEN_1752; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2815 = 2'h2 != last_proc_id ? _GEN_2343 : _GEN_1753; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2816 = 2'h2 != last_proc_id ? _GEN_2344 : _GEN_1754; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2817 = 2'h2 != last_proc_id ? _GEN_2345 : _GEN_1755; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2818 = 2'h2 != last_proc_id ? _GEN_2346 : _GEN_1756; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2819 = 2'h2 != last_proc_id ? _GEN_2347 : _GEN_1757; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2820 = 2'h2 != last_proc_id ? _GEN_2348 : _GEN_1758; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2821 = 2'h2 != last_proc_id ? _GEN_2349 : _GEN_1759; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2822 = 2'h2 != last_proc_id ? _GEN_2350 : _GEN_1760; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2823 = 2'h2 != last_proc_id ? _GEN_2351 : _GEN_1761; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2824 = 2'h2 != last_proc_id ? _GEN_2352 : _GEN_1762; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2825 = 2'h2 != last_proc_id ? _GEN_2353 : _GEN_1763; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2826 = 2'h2 != last_proc_id ? _GEN_2354 : _GEN_1764; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2827 = 2'h2 != last_proc_id ? _GEN_2355 : _GEN_1765; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2828 = 2'h2 != last_proc_id ? _GEN_2356 : _GEN_1766; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2829 = 2'h2 != last_proc_id ? _GEN_2357 : _GEN_1767; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2830 = 2'h2 != last_proc_id ? _GEN_2358 : _GEN_1768; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2831 = 2'h2 != last_proc_id ? _GEN_2359 : _GEN_1769; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2832 = 2'h2 != last_proc_id ? _GEN_2360 : _GEN_1770; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2833 = 2'h2 != last_proc_id ? _GEN_2361 : _GEN_1771; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2834 = 2'h2 != last_proc_id ? _GEN_2362 : _GEN_1772; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2835 = 2'h2 != last_proc_id ? _GEN_2363 : _GEN_1773; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2836 = 2'h2 != last_proc_id ? _GEN_2364 : _GEN_1774; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2837 = 2'h2 != last_proc_id ? _GEN_2365 : _GEN_1775; // @[ipsa.scala 94:65]
  wire  _GEN_2838 = 2'h2 != last_proc_id ? _GEN_2366 : _GEN_1776; // @[ipsa.scala 94:65]
  wire  _GEN_2839 = 2'h2 != last_proc_id ? _GEN_2367 : _GEN_1777; // @[ipsa.scala 94:65]
  wire [1:0] _GEN_2840 = 2'h2 != last_proc_id ? _GEN_2368 : _GEN_1778; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2841 = 2'h2 != last_proc_id ? _GEN_2369 : _GEN_1779; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2842 = 2'h2 != last_proc_id ? _GEN_2370 : _GEN_1780; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2843 = 2'h2 != last_proc_id ? _GEN_2371 : _GEN_1781; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2844 = 2'h2 != last_proc_id ? _GEN_2372 : _GEN_1782; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2845 = 2'h2 != last_proc_id ? _GEN_2373 : _GEN_1783; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2846 = 2'h2 != last_proc_id ? _GEN_2374 : _GEN_1784; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2847 = 2'h2 != last_proc_id ? _GEN_2375 : _GEN_1785; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2848 = 2'h2 != last_proc_id ? _GEN_2376 : _GEN_1786; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2849 = 2'h2 != last_proc_id ? _GEN_2377 : _GEN_1787; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2850 = 2'h2 != last_proc_id ? _GEN_2378 : _GEN_1788; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2851 = 2'h2 != last_proc_id ? _GEN_2379 : _GEN_1789; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2852 = 2'h2 != last_proc_id ? _GEN_2380 : _GEN_1790; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2853 = 2'h2 != last_proc_id ? _GEN_2381 : _GEN_1791; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2854 = 2'h2 != last_proc_id ? _GEN_2382 : _GEN_1792; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2855 = 2'h2 != last_proc_id ? _GEN_2383 : _GEN_1793; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2856 = 2'h2 != last_proc_id ? _GEN_2384 : _GEN_1794; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2857 = 2'h2 != last_proc_id ? _GEN_2385 : _GEN_1795; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2858 = 2'h2 != last_proc_id ? _GEN_2386 : _GEN_1796; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2859 = 2'h2 != last_proc_id ? _GEN_2387 : _GEN_1797; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2860 = 2'h2 != last_proc_id ? _GEN_2388 : _GEN_1798; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2861 = 2'h2 != last_proc_id ? _GEN_2389 : _GEN_1799; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2862 = 2'h2 != last_proc_id ? _GEN_2390 : _GEN_1800; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2863 = 2'h2 != last_proc_id ? _GEN_2391 : _GEN_1801; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2864 = 2'h2 != last_proc_id ? _GEN_2392 : _GEN_1802; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2865 = 2'h2 != last_proc_id ? _GEN_2393 : _GEN_1803; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2866 = 2'h2 != last_proc_id ? _GEN_2394 : _GEN_1804; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2867 = 2'h2 != last_proc_id ? _GEN_2395 : _GEN_1805; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2868 = 2'h2 != last_proc_id ? _GEN_2396 : _GEN_1806; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2869 = 2'h2 != last_proc_id ? _GEN_2397 : _GEN_1807; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2870 = 2'h2 != last_proc_id ? _GEN_2398 : _GEN_1808; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2871 = 2'h2 != last_proc_id ? _GEN_2399 : _GEN_1809; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2872 = 2'h2 != last_proc_id ? _GEN_2400 : _GEN_1810; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2873 = 2'h2 != last_proc_id ? _GEN_2401 : _GEN_1811; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2874 = 2'h2 != last_proc_id ? _GEN_2402 : _GEN_1812; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2875 = 2'h2 != last_proc_id ? _GEN_2403 : _GEN_1813; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2876 = 2'h2 != last_proc_id ? _GEN_2404 : _GEN_1814; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2877 = 2'h2 != last_proc_id ? _GEN_2405 : _GEN_1815; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2878 = 2'h2 != last_proc_id ? _GEN_2406 : _GEN_1816; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2879 = 2'h2 != last_proc_id ? _GEN_2407 : _GEN_1817; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2880 = 2'h2 != last_proc_id ? _GEN_2408 : _GEN_1818; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2881 = 2'h2 != last_proc_id ? _GEN_2409 : _GEN_1819; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2882 = 2'h2 != last_proc_id ? _GEN_2410 : _GEN_1820; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2883 = 2'h2 != last_proc_id ? _GEN_2411 : _GEN_1821; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2884 = 2'h2 != last_proc_id ? _GEN_2412 : _GEN_1822; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2885 = 2'h2 != last_proc_id ? _GEN_2413 : _GEN_1823; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2886 = 2'h2 != last_proc_id ? _GEN_2414 : _GEN_1824; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2887 = 2'h2 != last_proc_id ? _GEN_2415 : _GEN_1825; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2888 = 2'h2 != last_proc_id ? _GEN_2416 : _GEN_1826; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2889 = 2'h2 != last_proc_id ? _GEN_2417 : _GEN_1827; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2890 = 2'h2 != last_proc_id ? _GEN_2418 : _GEN_1828; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2891 = 2'h2 != last_proc_id ? _GEN_2419 : _GEN_1829; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2892 = 2'h2 != last_proc_id ? _GEN_2420 : _GEN_1830; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2893 = 2'h2 != last_proc_id ? _GEN_2421 : _GEN_1831; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2894 = 2'h2 != last_proc_id ? _GEN_2422 : _GEN_1832; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2895 = 2'h2 != last_proc_id ? _GEN_2423 : _GEN_1833; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2896 = 2'h2 != last_proc_id ? _GEN_2424 : _GEN_1834; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2897 = 2'h2 != last_proc_id ? _GEN_2425 : _GEN_1835; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2898 = 2'h2 != last_proc_id ? _GEN_2426 : _GEN_1836; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2899 = 2'h2 != last_proc_id ? _GEN_2427 : _GEN_1837; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2900 = 2'h2 != last_proc_id ? _GEN_2428 : _GEN_1838; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2901 = 2'h2 != last_proc_id ? _GEN_2429 : _GEN_1839; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2902 = 2'h2 != last_proc_id ? _GEN_2430 : _GEN_1840; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2903 = 2'h2 != last_proc_id ? _GEN_2431 : _GEN_1841; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2904 = 2'h2 != last_proc_id ? _GEN_2432 : _GEN_1842; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2905 = 2'h2 != last_proc_id ? _GEN_2433 : _GEN_1843; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2906 = 2'h2 != last_proc_id ? _GEN_2434 : _GEN_1844; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2907 = 2'h2 != last_proc_id ? _GEN_2435 : _GEN_1845; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2908 = 2'h2 != last_proc_id ? _GEN_2436 : _GEN_1846; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2909 = 2'h2 != last_proc_id ? _GEN_2437 : _GEN_1847; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2910 = 2'h2 != last_proc_id ? _GEN_2438 : _GEN_1848; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2911 = 2'h2 != last_proc_id ? _GEN_2439 : _GEN_1849; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2912 = 2'h2 != last_proc_id ? _GEN_2440 : _GEN_1850; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2913 = 2'h2 != last_proc_id ? _GEN_2441 : _GEN_1851; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2914 = 2'h2 != last_proc_id ? _GEN_2442 : _GEN_1852; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2915 = 2'h2 != last_proc_id ? _GEN_2443 : _GEN_1853; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2916 = 2'h2 != last_proc_id ? _GEN_2444 : _GEN_1854; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2917 = 2'h2 != last_proc_id ? _GEN_2445 : _GEN_1855; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2918 = 2'h2 != last_proc_id ? _GEN_2446 : _GEN_1856; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2919 = 2'h2 != last_proc_id ? _GEN_2447 : _GEN_1857; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2920 = 2'h2 != last_proc_id ? _GEN_2448 : _GEN_1858; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2921 = 2'h2 != last_proc_id ? _GEN_2449 : _GEN_1859; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2922 = 2'h2 != last_proc_id ? _GEN_2450 : _GEN_1860; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2923 = 2'h2 != last_proc_id ? _GEN_2451 : _GEN_1861; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2924 = 2'h2 != last_proc_id ? _GEN_2452 : _GEN_1862; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2925 = 2'h2 != last_proc_id ? _GEN_2453 : _GEN_1863; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2926 = 2'h2 != last_proc_id ? _GEN_2454 : _GEN_1864; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2927 = 2'h2 != last_proc_id ? _GEN_2455 : _GEN_1865; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2928 = 2'h2 != last_proc_id ? _GEN_2456 : _GEN_1866; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2929 = 2'h2 != last_proc_id ? _GEN_2457 : _GEN_1867; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2930 = 2'h2 != last_proc_id ? _GEN_2458 : _GEN_1868; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2931 = 2'h2 != last_proc_id ? _GEN_2459 : _GEN_1869; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2932 = 2'h2 != last_proc_id ? _GEN_2460 : _GEN_1870; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2933 = 2'h2 != last_proc_id ? _GEN_2461 : _GEN_1871; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2934 = 2'h2 != last_proc_id ? _GEN_2462 : _GEN_1872; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2935 = 2'h2 != last_proc_id ? _GEN_2463 : _GEN_1873; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2936 = 2'h2 != last_proc_id ? _GEN_2464 : _GEN_1874; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2937 = 2'h2 != last_proc_id ? _GEN_2465 : _GEN_1875; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2938 = 2'h2 != last_proc_id ? _GEN_2466 : _GEN_1876; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2939 = 2'h2 != last_proc_id ? _GEN_2467 : _GEN_1877; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2940 = 2'h2 != last_proc_id ? _GEN_2468 : _GEN_1878; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2941 = 2'h2 != last_proc_id ? _GEN_2469 : _GEN_1879; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2942 = 2'h2 != last_proc_id ? _GEN_2470 : _GEN_1880; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2943 = 2'h2 != last_proc_id ? _GEN_2471 : _GEN_1881; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2944 = 2'h2 != last_proc_id ? _GEN_2472 : _GEN_1882; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2945 = 2'h2 != last_proc_id ? _GEN_2473 : _GEN_1883; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2946 = 2'h2 != last_proc_id ? _GEN_2474 : _GEN_1884; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2947 = 2'h2 != last_proc_id ? _GEN_2475 : _GEN_1885; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2948 = 2'h2 != last_proc_id ? _GEN_2476 : _GEN_1886; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2949 = 2'h2 != last_proc_id ? _GEN_2477 : _GEN_1887; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2950 = 2'h2 != last_proc_id ? _GEN_2478 : _GEN_1888; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2951 = 2'h2 != last_proc_id ? _GEN_2479 : _GEN_1889; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2952 = 2'h2 != last_proc_id ? _GEN_2480 : _GEN_1890; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2953 = 2'h2 != last_proc_id ? _GEN_2481 : _GEN_1891; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2954 = 2'h2 != last_proc_id ? _GEN_2482 : _GEN_1892; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2955 = 2'h2 != last_proc_id ? _GEN_2483 : _GEN_1893; // @[ipsa.scala 94:65]
  wire  _GEN_2956 = 2'h2 != last_proc_id ? _GEN_2484 : _GEN_1894; // @[ipsa.scala 94:65]
  wire  _GEN_2957 = 2'h2 != last_proc_id ? _GEN_2485 : _GEN_1895; // @[ipsa.scala 94:65]
  wire [1:0] _GEN_2958 = 2'h2 != last_proc_id ? _GEN_2486 : _GEN_1896; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2959 = 2'h2 != last_proc_id ? _GEN_2487 : _GEN_1897; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2960 = 2'h2 != last_proc_id ? _GEN_2488 : _GEN_1898; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2961 = 2'h2 != last_proc_id ? _GEN_2489 : _GEN_1899; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2962 = 2'h2 != last_proc_id ? _GEN_2490 : _GEN_1900; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2963 = 2'h2 != last_proc_id ? _GEN_2491 : _GEN_1901; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2964 = 2'h2 != last_proc_id ? _GEN_2492 : _GEN_1902; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2965 = 2'h2 != last_proc_id ? _GEN_2493 : _GEN_1903; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2966 = 2'h2 != last_proc_id ? _GEN_2494 : _GEN_1904; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2967 = 2'h2 != last_proc_id ? _GEN_2495 : _GEN_1905; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2968 = 2'h2 != last_proc_id ? _GEN_2496 : _GEN_1906; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2969 = 2'h2 != last_proc_id ? _GEN_2497 : _GEN_1907; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2970 = 2'h2 != last_proc_id ? _GEN_2498 : _GEN_1908; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2971 = 2'h2 != last_proc_id ? _GEN_2499 : _GEN_1909; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2972 = 2'h2 != last_proc_id ? _GEN_2500 : _GEN_1910; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2973 = 2'h2 != last_proc_id ? _GEN_2501 : _GEN_1911; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2974 = 2'h2 != last_proc_id ? _GEN_2502 : _GEN_1912; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2975 = 2'h2 != last_proc_id ? _GEN_2503 : _GEN_1913; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2976 = 2'h2 != last_proc_id ? _GEN_2504 : _GEN_1914; // @[ipsa.scala 94:65]
  wire [15:0] _GEN_2977 = 2'h2 != last_proc_id ? _GEN_2505 : _GEN_1915; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2978 = 2'h2 != last_proc_id ? _GEN_2506 : _GEN_1916; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2979 = 2'h2 != last_proc_id ? _GEN_2507 : _GEN_1917; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2980 = 2'h2 != last_proc_id ? _GEN_2508 : _GEN_1918; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2981 = 2'h2 != last_proc_id ? _GEN_2509 : _GEN_1919; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2982 = 2'h2 != last_proc_id ? _GEN_2510 : _GEN_1920; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2983 = 2'h2 != last_proc_id ? _GEN_2511 : _GEN_1921; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2984 = 2'h2 != last_proc_id ? _GEN_2512 : _GEN_1922; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2985 = 2'h2 != last_proc_id ? _GEN_2513 : _GEN_1923; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2986 = 2'h2 != last_proc_id ? _GEN_2514 : _GEN_1924; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2987 = 2'h2 != last_proc_id ? _GEN_2515 : _GEN_1925; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2988 = 2'h2 != last_proc_id ? _GEN_2516 : _GEN_1926; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2989 = 2'h2 != last_proc_id ? _GEN_2517 : _GEN_1927; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2990 = 2'h2 != last_proc_id ? _GEN_2518 : _GEN_1928; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2991 = 2'h2 != last_proc_id ? _GEN_2519 : _GEN_1929; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2992 = 2'h2 != last_proc_id ? _GEN_2520 : _GEN_1930; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2993 = 2'h2 != last_proc_id ? _GEN_2521 : _GEN_1931; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2994 = 2'h2 != last_proc_id ? _GEN_2522 : _GEN_1932; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2995 = 2'h2 != last_proc_id ? _GEN_2523 : _GEN_1933; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2996 = 2'h2 != last_proc_id ? _GEN_2524 : _GEN_1934; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2997 = 2'h2 != last_proc_id ? _GEN_2525 : _GEN_1935; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2998 = 2'h2 != last_proc_id ? _GEN_2526 : _GEN_1936; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_2999 = 2'h2 != last_proc_id ? _GEN_2527 : _GEN_1937; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3000 = 2'h2 != last_proc_id ? _GEN_2528 : _GEN_1938; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3001 = 2'h2 != last_proc_id ? _GEN_2529 : _GEN_1939; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3002 = 2'h2 != last_proc_id ? _GEN_2530 : _GEN_1940; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3003 = 2'h2 != last_proc_id ? _GEN_2531 : _GEN_1941; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3004 = 2'h2 != last_proc_id ? _GEN_2532 : _GEN_1942; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3005 = 2'h2 != last_proc_id ? _GEN_2533 : _GEN_1943; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3006 = 2'h2 != last_proc_id ? _GEN_2534 : _GEN_1944; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3007 = 2'h2 != last_proc_id ? _GEN_2535 : _GEN_1945; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3008 = 2'h2 != last_proc_id ? _GEN_2536 : _GEN_1946; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3009 = 2'h2 != last_proc_id ? _GEN_2537 : _GEN_1947; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3010 = 2'h2 != last_proc_id ? _GEN_2538 : _GEN_1948; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3011 = 2'h2 != last_proc_id ? _GEN_2539 : _GEN_1949; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3012 = 2'h2 != last_proc_id ? _GEN_2540 : _GEN_1950; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3013 = 2'h2 != last_proc_id ? _GEN_2541 : _GEN_1951; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3014 = 2'h2 != last_proc_id ? _GEN_2542 : _GEN_1952; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3015 = 2'h2 != last_proc_id ? _GEN_2543 : _GEN_1953; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3016 = 2'h2 != last_proc_id ? _GEN_2544 : _GEN_1954; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3017 = 2'h2 != last_proc_id ? _GEN_2545 : _GEN_1955; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3018 = 2'h2 != last_proc_id ? _GEN_2546 : _GEN_1956; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3019 = 2'h2 != last_proc_id ? _GEN_2547 : _GEN_1957; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3020 = 2'h2 != last_proc_id ? _GEN_2548 : _GEN_1958; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3021 = 2'h2 != last_proc_id ? _GEN_2549 : _GEN_1959; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3022 = 2'h2 != last_proc_id ? _GEN_2550 : _GEN_1960; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3023 = 2'h2 != last_proc_id ? _GEN_2551 : _GEN_1961; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3024 = 2'h2 != last_proc_id ? _GEN_2552 : _GEN_1962; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3025 = 2'h2 != last_proc_id ? _GEN_2553 : _GEN_1963; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3026 = 2'h2 != last_proc_id ? _GEN_2554 : _GEN_1964; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3027 = 2'h2 != last_proc_id ? _GEN_2555 : _GEN_1965; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3028 = 2'h2 != last_proc_id ? _GEN_2556 : _GEN_1966; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3029 = 2'h2 != last_proc_id ? _GEN_2557 : _GEN_1967; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3030 = 2'h2 != last_proc_id ? _GEN_2558 : _GEN_1968; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3031 = 2'h2 != last_proc_id ? _GEN_2559 : _GEN_1969; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3032 = 2'h2 != last_proc_id ? _GEN_2560 : _GEN_1970; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3033 = 2'h2 != last_proc_id ? _GEN_2561 : _GEN_1971; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3034 = 2'h2 != last_proc_id ? _GEN_2562 : _GEN_1972; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3035 = 2'h2 != last_proc_id ? _GEN_2563 : _GEN_1973; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3036 = 2'h2 != last_proc_id ? _GEN_2564 : _GEN_1974; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3037 = 2'h2 != last_proc_id ? _GEN_2565 : _GEN_1975; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3038 = 2'h2 != last_proc_id ? _GEN_2566 : _GEN_1976; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3039 = 2'h2 != last_proc_id ? _GEN_2567 : _GEN_1977; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3040 = 2'h2 != last_proc_id ? _GEN_2568 : _GEN_1978; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3041 = 2'h2 != last_proc_id ? _GEN_2569 : _GEN_1979; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3042 = 2'h2 != last_proc_id ? _GEN_2570 : _GEN_1980; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3043 = 2'h2 != last_proc_id ? _GEN_2571 : _GEN_1981; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3044 = 2'h2 != last_proc_id ? _GEN_2572 : _GEN_1982; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3045 = 2'h2 != last_proc_id ? _GEN_2573 : _GEN_1983; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3046 = 2'h2 != last_proc_id ? _GEN_2574 : _GEN_1984; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3047 = 2'h2 != last_proc_id ? _GEN_2575 : _GEN_1985; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3048 = 2'h2 != last_proc_id ? _GEN_2576 : _GEN_1986; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3049 = 2'h2 != last_proc_id ? _GEN_2577 : _GEN_1987; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3050 = 2'h2 != last_proc_id ? _GEN_2578 : _GEN_1988; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3051 = 2'h2 != last_proc_id ? _GEN_2579 : _GEN_1989; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3052 = 2'h2 != last_proc_id ? _GEN_2580 : _GEN_1990; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3053 = 2'h2 != last_proc_id ? _GEN_2581 : _GEN_1991; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3054 = 2'h2 != last_proc_id ? _GEN_2582 : _GEN_1992; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3055 = 2'h2 != last_proc_id ? _GEN_2583 : _GEN_1993; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3056 = 2'h2 != last_proc_id ? _GEN_2584 : _GEN_1994; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3057 = 2'h2 != last_proc_id ? _GEN_2585 : _GEN_1995; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3058 = 2'h2 != last_proc_id ? _GEN_2586 : _GEN_1996; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3059 = 2'h2 != last_proc_id ? _GEN_2587 : _GEN_1997; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3060 = 2'h2 != last_proc_id ? _GEN_2588 : _GEN_1998; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3061 = 2'h2 != last_proc_id ? _GEN_2589 : _GEN_1999; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3062 = 2'h2 != last_proc_id ? _GEN_2590 : _GEN_2000; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3063 = 2'h2 != last_proc_id ? _GEN_2591 : _GEN_2001; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3064 = 2'h2 != last_proc_id ? _GEN_2592 : _GEN_2002; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3065 = 2'h2 != last_proc_id ? _GEN_2593 : _GEN_2003; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3066 = 2'h2 != last_proc_id ? _GEN_2594 : _GEN_2004; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3067 = 2'h2 != last_proc_id ? _GEN_2595 : _GEN_2005; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3068 = 2'h2 != last_proc_id ? _GEN_2596 : _GEN_2006; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3069 = 2'h2 != last_proc_id ? _GEN_2597 : _GEN_2007; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3070 = 2'h2 != last_proc_id ? _GEN_2598 : _GEN_2008; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3071 = 2'h2 != last_proc_id ? _GEN_2599 : _GEN_2009; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3072 = 2'h2 != last_proc_id ? _GEN_2600 : _GEN_2010; // @[ipsa.scala 94:65]
  wire [7:0] _GEN_3073 = 2'h2 != last_proc_id ? _GEN_2601 : _GEN_2011; // @[ipsa.scala 94:65]
  wire  _GEN_3074 = 2'h2 != last_proc_id ? _GEN_2012 : trans_2_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire  _GEN_3075 = 2'h2 != last_proc_id ? _GEN_2013 : trans_2_io_pipe_phv_out_next_config_id; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [1:0] _GEN_3076 = 2'h2 != last_proc_id ? _GEN_2014 : trans_2_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_3077 = 2'h2 != last_proc_id ? _GEN_2015 : trans_2_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3078 = 2'h2 != last_proc_id ? _GEN_2016 : trans_2_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3079 = 2'h2 != last_proc_id ? _GEN_2017 : trans_2_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_3080 = 2'h2 != last_proc_id ? _GEN_2018 : trans_2_io_pipe_phv_out_header_0; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_3081 = 2'h2 != last_proc_id ? _GEN_2019 : trans_2_io_pipe_phv_out_header_1; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_3082 = 2'h2 != last_proc_id ? _GEN_2020 : trans_2_io_pipe_phv_out_header_2; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_3083 = 2'h2 != last_proc_id ? _GEN_2021 : trans_2_io_pipe_phv_out_header_3; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_3084 = 2'h2 != last_proc_id ? _GEN_2022 : trans_2_io_pipe_phv_out_header_4; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_3085 = 2'h2 != last_proc_id ? _GEN_2023 : trans_2_io_pipe_phv_out_header_5; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_3086 = 2'h2 != last_proc_id ? _GEN_2024 : trans_2_io_pipe_phv_out_header_6; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_3087 = 2'h2 != last_proc_id ? _GEN_2025 : trans_2_io_pipe_phv_out_header_7; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_3088 = 2'h2 != last_proc_id ? _GEN_2026 : trans_2_io_pipe_phv_out_header_8; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_3089 = 2'h2 != last_proc_id ? _GEN_2027 : trans_2_io_pipe_phv_out_header_9; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_3090 = 2'h2 != last_proc_id ? _GEN_2028 : trans_2_io_pipe_phv_out_header_10; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_3091 = 2'h2 != last_proc_id ? _GEN_2029 : trans_2_io_pipe_phv_out_header_11; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_3092 = 2'h2 != last_proc_id ? _GEN_2030 : trans_2_io_pipe_phv_out_header_12; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_3093 = 2'h2 != last_proc_id ? _GEN_2031 : trans_2_io_pipe_phv_out_header_13; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_3094 = 2'h2 != last_proc_id ? _GEN_2032 : trans_2_io_pipe_phv_out_header_14; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [15:0] _GEN_3095 = 2'h2 != last_proc_id ? _GEN_2033 : trans_2_io_pipe_phv_out_header_15; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3096 = 2'h2 != last_proc_id ? _GEN_2034 : trans_2_io_pipe_phv_out_data_0; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3097 = 2'h2 != last_proc_id ? _GEN_2035 : trans_2_io_pipe_phv_out_data_1; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3098 = 2'h2 != last_proc_id ? _GEN_2036 : trans_2_io_pipe_phv_out_data_2; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3099 = 2'h2 != last_proc_id ? _GEN_2037 : trans_2_io_pipe_phv_out_data_3; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3100 = 2'h2 != last_proc_id ? _GEN_2038 : trans_2_io_pipe_phv_out_data_4; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3101 = 2'h2 != last_proc_id ? _GEN_2039 : trans_2_io_pipe_phv_out_data_5; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3102 = 2'h2 != last_proc_id ? _GEN_2040 : trans_2_io_pipe_phv_out_data_6; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3103 = 2'h2 != last_proc_id ? _GEN_2041 : trans_2_io_pipe_phv_out_data_7; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3104 = 2'h2 != last_proc_id ? _GEN_2042 : trans_2_io_pipe_phv_out_data_8; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3105 = 2'h2 != last_proc_id ? _GEN_2043 : trans_2_io_pipe_phv_out_data_9; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3106 = 2'h2 != last_proc_id ? _GEN_2044 : trans_2_io_pipe_phv_out_data_10; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3107 = 2'h2 != last_proc_id ? _GEN_2045 : trans_2_io_pipe_phv_out_data_11; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3108 = 2'h2 != last_proc_id ? _GEN_2046 : trans_2_io_pipe_phv_out_data_12; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3109 = 2'h2 != last_proc_id ? _GEN_2047 : trans_2_io_pipe_phv_out_data_13; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3110 = 2'h2 != last_proc_id ? _GEN_2048 : trans_2_io_pipe_phv_out_data_14; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3111 = 2'h2 != last_proc_id ? _GEN_2049 : trans_2_io_pipe_phv_out_data_15; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3112 = 2'h2 != last_proc_id ? _GEN_2050 : trans_2_io_pipe_phv_out_data_16; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3113 = 2'h2 != last_proc_id ? _GEN_2051 : trans_2_io_pipe_phv_out_data_17; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3114 = 2'h2 != last_proc_id ? _GEN_2052 : trans_2_io_pipe_phv_out_data_18; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3115 = 2'h2 != last_proc_id ? _GEN_2053 : trans_2_io_pipe_phv_out_data_19; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3116 = 2'h2 != last_proc_id ? _GEN_2054 : trans_2_io_pipe_phv_out_data_20; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3117 = 2'h2 != last_proc_id ? _GEN_2055 : trans_2_io_pipe_phv_out_data_21; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3118 = 2'h2 != last_proc_id ? _GEN_2056 : trans_2_io_pipe_phv_out_data_22; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3119 = 2'h2 != last_proc_id ? _GEN_2057 : trans_2_io_pipe_phv_out_data_23; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3120 = 2'h2 != last_proc_id ? _GEN_2058 : trans_2_io_pipe_phv_out_data_24; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3121 = 2'h2 != last_proc_id ? _GEN_2059 : trans_2_io_pipe_phv_out_data_25; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3122 = 2'h2 != last_proc_id ? _GEN_2060 : trans_2_io_pipe_phv_out_data_26; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3123 = 2'h2 != last_proc_id ? _GEN_2061 : trans_2_io_pipe_phv_out_data_27; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3124 = 2'h2 != last_proc_id ? _GEN_2062 : trans_2_io_pipe_phv_out_data_28; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3125 = 2'h2 != last_proc_id ? _GEN_2063 : trans_2_io_pipe_phv_out_data_29; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3126 = 2'h2 != last_proc_id ? _GEN_2064 : trans_2_io_pipe_phv_out_data_30; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3127 = 2'h2 != last_proc_id ? _GEN_2065 : trans_2_io_pipe_phv_out_data_31; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3128 = 2'h2 != last_proc_id ? _GEN_2066 : trans_2_io_pipe_phv_out_data_32; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3129 = 2'h2 != last_proc_id ? _GEN_2067 : trans_2_io_pipe_phv_out_data_33; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3130 = 2'h2 != last_proc_id ? _GEN_2068 : trans_2_io_pipe_phv_out_data_34; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3131 = 2'h2 != last_proc_id ? _GEN_2069 : trans_2_io_pipe_phv_out_data_35; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3132 = 2'h2 != last_proc_id ? _GEN_2070 : trans_2_io_pipe_phv_out_data_36; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3133 = 2'h2 != last_proc_id ? _GEN_2071 : trans_2_io_pipe_phv_out_data_37; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3134 = 2'h2 != last_proc_id ? _GEN_2072 : trans_2_io_pipe_phv_out_data_38; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3135 = 2'h2 != last_proc_id ? _GEN_2073 : trans_2_io_pipe_phv_out_data_39; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3136 = 2'h2 != last_proc_id ? _GEN_2074 : trans_2_io_pipe_phv_out_data_40; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3137 = 2'h2 != last_proc_id ? _GEN_2075 : trans_2_io_pipe_phv_out_data_41; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3138 = 2'h2 != last_proc_id ? _GEN_2076 : trans_2_io_pipe_phv_out_data_42; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3139 = 2'h2 != last_proc_id ? _GEN_2077 : trans_2_io_pipe_phv_out_data_43; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3140 = 2'h2 != last_proc_id ? _GEN_2078 : trans_2_io_pipe_phv_out_data_44; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3141 = 2'h2 != last_proc_id ? _GEN_2079 : trans_2_io_pipe_phv_out_data_45; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3142 = 2'h2 != last_proc_id ? _GEN_2080 : trans_2_io_pipe_phv_out_data_46; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3143 = 2'h2 != last_proc_id ? _GEN_2081 : trans_2_io_pipe_phv_out_data_47; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3144 = 2'h2 != last_proc_id ? _GEN_2082 : trans_2_io_pipe_phv_out_data_48; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3145 = 2'h2 != last_proc_id ? _GEN_2083 : trans_2_io_pipe_phv_out_data_49; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3146 = 2'h2 != last_proc_id ? _GEN_2084 : trans_2_io_pipe_phv_out_data_50; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3147 = 2'h2 != last_proc_id ? _GEN_2085 : trans_2_io_pipe_phv_out_data_51; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3148 = 2'h2 != last_proc_id ? _GEN_2086 : trans_2_io_pipe_phv_out_data_52; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3149 = 2'h2 != last_proc_id ? _GEN_2087 : trans_2_io_pipe_phv_out_data_53; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3150 = 2'h2 != last_proc_id ? _GEN_2088 : trans_2_io_pipe_phv_out_data_54; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3151 = 2'h2 != last_proc_id ? _GEN_2089 : trans_2_io_pipe_phv_out_data_55; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3152 = 2'h2 != last_proc_id ? _GEN_2090 : trans_2_io_pipe_phv_out_data_56; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3153 = 2'h2 != last_proc_id ? _GEN_2091 : trans_2_io_pipe_phv_out_data_57; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3154 = 2'h2 != last_proc_id ? _GEN_2092 : trans_2_io_pipe_phv_out_data_58; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3155 = 2'h2 != last_proc_id ? _GEN_2093 : trans_2_io_pipe_phv_out_data_59; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3156 = 2'h2 != last_proc_id ? _GEN_2094 : trans_2_io_pipe_phv_out_data_60; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3157 = 2'h2 != last_proc_id ? _GEN_2095 : trans_2_io_pipe_phv_out_data_61; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3158 = 2'h2 != last_proc_id ? _GEN_2096 : trans_2_io_pipe_phv_out_data_62; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3159 = 2'h2 != last_proc_id ? _GEN_2097 : trans_2_io_pipe_phv_out_data_63; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3160 = 2'h2 != last_proc_id ? _GEN_2098 : trans_2_io_pipe_phv_out_data_64; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3161 = 2'h2 != last_proc_id ? _GEN_2099 : trans_2_io_pipe_phv_out_data_65; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3162 = 2'h2 != last_proc_id ? _GEN_2100 : trans_2_io_pipe_phv_out_data_66; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3163 = 2'h2 != last_proc_id ? _GEN_2101 : trans_2_io_pipe_phv_out_data_67; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3164 = 2'h2 != last_proc_id ? _GEN_2102 : trans_2_io_pipe_phv_out_data_68; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3165 = 2'h2 != last_proc_id ? _GEN_2103 : trans_2_io_pipe_phv_out_data_69; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3166 = 2'h2 != last_proc_id ? _GEN_2104 : trans_2_io_pipe_phv_out_data_70; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3167 = 2'h2 != last_proc_id ? _GEN_2105 : trans_2_io_pipe_phv_out_data_71; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3168 = 2'h2 != last_proc_id ? _GEN_2106 : trans_2_io_pipe_phv_out_data_72; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3169 = 2'h2 != last_proc_id ? _GEN_2107 : trans_2_io_pipe_phv_out_data_73; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3170 = 2'h2 != last_proc_id ? _GEN_2108 : trans_2_io_pipe_phv_out_data_74; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3171 = 2'h2 != last_proc_id ? _GEN_2109 : trans_2_io_pipe_phv_out_data_75; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3172 = 2'h2 != last_proc_id ? _GEN_2110 : trans_2_io_pipe_phv_out_data_76; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3173 = 2'h2 != last_proc_id ? _GEN_2111 : trans_2_io_pipe_phv_out_data_77; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3174 = 2'h2 != last_proc_id ? _GEN_2112 : trans_2_io_pipe_phv_out_data_78; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3175 = 2'h2 != last_proc_id ? _GEN_2113 : trans_2_io_pipe_phv_out_data_79; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3176 = 2'h2 != last_proc_id ? _GEN_2114 : trans_2_io_pipe_phv_out_data_80; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3177 = 2'h2 != last_proc_id ? _GEN_2115 : trans_2_io_pipe_phv_out_data_81; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3178 = 2'h2 != last_proc_id ? _GEN_2116 : trans_2_io_pipe_phv_out_data_82; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3179 = 2'h2 != last_proc_id ? _GEN_2117 : trans_2_io_pipe_phv_out_data_83; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3180 = 2'h2 != last_proc_id ? _GEN_2118 : trans_2_io_pipe_phv_out_data_84; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3181 = 2'h2 != last_proc_id ? _GEN_2119 : trans_2_io_pipe_phv_out_data_85; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3182 = 2'h2 != last_proc_id ? _GEN_2120 : trans_2_io_pipe_phv_out_data_86; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3183 = 2'h2 != last_proc_id ? _GEN_2121 : trans_2_io_pipe_phv_out_data_87; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3184 = 2'h2 != last_proc_id ? _GEN_2122 : trans_2_io_pipe_phv_out_data_88; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3185 = 2'h2 != last_proc_id ? _GEN_2123 : trans_2_io_pipe_phv_out_data_89; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3186 = 2'h2 != last_proc_id ? _GEN_2124 : trans_2_io_pipe_phv_out_data_90; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3187 = 2'h2 != last_proc_id ? _GEN_2125 : trans_2_io_pipe_phv_out_data_91; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3188 = 2'h2 != last_proc_id ? _GEN_2126 : trans_2_io_pipe_phv_out_data_92; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3189 = 2'h2 != last_proc_id ? _GEN_2127 : trans_2_io_pipe_phv_out_data_93; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3190 = 2'h2 != last_proc_id ? _GEN_2128 : trans_2_io_pipe_phv_out_data_94; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire [7:0] _GEN_3191 = 2'h2 != last_proc_id ? _GEN_2129 : trans_2_io_pipe_phv_out_data_95; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  wire  _GEN_3192 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_is_valid_processor : _GEN_2602; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire  _GEN_3193 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_next_config_id : _GEN_2603; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [1:0] _GEN_3194 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_next_processor_id : _GEN_2604; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3195 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_parse_transition_field : _GEN_2605; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3196 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_parse_current_offset : _GEN_2606; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3197 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_parse_current_state : _GEN_2607; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3198 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_0 : _GEN_2608; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3199 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_1 : _GEN_2609; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3200 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_2 : _GEN_2610; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3201 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_3 : _GEN_2611; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3202 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_4 : _GEN_2612; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3203 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_5 : _GEN_2613; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3204 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_6 : _GEN_2614; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3205 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_7 : _GEN_2615; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3206 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_8 : _GEN_2616; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3207 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_9 : _GEN_2617; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3208 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_10 : _GEN_2618; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3209 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_11 : _GEN_2619; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3210 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_12 : _GEN_2620; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3211 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_13 : _GEN_2621; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3212 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_14 : _GEN_2622; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3213 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_15 : _GEN_2623; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3214 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_0 : _GEN_2624; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3215 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_1 : _GEN_2625; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3216 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_2 : _GEN_2626; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3217 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_3 : _GEN_2627; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3218 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_4 : _GEN_2628; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3219 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_5 : _GEN_2629; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3220 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_6 : _GEN_2630; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3221 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_7 : _GEN_2631; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3222 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_8 : _GEN_2632; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3223 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_9 : _GEN_2633; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3224 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_10 : _GEN_2634; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3225 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_11 : _GEN_2635; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3226 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_12 : _GEN_2636; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3227 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_13 : _GEN_2637; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3228 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_14 : _GEN_2638; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3229 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_15 : _GEN_2639; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3230 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_16 : _GEN_2640; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3231 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_17 : _GEN_2641; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3232 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_18 : _GEN_2642; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3233 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_19 : _GEN_2643; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3234 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_20 : _GEN_2644; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3235 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_21 : _GEN_2645; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3236 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_22 : _GEN_2646; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3237 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_23 : _GEN_2647; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3238 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_24 : _GEN_2648; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3239 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_25 : _GEN_2649; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3240 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_26 : _GEN_2650; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3241 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_27 : _GEN_2651; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3242 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_28 : _GEN_2652; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3243 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_29 : _GEN_2653; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3244 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_30 : _GEN_2654; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3245 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_31 : _GEN_2655; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3246 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_32 : _GEN_2656; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3247 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_33 : _GEN_2657; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3248 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_34 : _GEN_2658; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3249 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_35 : _GEN_2659; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3250 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_36 : _GEN_2660; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3251 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_37 : _GEN_2661; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3252 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_38 : _GEN_2662; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3253 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_39 : _GEN_2663; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3254 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_40 : _GEN_2664; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3255 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_41 : _GEN_2665; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3256 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_42 : _GEN_2666; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3257 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_43 : _GEN_2667; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3258 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_44 : _GEN_2668; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3259 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_45 : _GEN_2669; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3260 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_46 : _GEN_2670; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3261 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_47 : _GEN_2671; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3262 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_48 : _GEN_2672; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3263 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_49 : _GEN_2673; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3264 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_50 : _GEN_2674; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3265 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_51 : _GEN_2675; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3266 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_52 : _GEN_2676; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3267 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_53 : _GEN_2677; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3268 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_54 : _GEN_2678; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3269 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_55 : _GEN_2679; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3270 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_56 : _GEN_2680; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3271 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_57 : _GEN_2681; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3272 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_58 : _GEN_2682; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3273 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_59 : _GEN_2683; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3274 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_60 : _GEN_2684; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3275 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_61 : _GEN_2685; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3276 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_62 : _GEN_2686; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3277 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_63 : _GEN_2687; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3278 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_64 : _GEN_2688; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3279 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_65 : _GEN_2689; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3280 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_66 : _GEN_2690; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3281 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_67 : _GEN_2691; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3282 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_68 : _GEN_2692; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3283 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_69 : _GEN_2693; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3284 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_70 : _GEN_2694; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3285 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_71 : _GEN_2695; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3286 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_72 : _GEN_2696; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3287 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_73 : _GEN_2697; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3288 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_74 : _GEN_2698; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3289 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_75 : _GEN_2699; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3290 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_76 : _GEN_2700; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3291 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_77 : _GEN_2701; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3292 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_78 : _GEN_2702; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3293 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_79 : _GEN_2703; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3294 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_80 : _GEN_2704; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3295 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_81 : _GEN_2705; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3296 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_82 : _GEN_2706; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3297 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_83 : _GEN_2707; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3298 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_84 : _GEN_2708; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3299 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_85 : _GEN_2709; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3300 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_86 : _GEN_2710; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3301 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_87 : _GEN_2711; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3302 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_88 : _GEN_2712; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3303 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_89 : _GEN_2713; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3304 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_90 : _GEN_2714; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3305 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_91 : _GEN_2715; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3306 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_92 : _GEN_2716; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3307 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_93 : _GEN_2717; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3308 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_94 : _GEN_2718; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3309 = 2'h0 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_95 : _GEN_2719; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire  _GEN_3310 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_is_valid_processor : _GEN_2720; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire  _GEN_3311 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_next_config_id : _GEN_2721; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [1:0] _GEN_3312 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_next_processor_id : _GEN_2722; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3313 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_parse_transition_field : _GEN_2723; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3314 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_parse_current_offset : _GEN_2724; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3315 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_parse_current_state : _GEN_2725; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3316 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_0 : _GEN_2726; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3317 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_1 : _GEN_2727; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3318 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_2 : _GEN_2728; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3319 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_3 : _GEN_2729; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3320 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_4 : _GEN_2730; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3321 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_5 : _GEN_2731; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3322 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_6 : _GEN_2732; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3323 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_7 : _GEN_2733; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3324 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_8 : _GEN_2734; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3325 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_9 : _GEN_2735; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3326 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_10 : _GEN_2736; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3327 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_11 : _GEN_2737; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3328 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_12 : _GEN_2738; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3329 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_13 : _GEN_2739; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3330 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_14 : _GEN_2740; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3331 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_15 : _GEN_2741; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3332 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_0 : _GEN_2742; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3333 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_1 : _GEN_2743; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3334 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_2 : _GEN_2744; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3335 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_3 : _GEN_2745; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3336 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_4 : _GEN_2746; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3337 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_5 : _GEN_2747; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3338 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_6 : _GEN_2748; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3339 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_7 : _GEN_2749; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3340 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_8 : _GEN_2750; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3341 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_9 : _GEN_2751; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3342 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_10 : _GEN_2752; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3343 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_11 : _GEN_2753; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3344 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_12 : _GEN_2754; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3345 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_13 : _GEN_2755; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3346 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_14 : _GEN_2756; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3347 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_15 : _GEN_2757; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3348 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_16 : _GEN_2758; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3349 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_17 : _GEN_2759; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3350 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_18 : _GEN_2760; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3351 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_19 : _GEN_2761; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3352 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_20 : _GEN_2762; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3353 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_21 : _GEN_2763; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3354 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_22 : _GEN_2764; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3355 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_23 : _GEN_2765; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3356 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_24 : _GEN_2766; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3357 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_25 : _GEN_2767; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3358 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_26 : _GEN_2768; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3359 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_27 : _GEN_2769; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3360 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_28 : _GEN_2770; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3361 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_29 : _GEN_2771; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3362 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_30 : _GEN_2772; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3363 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_31 : _GEN_2773; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3364 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_32 : _GEN_2774; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3365 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_33 : _GEN_2775; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3366 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_34 : _GEN_2776; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3367 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_35 : _GEN_2777; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3368 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_36 : _GEN_2778; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3369 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_37 : _GEN_2779; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3370 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_38 : _GEN_2780; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3371 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_39 : _GEN_2781; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3372 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_40 : _GEN_2782; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3373 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_41 : _GEN_2783; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3374 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_42 : _GEN_2784; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3375 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_43 : _GEN_2785; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3376 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_44 : _GEN_2786; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3377 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_45 : _GEN_2787; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3378 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_46 : _GEN_2788; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3379 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_47 : _GEN_2789; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3380 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_48 : _GEN_2790; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3381 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_49 : _GEN_2791; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3382 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_50 : _GEN_2792; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3383 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_51 : _GEN_2793; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3384 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_52 : _GEN_2794; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3385 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_53 : _GEN_2795; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3386 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_54 : _GEN_2796; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3387 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_55 : _GEN_2797; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3388 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_56 : _GEN_2798; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3389 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_57 : _GEN_2799; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3390 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_58 : _GEN_2800; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3391 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_59 : _GEN_2801; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3392 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_60 : _GEN_2802; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3393 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_61 : _GEN_2803; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3394 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_62 : _GEN_2804; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3395 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_63 : _GEN_2805; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3396 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_64 : _GEN_2806; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3397 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_65 : _GEN_2807; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3398 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_66 : _GEN_2808; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3399 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_67 : _GEN_2809; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3400 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_68 : _GEN_2810; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3401 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_69 : _GEN_2811; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3402 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_70 : _GEN_2812; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3403 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_71 : _GEN_2813; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3404 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_72 : _GEN_2814; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3405 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_73 : _GEN_2815; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3406 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_74 : _GEN_2816; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3407 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_75 : _GEN_2817; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3408 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_76 : _GEN_2818; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3409 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_77 : _GEN_2819; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3410 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_78 : _GEN_2820; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3411 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_79 : _GEN_2821; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3412 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_80 : _GEN_2822; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3413 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_81 : _GEN_2823; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3414 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_82 : _GEN_2824; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3415 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_83 : _GEN_2825; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3416 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_84 : _GEN_2826; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3417 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_85 : _GEN_2827; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3418 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_86 : _GEN_2828; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3419 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_87 : _GEN_2829; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3420 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_88 : _GEN_2830; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3421 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_89 : _GEN_2831; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3422 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_90 : _GEN_2832; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3423 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_91 : _GEN_2833; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3424 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_92 : _GEN_2834; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3425 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_93 : _GEN_2835; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3426 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_94 : _GEN_2836; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3427 = 2'h1 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_95 : _GEN_2837; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire  _GEN_3428 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_is_valid_processor : _GEN_2838; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire  _GEN_3429 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_next_config_id : _GEN_2839; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [1:0] _GEN_3430 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_next_processor_id : _GEN_2840; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3431 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_parse_transition_field : _GEN_2841; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3432 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_parse_current_offset : _GEN_2842; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3433 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_parse_current_state : _GEN_2843; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3434 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_0 : _GEN_2844; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3435 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_1 : _GEN_2845; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3436 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_2 : _GEN_2846; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3437 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_3 : _GEN_2847; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3438 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_4 : _GEN_2848; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3439 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_5 : _GEN_2849; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3440 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_6 : _GEN_2850; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3441 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_7 : _GEN_2851; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3442 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_8 : _GEN_2852; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3443 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_9 : _GEN_2853; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3444 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_10 : _GEN_2854; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3445 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_11 : _GEN_2855; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3446 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_12 : _GEN_2856; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3447 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_13 : _GEN_2857; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3448 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_14 : _GEN_2858; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3449 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_15 : _GEN_2859; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3450 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_0 : _GEN_2860; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3451 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_1 : _GEN_2861; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3452 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_2 : _GEN_2862; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3453 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_3 : _GEN_2863; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3454 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_4 : _GEN_2864; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3455 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_5 : _GEN_2865; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3456 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_6 : _GEN_2866; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3457 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_7 : _GEN_2867; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3458 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_8 : _GEN_2868; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3459 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_9 : _GEN_2869; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3460 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_10 : _GEN_2870; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3461 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_11 : _GEN_2871; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3462 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_12 : _GEN_2872; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3463 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_13 : _GEN_2873; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3464 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_14 : _GEN_2874; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3465 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_15 : _GEN_2875; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3466 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_16 : _GEN_2876; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3467 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_17 : _GEN_2877; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3468 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_18 : _GEN_2878; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3469 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_19 : _GEN_2879; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3470 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_20 : _GEN_2880; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3471 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_21 : _GEN_2881; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3472 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_22 : _GEN_2882; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3473 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_23 : _GEN_2883; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3474 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_24 : _GEN_2884; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3475 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_25 : _GEN_2885; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3476 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_26 : _GEN_2886; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3477 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_27 : _GEN_2887; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3478 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_28 : _GEN_2888; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3479 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_29 : _GEN_2889; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3480 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_30 : _GEN_2890; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3481 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_31 : _GEN_2891; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3482 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_32 : _GEN_2892; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3483 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_33 : _GEN_2893; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3484 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_34 : _GEN_2894; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3485 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_35 : _GEN_2895; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3486 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_36 : _GEN_2896; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3487 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_37 : _GEN_2897; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3488 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_38 : _GEN_2898; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3489 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_39 : _GEN_2899; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3490 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_40 : _GEN_2900; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3491 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_41 : _GEN_2901; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3492 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_42 : _GEN_2902; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3493 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_43 : _GEN_2903; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3494 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_44 : _GEN_2904; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3495 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_45 : _GEN_2905; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3496 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_46 : _GEN_2906; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3497 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_47 : _GEN_2907; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3498 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_48 : _GEN_2908; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3499 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_49 : _GEN_2909; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3500 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_50 : _GEN_2910; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3501 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_51 : _GEN_2911; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3502 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_52 : _GEN_2912; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3503 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_53 : _GEN_2913; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3504 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_54 : _GEN_2914; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3505 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_55 : _GEN_2915; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3506 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_56 : _GEN_2916; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3507 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_57 : _GEN_2917; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3508 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_58 : _GEN_2918; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3509 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_59 : _GEN_2919; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3510 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_60 : _GEN_2920; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3511 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_61 : _GEN_2921; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3512 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_62 : _GEN_2922; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3513 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_63 : _GEN_2923; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3514 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_64 : _GEN_2924; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3515 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_65 : _GEN_2925; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3516 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_66 : _GEN_2926; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3517 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_67 : _GEN_2927; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3518 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_68 : _GEN_2928; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3519 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_69 : _GEN_2929; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3520 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_70 : _GEN_2930; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3521 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_71 : _GEN_2931; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3522 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_72 : _GEN_2932; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3523 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_73 : _GEN_2933; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3524 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_74 : _GEN_2934; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3525 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_75 : _GEN_2935; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3526 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_76 : _GEN_2936; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3527 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_77 : _GEN_2937; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3528 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_78 : _GEN_2938; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3529 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_79 : _GEN_2939; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3530 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_80 : _GEN_2940; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3531 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_81 : _GEN_2941; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3532 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_82 : _GEN_2942; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3533 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_83 : _GEN_2943; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3534 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_84 : _GEN_2944; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3535 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_85 : _GEN_2945; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3536 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_86 : _GEN_2946; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3537 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_87 : _GEN_2947; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3538 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_88 : _GEN_2948; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3539 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_89 : _GEN_2949; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3540 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_90 : _GEN_2950; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3541 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_91 : _GEN_2951; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3542 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_92 : _GEN_2952; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3543 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_93 : _GEN_2953; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3544 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_94 : _GEN_2954; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3545 = 2'h2 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_95 : _GEN_2955; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire  _GEN_3546 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_is_valid_processor : _GEN_2956; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire  _GEN_3547 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_next_config_id : _GEN_2957; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [1:0] _GEN_3548 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_next_processor_id : _GEN_2958; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3549 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_parse_transition_field : _GEN_2959; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3550 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_parse_current_offset : _GEN_2960; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3551 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_parse_current_state : _GEN_2961; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3552 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_0 : _GEN_2962; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3553 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_1 : _GEN_2963; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3554 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_2 : _GEN_2964; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3555 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_3 : _GEN_2965; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3556 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_4 : _GEN_2966; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3557 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_5 : _GEN_2967; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3558 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_6 : _GEN_2968; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3559 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_7 : _GEN_2969; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3560 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_8 : _GEN_2970; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3561 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_9 : _GEN_2971; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3562 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_10 : _GEN_2972; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3563 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_11 : _GEN_2973; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3564 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_12 : _GEN_2974; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3565 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_13 : _GEN_2975; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3566 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_14 : _GEN_2976; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [15:0] _GEN_3567 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_header_15 : _GEN_2977; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3568 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_0 : _GEN_2978; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3569 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_1 : _GEN_2979; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3570 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_2 : _GEN_2980; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3571 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_3 : _GEN_2981; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3572 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_4 : _GEN_2982; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3573 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_5 : _GEN_2983; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3574 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_6 : _GEN_2984; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3575 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_7 : _GEN_2985; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3576 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_8 : _GEN_2986; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3577 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_9 : _GEN_2987; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3578 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_10 : _GEN_2988; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3579 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_11 : _GEN_2989; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3580 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_12 : _GEN_2990; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3581 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_13 : _GEN_2991; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3582 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_14 : _GEN_2992; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3583 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_15 : _GEN_2993; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3584 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_16 : _GEN_2994; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3585 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_17 : _GEN_2995; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3586 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_18 : _GEN_2996; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3587 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_19 : _GEN_2997; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3588 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_20 : _GEN_2998; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3589 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_21 : _GEN_2999; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3590 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_22 : _GEN_3000; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3591 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_23 : _GEN_3001; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3592 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_24 : _GEN_3002; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3593 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_25 : _GEN_3003; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3594 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_26 : _GEN_3004; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3595 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_27 : _GEN_3005; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3596 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_28 : _GEN_3006; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3597 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_29 : _GEN_3007; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3598 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_30 : _GEN_3008; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3599 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_31 : _GEN_3009; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3600 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_32 : _GEN_3010; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3601 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_33 : _GEN_3011; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3602 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_34 : _GEN_3012; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3603 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_35 : _GEN_3013; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3604 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_36 : _GEN_3014; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3605 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_37 : _GEN_3015; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3606 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_38 : _GEN_3016; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3607 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_39 : _GEN_3017; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3608 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_40 : _GEN_3018; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3609 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_41 : _GEN_3019; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3610 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_42 : _GEN_3020; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3611 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_43 : _GEN_3021; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3612 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_44 : _GEN_3022; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3613 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_45 : _GEN_3023; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3614 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_46 : _GEN_3024; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3615 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_47 : _GEN_3025; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3616 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_48 : _GEN_3026; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3617 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_49 : _GEN_3027; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3618 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_50 : _GEN_3028; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3619 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_51 : _GEN_3029; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3620 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_52 : _GEN_3030; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3621 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_53 : _GEN_3031; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3622 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_54 : _GEN_3032; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3623 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_55 : _GEN_3033; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3624 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_56 : _GEN_3034; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3625 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_57 : _GEN_3035; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3626 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_58 : _GEN_3036; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3627 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_59 : _GEN_3037; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3628 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_60 : _GEN_3038; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3629 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_61 : _GEN_3039; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3630 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_62 : _GEN_3040; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3631 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_63 : _GEN_3041; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3632 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_64 : _GEN_3042; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3633 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_65 : _GEN_3043; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3634 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_66 : _GEN_3044; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3635 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_67 : _GEN_3045; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3636 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_68 : _GEN_3046; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3637 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_69 : _GEN_3047; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3638 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_70 : _GEN_3048; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3639 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_71 : _GEN_3049; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3640 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_72 : _GEN_3050; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3641 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_73 : _GEN_3051; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3642 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_74 : _GEN_3052; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3643 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_75 : _GEN_3053; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3644 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_76 : _GEN_3054; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3645 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_77 : _GEN_3055; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3646 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_78 : _GEN_3056; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3647 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_79 : _GEN_3057; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3648 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_80 : _GEN_3058; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3649 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_81 : _GEN_3059; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3650 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_82 : _GEN_3060; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3651 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_83 : _GEN_3061; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3652 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_84 : _GEN_3062; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3653 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_85 : _GEN_3063; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3654 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_86 : _GEN_3064; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3655 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_87 : _GEN_3065; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3656 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_88 : _GEN_3066; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3657 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_89 : _GEN_3067; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3658 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_90 : _GEN_3068; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3659 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_91 : _GEN_3069; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3660 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_92 : _GEN_3070; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3661 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_93 : _GEN_3071; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3662 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_94 : _GEN_3072; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  wire [7:0] _GEN_3663 = 2'h3 == next_proc_id_3 ? trans_3_io_pipe_phv_out_data_95 : _GEN_3073; // @[ipsa.scala 96:76 ipsa.scala 97:44]
  Processor proc_0 ( // @[ipsa.scala 56:25]
    .clock(proc_0_clock),
    .io_pipe_phv_in_data_0(proc_0_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_0_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_0_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_0_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_0_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_0_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_0_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_0_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_0_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_0_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_0_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_0_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_0_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_0_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_0_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_0_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_0_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_0_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_0_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_0_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_0_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_0_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_0_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_0_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_0_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_0_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_0_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_0_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_0_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_0_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_0_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_0_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_0_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_0_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_0_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_0_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_0_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_0_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_0_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_0_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_0_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_0_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_0_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_0_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_0_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_0_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_0_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_0_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_0_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_0_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_0_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_0_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_0_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_0_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_0_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_0_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_0_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_0_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_0_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_0_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_0_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_0_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_0_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_0_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_0_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_0_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_0_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_0_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_0_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_0_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_0_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_0_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_0_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_0_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_0_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_0_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_0_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_0_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_0_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_0_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_0_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_0_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_0_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_0_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_0_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_0_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_0_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_0_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_0_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_0_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_0_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_0_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_0_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_0_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_0_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_0_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(proc_0_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(proc_0_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(proc_0_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(proc_0_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(proc_0_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(proc_0_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(proc_0_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(proc_0_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(proc_0_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(proc_0_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(proc_0_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(proc_0_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(proc_0_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(proc_0_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(proc_0_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(proc_0_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(proc_0_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(proc_0_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(proc_0_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(proc_0_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_0_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_0_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(proc_0_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_0_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_0_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_0_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_0_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_0_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_0_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_0_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_0_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_0_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_0_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_0_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_0_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_0_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_0_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_0_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_0_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_0_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_0_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_0_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_0_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_0_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_0_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_0_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_0_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_0_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_0_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_0_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_0_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_0_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_0_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_0_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_0_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_0_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_0_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_0_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_0_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_0_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_0_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_0_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_0_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_0_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_0_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_0_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_0_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_0_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_0_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_0_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_0_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_0_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_0_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_0_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_0_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_0_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_0_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_0_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_0_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_0_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_0_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_0_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_0_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_0_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_0_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_0_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_0_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_0_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_0_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_0_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_0_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_0_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_0_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_0_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_0_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_0_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_0_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_0_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_0_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_0_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_0_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_0_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_0_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_0_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_0_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_0_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_0_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_0_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_0_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_0_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_0_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_0_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_0_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_0_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_0_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_0_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_0_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_0_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(proc_0_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(proc_0_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(proc_0_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(proc_0_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(proc_0_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(proc_0_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(proc_0_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(proc_0_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(proc_0_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(proc_0_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(proc_0_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(proc_0_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(proc_0_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(proc_0_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(proc_0_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(proc_0_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(proc_0_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(proc_0_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(proc_0_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(proc_0_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_0_io_pipe_phv_out_next_config_id),
    .io_mod_par_mod_en(proc_0_io_mod_par_mod_en),
    .io_mod_par_mod_last_mau_id_mod(proc_0_io_mod_par_mod_last_mau_id_mod),
    .io_mod_par_mod_last_mau_id(proc_0_io_mod_par_mod_last_mau_id),
    .io_mod_par_mod_cs(proc_0_io_mod_par_mod_cs),
    .io_mod_par_mod_module_mod_state_id_mod(proc_0_io_mod_par_mod_module_mod_state_id_mod),
    .io_mod_par_mod_module_mod_state_id(proc_0_io_mod_par_mod_module_mod_state_id),
    .io_mod_par_mod_module_mod_sram_w_cs(proc_0_io_mod_par_mod_module_mod_sram_w_cs),
    .io_mod_par_mod_module_mod_sram_w_addr(proc_0_io_mod_par_mod_module_mod_sram_w_addr),
    .io_mod_par_mod_module_mod_sram_w_data(proc_0_io_mod_par_mod_module_mod_sram_w_data),
    .io_mod_mat_mod_en(proc_0_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_0_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_header_id(proc_0_io_mod_mat_mod_key_mod_header_id),
    .io_mod_mat_mod_key_mod_internal_offset(proc_0_io_mod_mat_mod_key_mod_internal_offset),
    .io_mod_mat_mod_key_mod_key_length(proc_0_io_mod_mat_mod_key_mod_key_length),
    .io_mod_mat_mod_table_mod_table_width(proc_0_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_table_mod_table_depth(proc_0_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_act_mod_en(proc_0_io_mod_act_mod_en),
    .io_mod_act_mod_addr(proc_0_io_mod_act_mod_addr),
    .io_mod_act_mod_data_0(proc_0_io_mod_act_mod_data_0),
    .io_mod_act_mod_data_1(proc_0_io_mod_act_mod_data_1),
    .io_mem_cluster_0_en(proc_0_io_mem_cluster_0_en),
    .io_mem_cluster_0_addr(proc_0_io_mem_cluster_0_addr),
    .io_mem_cluster_0_data(proc_0_io_mem_cluster_0_data),
    .io_mem_cluster_1_en(proc_0_io_mem_cluster_1_en),
    .io_mem_cluster_1_addr(proc_0_io_mem_cluster_1_addr),
    .io_mem_cluster_1_data(proc_0_io_mem_cluster_1_data),
    .io_mem_cluster_2_en(proc_0_io_mem_cluster_2_en),
    .io_mem_cluster_2_addr(proc_0_io_mem_cluster_2_addr),
    .io_mem_cluster_2_data(proc_0_io_mem_cluster_2_data),
    .io_mem_cluster_3_en(proc_0_io_mem_cluster_3_en),
    .io_mem_cluster_3_addr(proc_0_io_mem_cluster_3_addr),
    .io_mem_cluster_3_data(proc_0_io_mem_cluster_3_data),
    .io_mem_cluster_4_en(proc_0_io_mem_cluster_4_en),
    .io_mem_cluster_4_addr(proc_0_io_mem_cluster_4_addr),
    .io_mem_cluster_4_data(proc_0_io_mem_cluster_4_data),
    .io_mem_cluster_5_en(proc_0_io_mem_cluster_5_en),
    .io_mem_cluster_5_addr(proc_0_io_mem_cluster_5_addr),
    .io_mem_cluster_5_data(proc_0_io_mem_cluster_5_data),
    .io_mem_cluster_6_en(proc_0_io_mem_cluster_6_en),
    .io_mem_cluster_6_addr(proc_0_io_mem_cluster_6_addr),
    .io_mem_cluster_6_data(proc_0_io_mem_cluster_6_data),
    .io_mem_cluster_7_en(proc_0_io_mem_cluster_7_en),
    .io_mem_cluster_7_addr(proc_0_io_mem_cluster_7_addr),
    .io_mem_cluster_7_data(proc_0_io_mem_cluster_7_data)
  );
  Processor proc_1 ( // @[ipsa.scala 56:25]
    .clock(proc_1_clock),
    .io_pipe_phv_in_data_0(proc_1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(proc_1_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(proc_1_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(proc_1_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(proc_1_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(proc_1_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(proc_1_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(proc_1_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(proc_1_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(proc_1_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(proc_1_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(proc_1_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(proc_1_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(proc_1_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(proc_1_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(proc_1_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(proc_1_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(proc_1_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(proc_1_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(proc_1_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(proc_1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_1_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(proc_1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(proc_1_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(proc_1_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(proc_1_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(proc_1_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(proc_1_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(proc_1_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(proc_1_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(proc_1_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(proc_1_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(proc_1_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(proc_1_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(proc_1_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(proc_1_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(proc_1_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(proc_1_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(proc_1_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(proc_1_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(proc_1_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(proc_1_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(proc_1_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_1_io_pipe_phv_out_next_config_id),
    .io_mod_par_mod_en(proc_1_io_mod_par_mod_en),
    .io_mod_par_mod_last_mau_id_mod(proc_1_io_mod_par_mod_last_mau_id_mod),
    .io_mod_par_mod_last_mau_id(proc_1_io_mod_par_mod_last_mau_id),
    .io_mod_par_mod_cs(proc_1_io_mod_par_mod_cs),
    .io_mod_par_mod_module_mod_state_id_mod(proc_1_io_mod_par_mod_module_mod_state_id_mod),
    .io_mod_par_mod_module_mod_state_id(proc_1_io_mod_par_mod_module_mod_state_id),
    .io_mod_par_mod_module_mod_sram_w_cs(proc_1_io_mod_par_mod_module_mod_sram_w_cs),
    .io_mod_par_mod_module_mod_sram_w_addr(proc_1_io_mod_par_mod_module_mod_sram_w_addr),
    .io_mod_par_mod_module_mod_sram_w_data(proc_1_io_mod_par_mod_module_mod_sram_w_data),
    .io_mod_mat_mod_en(proc_1_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_1_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_header_id(proc_1_io_mod_mat_mod_key_mod_header_id),
    .io_mod_mat_mod_key_mod_internal_offset(proc_1_io_mod_mat_mod_key_mod_internal_offset),
    .io_mod_mat_mod_key_mod_key_length(proc_1_io_mod_mat_mod_key_mod_key_length),
    .io_mod_mat_mod_table_mod_table_width(proc_1_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_table_mod_table_depth(proc_1_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_act_mod_en(proc_1_io_mod_act_mod_en),
    .io_mod_act_mod_addr(proc_1_io_mod_act_mod_addr),
    .io_mod_act_mod_data_0(proc_1_io_mod_act_mod_data_0),
    .io_mod_act_mod_data_1(proc_1_io_mod_act_mod_data_1),
    .io_mem_cluster_0_en(proc_1_io_mem_cluster_0_en),
    .io_mem_cluster_0_addr(proc_1_io_mem_cluster_0_addr),
    .io_mem_cluster_0_data(proc_1_io_mem_cluster_0_data),
    .io_mem_cluster_1_en(proc_1_io_mem_cluster_1_en),
    .io_mem_cluster_1_addr(proc_1_io_mem_cluster_1_addr),
    .io_mem_cluster_1_data(proc_1_io_mem_cluster_1_data),
    .io_mem_cluster_2_en(proc_1_io_mem_cluster_2_en),
    .io_mem_cluster_2_addr(proc_1_io_mem_cluster_2_addr),
    .io_mem_cluster_2_data(proc_1_io_mem_cluster_2_data),
    .io_mem_cluster_3_en(proc_1_io_mem_cluster_3_en),
    .io_mem_cluster_3_addr(proc_1_io_mem_cluster_3_addr),
    .io_mem_cluster_3_data(proc_1_io_mem_cluster_3_data),
    .io_mem_cluster_4_en(proc_1_io_mem_cluster_4_en),
    .io_mem_cluster_4_addr(proc_1_io_mem_cluster_4_addr),
    .io_mem_cluster_4_data(proc_1_io_mem_cluster_4_data),
    .io_mem_cluster_5_en(proc_1_io_mem_cluster_5_en),
    .io_mem_cluster_5_addr(proc_1_io_mem_cluster_5_addr),
    .io_mem_cluster_5_data(proc_1_io_mem_cluster_5_data),
    .io_mem_cluster_6_en(proc_1_io_mem_cluster_6_en),
    .io_mem_cluster_6_addr(proc_1_io_mem_cluster_6_addr),
    .io_mem_cluster_6_data(proc_1_io_mem_cluster_6_data),
    .io_mem_cluster_7_en(proc_1_io_mem_cluster_7_en),
    .io_mem_cluster_7_addr(proc_1_io_mem_cluster_7_addr),
    .io_mem_cluster_7_data(proc_1_io_mem_cluster_7_data)
  );
  Processor proc_2 ( // @[ipsa.scala 56:25]
    .clock(proc_2_clock),
    .io_pipe_phv_in_data_0(proc_2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(proc_2_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(proc_2_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(proc_2_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(proc_2_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(proc_2_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(proc_2_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(proc_2_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(proc_2_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(proc_2_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(proc_2_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(proc_2_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(proc_2_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(proc_2_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(proc_2_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(proc_2_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(proc_2_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(proc_2_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(proc_2_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(proc_2_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(proc_2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_2_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(proc_2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(proc_2_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(proc_2_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(proc_2_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(proc_2_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(proc_2_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(proc_2_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(proc_2_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(proc_2_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(proc_2_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(proc_2_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(proc_2_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(proc_2_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(proc_2_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(proc_2_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(proc_2_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(proc_2_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(proc_2_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(proc_2_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(proc_2_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(proc_2_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_2_io_pipe_phv_out_next_config_id),
    .io_mod_par_mod_en(proc_2_io_mod_par_mod_en),
    .io_mod_par_mod_last_mau_id_mod(proc_2_io_mod_par_mod_last_mau_id_mod),
    .io_mod_par_mod_last_mau_id(proc_2_io_mod_par_mod_last_mau_id),
    .io_mod_par_mod_cs(proc_2_io_mod_par_mod_cs),
    .io_mod_par_mod_module_mod_state_id_mod(proc_2_io_mod_par_mod_module_mod_state_id_mod),
    .io_mod_par_mod_module_mod_state_id(proc_2_io_mod_par_mod_module_mod_state_id),
    .io_mod_par_mod_module_mod_sram_w_cs(proc_2_io_mod_par_mod_module_mod_sram_w_cs),
    .io_mod_par_mod_module_mod_sram_w_addr(proc_2_io_mod_par_mod_module_mod_sram_w_addr),
    .io_mod_par_mod_module_mod_sram_w_data(proc_2_io_mod_par_mod_module_mod_sram_w_data),
    .io_mod_mat_mod_en(proc_2_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_2_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_header_id(proc_2_io_mod_mat_mod_key_mod_header_id),
    .io_mod_mat_mod_key_mod_internal_offset(proc_2_io_mod_mat_mod_key_mod_internal_offset),
    .io_mod_mat_mod_key_mod_key_length(proc_2_io_mod_mat_mod_key_mod_key_length),
    .io_mod_mat_mod_table_mod_table_width(proc_2_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_table_mod_table_depth(proc_2_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_act_mod_en(proc_2_io_mod_act_mod_en),
    .io_mod_act_mod_addr(proc_2_io_mod_act_mod_addr),
    .io_mod_act_mod_data_0(proc_2_io_mod_act_mod_data_0),
    .io_mod_act_mod_data_1(proc_2_io_mod_act_mod_data_1),
    .io_mem_cluster_0_en(proc_2_io_mem_cluster_0_en),
    .io_mem_cluster_0_addr(proc_2_io_mem_cluster_0_addr),
    .io_mem_cluster_0_data(proc_2_io_mem_cluster_0_data),
    .io_mem_cluster_1_en(proc_2_io_mem_cluster_1_en),
    .io_mem_cluster_1_addr(proc_2_io_mem_cluster_1_addr),
    .io_mem_cluster_1_data(proc_2_io_mem_cluster_1_data),
    .io_mem_cluster_2_en(proc_2_io_mem_cluster_2_en),
    .io_mem_cluster_2_addr(proc_2_io_mem_cluster_2_addr),
    .io_mem_cluster_2_data(proc_2_io_mem_cluster_2_data),
    .io_mem_cluster_3_en(proc_2_io_mem_cluster_3_en),
    .io_mem_cluster_3_addr(proc_2_io_mem_cluster_3_addr),
    .io_mem_cluster_3_data(proc_2_io_mem_cluster_3_data),
    .io_mem_cluster_4_en(proc_2_io_mem_cluster_4_en),
    .io_mem_cluster_4_addr(proc_2_io_mem_cluster_4_addr),
    .io_mem_cluster_4_data(proc_2_io_mem_cluster_4_data),
    .io_mem_cluster_5_en(proc_2_io_mem_cluster_5_en),
    .io_mem_cluster_5_addr(proc_2_io_mem_cluster_5_addr),
    .io_mem_cluster_5_data(proc_2_io_mem_cluster_5_data),
    .io_mem_cluster_6_en(proc_2_io_mem_cluster_6_en),
    .io_mem_cluster_6_addr(proc_2_io_mem_cluster_6_addr),
    .io_mem_cluster_6_data(proc_2_io_mem_cluster_6_data),
    .io_mem_cluster_7_en(proc_2_io_mem_cluster_7_en),
    .io_mem_cluster_7_addr(proc_2_io_mem_cluster_7_addr),
    .io_mem_cluster_7_data(proc_2_io_mem_cluster_7_data)
  );
  Processor proc_3 ( // @[ipsa.scala 56:25]
    .clock(proc_3_clock),
    .io_pipe_phv_in_data_0(proc_3_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_3_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_3_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_3_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_3_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_3_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_3_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_3_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_3_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_3_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_3_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_3_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_3_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_3_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_3_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_3_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_3_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_3_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_3_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_3_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_3_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_3_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_3_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_3_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_3_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_3_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_3_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_3_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_3_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_3_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_3_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_3_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_3_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_3_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_3_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_3_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_3_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_3_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_3_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_3_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_3_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_3_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_3_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_3_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_3_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_3_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_3_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_3_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_3_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_3_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_3_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_3_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_3_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_3_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_3_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_3_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_3_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_3_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_3_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_3_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_3_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_3_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_3_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_3_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_3_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_3_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_3_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_3_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_3_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_3_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_3_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_3_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_3_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_3_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_3_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_3_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_3_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_3_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_3_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_3_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_3_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_3_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_3_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_3_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_3_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_3_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_3_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_3_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_3_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_3_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_3_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_3_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_3_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_3_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_3_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_3_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(proc_3_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(proc_3_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(proc_3_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(proc_3_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(proc_3_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(proc_3_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(proc_3_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(proc_3_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(proc_3_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(proc_3_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(proc_3_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(proc_3_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(proc_3_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(proc_3_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(proc_3_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(proc_3_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(proc_3_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(proc_3_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(proc_3_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(proc_3_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_3_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_3_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(proc_3_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_3_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_3_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_3_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_3_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_3_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_3_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_3_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_3_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_3_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_3_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_3_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_3_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_3_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_3_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_3_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_3_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_3_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_3_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_3_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_3_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_3_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_3_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_3_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_3_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_3_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_3_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_3_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_3_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_3_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_3_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_3_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_3_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_3_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_3_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_3_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_3_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_3_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_3_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_3_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_3_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_3_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_3_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_3_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_3_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_3_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_3_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_3_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_3_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_3_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_3_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_3_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_3_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_3_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_3_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_3_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_3_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_3_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_3_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_3_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_3_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_3_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_3_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_3_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_3_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_3_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_3_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_3_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_3_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_3_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_3_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_3_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_3_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_3_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_3_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_3_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_3_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_3_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_3_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_3_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_3_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_3_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_3_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_3_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_3_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_3_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_3_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_3_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_3_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_3_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_3_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_3_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_3_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_3_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_3_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_3_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(proc_3_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(proc_3_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(proc_3_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(proc_3_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(proc_3_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(proc_3_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(proc_3_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(proc_3_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(proc_3_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(proc_3_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(proc_3_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(proc_3_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(proc_3_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(proc_3_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(proc_3_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(proc_3_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(proc_3_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(proc_3_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(proc_3_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(proc_3_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_3_io_pipe_phv_out_next_config_id),
    .io_mod_par_mod_en(proc_3_io_mod_par_mod_en),
    .io_mod_par_mod_last_mau_id_mod(proc_3_io_mod_par_mod_last_mau_id_mod),
    .io_mod_par_mod_last_mau_id(proc_3_io_mod_par_mod_last_mau_id),
    .io_mod_par_mod_cs(proc_3_io_mod_par_mod_cs),
    .io_mod_par_mod_module_mod_state_id_mod(proc_3_io_mod_par_mod_module_mod_state_id_mod),
    .io_mod_par_mod_module_mod_state_id(proc_3_io_mod_par_mod_module_mod_state_id),
    .io_mod_par_mod_module_mod_sram_w_cs(proc_3_io_mod_par_mod_module_mod_sram_w_cs),
    .io_mod_par_mod_module_mod_sram_w_addr(proc_3_io_mod_par_mod_module_mod_sram_w_addr),
    .io_mod_par_mod_module_mod_sram_w_data(proc_3_io_mod_par_mod_module_mod_sram_w_data),
    .io_mod_mat_mod_en(proc_3_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_3_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_header_id(proc_3_io_mod_mat_mod_key_mod_header_id),
    .io_mod_mat_mod_key_mod_internal_offset(proc_3_io_mod_mat_mod_key_mod_internal_offset),
    .io_mod_mat_mod_key_mod_key_length(proc_3_io_mod_mat_mod_key_mod_key_length),
    .io_mod_mat_mod_table_mod_table_width(proc_3_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_table_mod_table_depth(proc_3_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_act_mod_en(proc_3_io_mod_act_mod_en),
    .io_mod_act_mod_addr(proc_3_io_mod_act_mod_addr),
    .io_mod_act_mod_data_0(proc_3_io_mod_act_mod_data_0),
    .io_mod_act_mod_data_1(proc_3_io_mod_act_mod_data_1),
    .io_mem_cluster_0_en(proc_3_io_mem_cluster_0_en),
    .io_mem_cluster_0_addr(proc_3_io_mem_cluster_0_addr),
    .io_mem_cluster_0_data(proc_3_io_mem_cluster_0_data),
    .io_mem_cluster_1_en(proc_3_io_mem_cluster_1_en),
    .io_mem_cluster_1_addr(proc_3_io_mem_cluster_1_addr),
    .io_mem_cluster_1_data(proc_3_io_mem_cluster_1_data),
    .io_mem_cluster_2_en(proc_3_io_mem_cluster_2_en),
    .io_mem_cluster_2_addr(proc_3_io_mem_cluster_2_addr),
    .io_mem_cluster_2_data(proc_3_io_mem_cluster_2_data),
    .io_mem_cluster_3_en(proc_3_io_mem_cluster_3_en),
    .io_mem_cluster_3_addr(proc_3_io_mem_cluster_3_addr),
    .io_mem_cluster_3_data(proc_3_io_mem_cluster_3_data),
    .io_mem_cluster_4_en(proc_3_io_mem_cluster_4_en),
    .io_mem_cluster_4_addr(proc_3_io_mem_cluster_4_addr),
    .io_mem_cluster_4_data(proc_3_io_mem_cluster_4_data),
    .io_mem_cluster_5_en(proc_3_io_mem_cluster_5_en),
    .io_mem_cluster_5_addr(proc_3_io_mem_cluster_5_addr),
    .io_mem_cluster_5_data(proc_3_io_mem_cluster_5_data),
    .io_mem_cluster_6_en(proc_3_io_mem_cluster_6_en),
    .io_mem_cluster_6_addr(proc_3_io_mem_cluster_6_addr),
    .io_mem_cluster_6_data(proc_3_io_mem_cluster_6_data),
    .io_mem_cluster_7_en(proc_3_io_mem_cluster_7_en),
    .io_mem_cluster_7_addr(proc_3_io_mem_cluster_7_addr),
    .io_mem_cluster_7_data(proc_3_io_mem_cluster_7_data)
  );
  SRAMCluster sram_cluster_0 ( // @[ipsa.scala 62:25]
    .clock(sram_cluster_0_clock),
    .io_w_wcs(sram_cluster_0_io_w_wcs),
    .io_w_w_en(sram_cluster_0_io_w_w_en),
    .io_w_w_addr(sram_cluster_0_io_w_w_addr),
    .io_w_w_data(sram_cluster_0_io_w_w_data),
    .io_r_0_cluster_0_en(sram_cluster_0_io_r_0_cluster_0_en),
    .io_r_0_cluster_0_addr(sram_cluster_0_io_r_0_cluster_0_addr),
    .io_r_0_cluster_0_data(sram_cluster_0_io_r_0_cluster_0_data),
    .io_r_0_cluster_1_en(sram_cluster_0_io_r_0_cluster_1_en),
    .io_r_0_cluster_1_addr(sram_cluster_0_io_r_0_cluster_1_addr),
    .io_r_0_cluster_1_data(sram_cluster_0_io_r_0_cluster_1_data),
    .io_r_0_cluster_2_en(sram_cluster_0_io_r_0_cluster_2_en),
    .io_r_0_cluster_2_addr(sram_cluster_0_io_r_0_cluster_2_addr),
    .io_r_0_cluster_2_data(sram_cluster_0_io_r_0_cluster_2_data),
    .io_r_0_cluster_3_en(sram_cluster_0_io_r_0_cluster_3_en),
    .io_r_0_cluster_3_addr(sram_cluster_0_io_r_0_cluster_3_addr),
    .io_r_0_cluster_3_data(sram_cluster_0_io_r_0_cluster_3_data),
    .io_r_0_cluster_4_en(sram_cluster_0_io_r_0_cluster_4_en),
    .io_r_0_cluster_4_addr(sram_cluster_0_io_r_0_cluster_4_addr),
    .io_r_0_cluster_4_data(sram_cluster_0_io_r_0_cluster_4_data),
    .io_r_0_cluster_5_en(sram_cluster_0_io_r_0_cluster_5_en),
    .io_r_0_cluster_5_addr(sram_cluster_0_io_r_0_cluster_5_addr),
    .io_r_0_cluster_5_data(sram_cluster_0_io_r_0_cluster_5_data),
    .io_r_0_cluster_6_en(sram_cluster_0_io_r_0_cluster_6_en),
    .io_r_0_cluster_6_addr(sram_cluster_0_io_r_0_cluster_6_addr),
    .io_r_0_cluster_6_data(sram_cluster_0_io_r_0_cluster_6_data),
    .io_r_0_cluster_7_en(sram_cluster_0_io_r_0_cluster_7_en),
    .io_r_0_cluster_7_addr(sram_cluster_0_io_r_0_cluster_7_addr),
    .io_r_0_cluster_7_data(sram_cluster_0_io_r_0_cluster_7_data),
    .io_r_1_cluster_0_en(sram_cluster_0_io_r_1_cluster_0_en),
    .io_r_1_cluster_0_addr(sram_cluster_0_io_r_1_cluster_0_addr),
    .io_r_1_cluster_0_data(sram_cluster_0_io_r_1_cluster_0_data),
    .io_r_1_cluster_1_en(sram_cluster_0_io_r_1_cluster_1_en),
    .io_r_1_cluster_1_addr(sram_cluster_0_io_r_1_cluster_1_addr),
    .io_r_1_cluster_1_data(sram_cluster_0_io_r_1_cluster_1_data),
    .io_r_1_cluster_2_en(sram_cluster_0_io_r_1_cluster_2_en),
    .io_r_1_cluster_2_addr(sram_cluster_0_io_r_1_cluster_2_addr),
    .io_r_1_cluster_2_data(sram_cluster_0_io_r_1_cluster_2_data),
    .io_r_1_cluster_3_en(sram_cluster_0_io_r_1_cluster_3_en),
    .io_r_1_cluster_3_addr(sram_cluster_0_io_r_1_cluster_3_addr),
    .io_r_1_cluster_3_data(sram_cluster_0_io_r_1_cluster_3_data),
    .io_r_1_cluster_4_en(sram_cluster_0_io_r_1_cluster_4_en),
    .io_r_1_cluster_4_addr(sram_cluster_0_io_r_1_cluster_4_addr),
    .io_r_1_cluster_4_data(sram_cluster_0_io_r_1_cluster_4_data),
    .io_r_1_cluster_5_en(sram_cluster_0_io_r_1_cluster_5_en),
    .io_r_1_cluster_5_addr(sram_cluster_0_io_r_1_cluster_5_addr),
    .io_r_1_cluster_5_data(sram_cluster_0_io_r_1_cluster_5_data),
    .io_r_1_cluster_6_en(sram_cluster_0_io_r_1_cluster_6_en),
    .io_r_1_cluster_6_addr(sram_cluster_0_io_r_1_cluster_6_addr),
    .io_r_1_cluster_6_data(sram_cluster_0_io_r_1_cluster_6_data),
    .io_r_1_cluster_7_en(sram_cluster_0_io_r_1_cluster_7_en),
    .io_r_1_cluster_7_addr(sram_cluster_0_io_r_1_cluster_7_addr),
    .io_r_1_cluster_7_data(sram_cluster_0_io_r_1_cluster_7_data),
    .io_r_2_cluster_0_en(sram_cluster_0_io_r_2_cluster_0_en),
    .io_r_2_cluster_0_addr(sram_cluster_0_io_r_2_cluster_0_addr),
    .io_r_2_cluster_0_data(sram_cluster_0_io_r_2_cluster_0_data),
    .io_r_2_cluster_1_en(sram_cluster_0_io_r_2_cluster_1_en),
    .io_r_2_cluster_1_addr(sram_cluster_0_io_r_2_cluster_1_addr),
    .io_r_2_cluster_1_data(sram_cluster_0_io_r_2_cluster_1_data),
    .io_r_2_cluster_2_en(sram_cluster_0_io_r_2_cluster_2_en),
    .io_r_2_cluster_2_addr(sram_cluster_0_io_r_2_cluster_2_addr),
    .io_r_2_cluster_2_data(sram_cluster_0_io_r_2_cluster_2_data),
    .io_r_2_cluster_3_en(sram_cluster_0_io_r_2_cluster_3_en),
    .io_r_2_cluster_3_addr(sram_cluster_0_io_r_2_cluster_3_addr),
    .io_r_2_cluster_3_data(sram_cluster_0_io_r_2_cluster_3_data),
    .io_r_2_cluster_4_en(sram_cluster_0_io_r_2_cluster_4_en),
    .io_r_2_cluster_4_addr(sram_cluster_0_io_r_2_cluster_4_addr),
    .io_r_2_cluster_4_data(sram_cluster_0_io_r_2_cluster_4_data),
    .io_r_2_cluster_5_en(sram_cluster_0_io_r_2_cluster_5_en),
    .io_r_2_cluster_5_addr(sram_cluster_0_io_r_2_cluster_5_addr),
    .io_r_2_cluster_5_data(sram_cluster_0_io_r_2_cluster_5_data),
    .io_r_2_cluster_6_en(sram_cluster_0_io_r_2_cluster_6_en),
    .io_r_2_cluster_6_addr(sram_cluster_0_io_r_2_cluster_6_addr),
    .io_r_2_cluster_6_data(sram_cluster_0_io_r_2_cluster_6_data),
    .io_r_2_cluster_7_en(sram_cluster_0_io_r_2_cluster_7_en),
    .io_r_2_cluster_7_addr(sram_cluster_0_io_r_2_cluster_7_addr),
    .io_r_2_cluster_7_data(sram_cluster_0_io_r_2_cluster_7_data),
    .io_r_3_cluster_0_en(sram_cluster_0_io_r_3_cluster_0_en),
    .io_r_3_cluster_0_addr(sram_cluster_0_io_r_3_cluster_0_addr),
    .io_r_3_cluster_0_data(sram_cluster_0_io_r_3_cluster_0_data),
    .io_r_3_cluster_1_en(sram_cluster_0_io_r_3_cluster_1_en),
    .io_r_3_cluster_1_addr(sram_cluster_0_io_r_3_cluster_1_addr),
    .io_r_3_cluster_1_data(sram_cluster_0_io_r_3_cluster_1_data),
    .io_r_3_cluster_2_en(sram_cluster_0_io_r_3_cluster_2_en),
    .io_r_3_cluster_2_addr(sram_cluster_0_io_r_3_cluster_2_addr),
    .io_r_3_cluster_2_data(sram_cluster_0_io_r_3_cluster_2_data),
    .io_r_3_cluster_3_en(sram_cluster_0_io_r_3_cluster_3_en),
    .io_r_3_cluster_3_addr(sram_cluster_0_io_r_3_cluster_3_addr),
    .io_r_3_cluster_3_data(sram_cluster_0_io_r_3_cluster_3_data),
    .io_r_3_cluster_4_en(sram_cluster_0_io_r_3_cluster_4_en),
    .io_r_3_cluster_4_addr(sram_cluster_0_io_r_3_cluster_4_addr),
    .io_r_3_cluster_4_data(sram_cluster_0_io_r_3_cluster_4_data),
    .io_r_3_cluster_5_en(sram_cluster_0_io_r_3_cluster_5_en),
    .io_r_3_cluster_5_addr(sram_cluster_0_io_r_3_cluster_5_addr),
    .io_r_3_cluster_5_data(sram_cluster_0_io_r_3_cluster_5_data),
    .io_r_3_cluster_6_en(sram_cluster_0_io_r_3_cluster_6_en),
    .io_r_3_cluster_6_addr(sram_cluster_0_io_r_3_cluster_6_addr),
    .io_r_3_cluster_6_data(sram_cluster_0_io_r_3_cluster_6_data),
    .io_r_3_cluster_7_en(sram_cluster_0_io_r_3_cluster_7_en),
    .io_r_3_cluster_7_addr(sram_cluster_0_io_r_3_cluster_7_addr),
    .io_r_3_cluster_7_data(sram_cluster_0_io_r_3_cluster_7_data)
  );
  Initializer init ( // @[ipsa.scala 74:22]
    .clock(init_clock),
    .io_pipe_phv_in_data_0(init_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(init_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(init_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(init_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(init_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(init_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(init_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(init_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(init_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(init_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(init_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(init_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(init_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(init_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(init_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(init_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(init_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(init_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(init_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(init_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(init_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(init_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(init_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(init_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(init_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(init_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(init_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(init_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(init_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(init_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(init_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(init_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(init_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(init_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(init_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(init_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(init_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(init_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(init_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(init_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(init_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(init_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(init_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(init_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(init_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(init_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(init_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(init_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(init_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(init_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(init_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(init_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(init_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(init_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(init_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(init_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(init_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(init_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(init_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(init_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(init_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(init_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(init_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(init_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(init_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(init_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(init_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(init_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(init_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(init_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(init_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(init_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(init_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(init_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(init_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(init_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(init_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(init_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(init_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(init_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(init_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(init_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(init_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(init_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(init_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(init_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(init_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(init_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(init_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(init_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(init_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(init_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(init_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(init_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(init_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(init_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(init_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(init_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(init_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(init_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(init_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(init_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(init_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(init_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(init_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(init_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(init_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(init_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(init_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(init_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(init_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(init_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(init_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(init_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(init_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_out_data_0(init_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(init_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(init_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(init_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(init_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(init_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(init_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(init_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(init_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(init_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(init_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(init_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(init_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(init_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(init_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(init_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(init_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(init_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(init_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(init_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(init_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(init_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(init_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(init_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(init_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(init_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(init_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(init_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(init_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(init_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(init_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(init_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(init_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(init_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(init_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(init_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(init_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(init_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(init_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(init_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(init_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(init_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(init_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(init_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(init_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(init_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(init_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(init_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(init_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(init_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(init_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(init_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(init_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(init_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(init_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(init_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(init_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(init_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(init_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(init_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(init_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(init_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(init_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(init_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(init_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(init_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(init_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(init_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(init_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(init_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(init_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(init_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(init_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(init_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(init_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(init_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(init_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(init_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(init_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(init_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(init_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(init_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(init_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(init_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(init_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(init_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(init_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(init_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(init_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(init_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(init_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(init_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(init_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(init_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(init_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(init_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(init_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(init_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(init_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(init_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(init_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(init_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(init_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(init_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(init_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(init_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(init_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(init_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(init_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(init_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(init_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(init_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(init_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(init_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(init_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(init_io_pipe_phv_out_next_processor_id),
    .io_first_proc_id(init_io_first_proc_id)
  );
  InterProcessorTransfer trans_0 ( // @[ipsa.scala 79:25]
    .clock(trans_0_clock),
    .io_pipe_phv_in_data_0(trans_0_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(trans_0_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(trans_0_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(trans_0_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(trans_0_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(trans_0_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(trans_0_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(trans_0_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(trans_0_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(trans_0_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(trans_0_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(trans_0_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(trans_0_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(trans_0_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(trans_0_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(trans_0_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(trans_0_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(trans_0_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(trans_0_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(trans_0_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(trans_0_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(trans_0_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(trans_0_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(trans_0_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(trans_0_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(trans_0_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(trans_0_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(trans_0_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(trans_0_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(trans_0_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(trans_0_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(trans_0_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(trans_0_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(trans_0_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(trans_0_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(trans_0_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(trans_0_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(trans_0_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(trans_0_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(trans_0_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(trans_0_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(trans_0_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(trans_0_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(trans_0_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(trans_0_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(trans_0_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(trans_0_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(trans_0_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(trans_0_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(trans_0_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(trans_0_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(trans_0_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(trans_0_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(trans_0_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(trans_0_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(trans_0_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(trans_0_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(trans_0_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(trans_0_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(trans_0_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(trans_0_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(trans_0_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(trans_0_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(trans_0_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(trans_0_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(trans_0_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(trans_0_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(trans_0_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(trans_0_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(trans_0_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(trans_0_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(trans_0_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(trans_0_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(trans_0_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(trans_0_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(trans_0_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(trans_0_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(trans_0_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(trans_0_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(trans_0_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(trans_0_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(trans_0_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(trans_0_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(trans_0_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(trans_0_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(trans_0_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(trans_0_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(trans_0_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(trans_0_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(trans_0_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(trans_0_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(trans_0_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(trans_0_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(trans_0_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(trans_0_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(trans_0_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(trans_0_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(trans_0_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(trans_0_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(trans_0_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(trans_0_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(trans_0_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(trans_0_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(trans_0_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(trans_0_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(trans_0_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(trans_0_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(trans_0_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(trans_0_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(trans_0_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(trans_0_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(trans_0_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(trans_0_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(trans_0_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(trans_0_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(trans_0_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(trans_0_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_out_data_0(trans_0_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(trans_0_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(trans_0_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(trans_0_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(trans_0_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(trans_0_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(trans_0_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(trans_0_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(trans_0_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(trans_0_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(trans_0_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(trans_0_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(trans_0_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(trans_0_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(trans_0_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(trans_0_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(trans_0_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(trans_0_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(trans_0_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(trans_0_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(trans_0_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(trans_0_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(trans_0_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(trans_0_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(trans_0_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(trans_0_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(trans_0_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(trans_0_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(trans_0_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(trans_0_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(trans_0_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(trans_0_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(trans_0_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(trans_0_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(trans_0_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(trans_0_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(trans_0_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(trans_0_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(trans_0_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(trans_0_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(trans_0_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(trans_0_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(trans_0_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(trans_0_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(trans_0_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(trans_0_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(trans_0_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(trans_0_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(trans_0_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(trans_0_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(trans_0_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(trans_0_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(trans_0_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(trans_0_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(trans_0_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(trans_0_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(trans_0_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(trans_0_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(trans_0_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(trans_0_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(trans_0_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(trans_0_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(trans_0_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(trans_0_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(trans_0_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(trans_0_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(trans_0_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(trans_0_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(trans_0_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(trans_0_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(trans_0_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(trans_0_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(trans_0_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(trans_0_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(trans_0_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(trans_0_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(trans_0_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(trans_0_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(trans_0_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(trans_0_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(trans_0_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(trans_0_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(trans_0_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(trans_0_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(trans_0_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(trans_0_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(trans_0_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(trans_0_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(trans_0_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(trans_0_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(trans_0_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(trans_0_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(trans_0_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(trans_0_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(trans_0_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(trans_0_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(trans_0_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(trans_0_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(trans_0_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(trans_0_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(trans_0_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(trans_0_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(trans_0_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(trans_0_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(trans_0_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(trans_0_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(trans_0_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(trans_0_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(trans_0_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(trans_0_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(trans_0_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(trans_0_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(trans_0_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(trans_0_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(trans_0_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(trans_0_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(trans_0_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(trans_0_io_pipe_phv_out_is_valid_processor),
    .io_next_proc_exist(trans_0_io_next_proc_exist),
    .io_next_proc_id(trans_0_io_next_proc_id)
  );
  InterProcessorTransfer trans_1 ( // @[ipsa.scala 79:25]
    .clock(trans_1_clock),
    .io_pipe_phv_in_data_0(trans_1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(trans_1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(trans_1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(trans_1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(trans_1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(trans_1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(trans_1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(trans_1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(trans_1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(trans_1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(trans_1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(trans_1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(trans_1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(trans_1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(trans_1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(trans_1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(trans_1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(trans_1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(trans_1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(trans_1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(trans_1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(trans_1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(trans_1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(trans_1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(trans_1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(trans_1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(trans_1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(trans_1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(trans_1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(trans_1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(trans_1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(trans_1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(trans_1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(trans_1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(trans_1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(trans_1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(trans_1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(trans_1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(trans_1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(trans_1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(trans_1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(trans_1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(trans_1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(trans_1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(trans_1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(trans_1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(trans_1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(trans_1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(trans_1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(trans_1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(trans_1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(trans_1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(trans_1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(trans_1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(trans_1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(trans_1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(trans_1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(trans_1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(trans_1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(trans_1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(trans_1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(trans_1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(trans_1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(trans_1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(trans_1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(trans_1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(trans_1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(trans_1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(trans_1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(trans_1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(trans_1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(trans_1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(trans_1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(trans_1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(trans_1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(trans_1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(trans_1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(trans_1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(trans_1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(trans_1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(trans_1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(trans_1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(trans_1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(trans_1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(trans_1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(trans_1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(trans_1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(trans_1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(trans_1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(trans_1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(trans_1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(trans_1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(trans_1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(trans_1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(trans_1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(trans_1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(trans_1_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(trans_1_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(trans_1_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(trans_1_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(trans_1_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(trans_1_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(trans_1_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(trans_1_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(trans_1_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(trans_1_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(trans_1_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(trans_1_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(trans_1_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(trans_1_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(trans_1_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(trans_1_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(trans_1_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(trans_1_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(trans_1_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(trans_1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(trans_1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_out_data_0(trans_1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(trans_1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(trans_1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(trans_1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(trans_1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(trans_1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(trans_1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(trans_1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(trans_1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(trans_1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(trans_1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(trans_1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(trans_1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(trans_1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(trans_1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(trans_1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(trans_1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(trans_1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(trans_1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(trans_1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(trans_1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(trans_1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(trans_1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(trans_1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(trans_1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(trans_1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(trans_1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(trans_1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(trans_1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(trans_1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(trans_1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(trans_1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(trans_1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(trans_1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(trans_1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(trans_1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(trans_1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(trans_1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(trans_1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(trans_1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(trans_1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(trans_1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(trans_1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(trans_1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(trans_1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(trans_1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(trans_1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(trans_1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(trans_1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(trans_1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(trans_1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(trans_1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(trans_1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(trans_1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(trans_1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(trans_1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(trans_1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(trans_1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(trans_1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(trans_1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(trans_1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(trans_1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(trans_1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(trans_1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(trans_1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(trans_1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(trans_1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(trans_1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(trans_1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(trans_1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(trans_1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(trans_1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(trans_1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(trans_1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(trans_1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(trans_1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(trans_1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(trans_1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(trans_1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(trans_1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(trans_1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(trans_1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(trans_1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(trans_1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(trans_1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(trans_1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(trans_1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(trans_1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(trans_1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(trans_1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(trans_1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(trans_1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(trans_1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(trans_1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(trans_1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(trans_1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(trans_1_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(trans_1_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(trans_1_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(trans_1_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(trans_1_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(trans_1_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(trans_1_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(trans_1_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(trans_1_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(trans_1_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(trans_1_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(trans_1_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(trans_1_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(trans_1_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(trans_1_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(trans_1_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(trans_1_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(trans_1_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(trans_1_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(trans_1_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(trans_1_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(trans_1_io_pipe_phv_out_is_valid_processor),
    .io_next_proc_exist(trans_1_io_next_proc_exist),
    .io_next_proc_id(trans_1_io_next_proc_id)
  );
  InterProcessorTransfer trans_2 ( // @[ipsa.scala 79:25]
    .clock(trans_2_clock),
    .io_pipe_phv_in_data_0(trans_2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(trans_2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(trans_2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(trans_2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(trans_2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(trans_2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(trans_2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(trans_2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(trans_2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(trans_2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(trans_2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(trans_2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(trans_2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(trans_2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(trans_2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(trans_2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(trans_2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(trans_2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(trans_2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(trans_2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(trans_2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(trans_2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(trans_2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(trans_2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(trans_2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(trans_2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(trans_2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(trans_2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(trans_2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(trans_2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(trans_2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(trans_2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(trans_2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(trans_2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(trans_2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(trans_2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(trans_2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(trans_2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(trans_2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(trans_2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(trans_2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(trans_2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(trans_2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(trans_2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(trans_2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(trans_2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(trans_2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(trans_2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(trans_2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(trans_2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(trans_2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(trans_2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(trans_2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(trans_2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(trans_2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(trans_2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(trans_2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(trans_2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(trans_2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(trans_2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(trans_2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(trans_2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(trans_2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(trans_2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(trans_2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(trans_2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(trans_2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(trans_2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(trans_2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(trans_2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(trans_2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(trans_2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(trans_2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(trans_2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(trans_2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(trans_2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(trans_2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(trans_2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(trans_2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(trans_2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(trans_2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(trans_2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(trans_2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(trans_2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(trans_2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(trans_2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(trans_2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(trans_2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(trans_2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(trans_2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(trans_2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(trans_2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(trans_2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(trans_2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(trans_2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(trans_2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(trans_2_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(trans_2_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(trans_2_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(trans_2_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(trans_2_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(trans_2_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(trans_2_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(trans_2_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(trans_2_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(trans_2_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(trans_2_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(trans_2_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(trans_2_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(trans_2_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(trans_2_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(trans_2_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(trans_2_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(trans_2_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(trans_2_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(trans_2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(trans_2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_out_data_0(trans_2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(trans_2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(trans_2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(trans_2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(trans_2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(trans_2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(trans_2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(trans_2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(trans_2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(trans_2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(trans_2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(trans_2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(trans_2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(trans_2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(trans_2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(trans_2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(trans_2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(trans_2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(trans_2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(trans_2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(trans_2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(trans_2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(trans_2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(trans_2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(trans_2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(trans_2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(trans_2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(trans_2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(trans_2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(trans_2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(trans_2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(trans_2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(trans_2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(trans_2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(trans_2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(trans_2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(trans_2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(trans_2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(trans_2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(trans_2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(trans_2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(trans_2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(trans_2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(trans_2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(trans_2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(trans_2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(trans_2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(trans_2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(trans_2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(trans_2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(trans_2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(trans_2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(trans_2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(trans_2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(trans_2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(trans_2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(trans_2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(trans_2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(trans_2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(trans_2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(trans_2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(trans_2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(trans_2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(trans_2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(trans_2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(trans_2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(trans_2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(trans_2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(trans_2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(trans_2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(trans_2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(trans_2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(trans_2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(trans_2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(trans_2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(trans_2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(trans_2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(trans_2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(trans_2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(trans_2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(trans_2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(trans_2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(trans_2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(trans_2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(trans_2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(trans_2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(trans_2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(trans_2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(trans_2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(trans_2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(trans_2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(trans_2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(trans_2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(trans_2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(trans_2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(trans_2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(trans_2_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(trans_2_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(trans_2_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(trans_2_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(trans_2_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(trans_2_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(trans_2_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(trans_2_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(trans_2_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(trans_2_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(trans_2_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(trans_2_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(trans_2_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(trans_2_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(trans_2_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(trans_2_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(trans_2_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(trans_2_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(trans_2_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(trans_2_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(trans_2_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(trans_2_io_pipe_phv_out_is_valid_processor),
    .io_next_proc_exist(trans_2_io_next_proc_exist),
    .io_next_proc_id(trans_2_io_next_proc_id)
  );
  InterProcessorTransfer trans_3 ( // @[ipsa.scala 79:25]
    .clock(trans_3_clock),
    .io_pipe_phv_in_data_0(trans_3_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(trans_3_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(trans_3_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(trans_3_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(trans_3_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(trans_3_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(trans_3_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(trans_3_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(trans_3_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(trans_3_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(trans_3_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(trans_3_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(trans_3_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(trans_3_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(trans_3_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(trans_3_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(trans_3_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(trans_3_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(trans_3_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(trans_3_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(trans_3_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(trans_3_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(trans_3_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(trans_3_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(trans_3_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(trans_3_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(trans_3_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(trans_3_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(trans_3_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(trans_3_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(trans_3_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(trans_3_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(trans_3_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(trans_3_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(trans_3_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(trans_3_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(trans_3_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(trans_3_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(trans_3_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(trans_3_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(trans_3_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(trans_3_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(trans_3_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(trans_3_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(trans_3_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(trans_3_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(trans_3_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(trans_3_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(trans_3_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(trans_3_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(trans_3_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(trans_3_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(trans_3_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(trans_3_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(trans_3_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(trans_3_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(trans_3_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(trans_3_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(trans_3_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(trans_3_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(trans_3_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(trans_3_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(trans_3_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(trans_3_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(trans_3_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(trans_3_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(trans_3_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(trans_3_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(trans_3_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(trans_3_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(trans_3_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(trans_3_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(trans_3_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(trans_3_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(trans_3_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(trans_3_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(trans_3_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(trans_3_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(trans_3_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(trans_3_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(trans_3_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(trans_3_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(trans_3_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(trans_3_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(trans_3_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(trans_3_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(trans_3_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(trans_3_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(trans_3_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(trans_3_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(trans_3_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(trans_3_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(trans_3_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(trans_3_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(trans_3_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(trans_3_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(trans_3_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(trans_3_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(trans_3_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(trans_3_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(trans_3_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(trans_3_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(trans_3_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(trans_3_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(trans_3_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(trans_3_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(trans_3_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(trans_3_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(trans_3_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(trans_3_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(trans_3_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(trans_3_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(trans_3_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(trans_3_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(trans_3_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(trans_3_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(trans_3_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_out_data_0(trans_3_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(trans_3_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(trans_3_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(trans_3_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(trans_3_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(trans_3_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(trans_3_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(trans_3_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(trans_3_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(trans_3_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(trans_3_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(trans_3_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(trans_3_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(trans_3_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(trans_3_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(trans_3_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(trans_3_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(trans_3_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(trans_3_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(trans_3_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(trans_3_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(trans_3_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(trans_3_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(trans_3_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(trans_3_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(trans_3_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(trans_3_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(trans_3_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(trans_3_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(trans_3_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(trans_3_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(trans_3_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(trans_3_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(trans_3_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(trans_3_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(trans_3_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(trans_3_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(trans_3_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(trans_3_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(trans_3_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(trans_3_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(trans_3_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(trans_3_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(trans_3_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(trans_3_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(trans_3_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(trans_3_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(trans_3_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(trans_3_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(trans_3_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(trans_3_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(trans_3_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(trans_3_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(trans_3_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(trans_3_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(trans_3_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(trans_3_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(trans_3_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(trans_3_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(trans_3_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(trans_3_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(trans_3_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(trans_3_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(trans_3_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(trans_3_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(trans_3_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(trans_3_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(trans_3_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(trans_3_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(trans_3_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(trans_3_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(trans_3_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(trans_3_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(trans_3_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(trans_3_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(trans_3_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(trans_3_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(trans_3_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(trans_3_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(trans_3_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(trans_3_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(trans_3_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(trans_3_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(trans_3_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(trans_3_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(trans_3_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(trans_3_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(trans_3_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(trans_3_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(trans_3_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(trans_3_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(trans_3_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(trans_3_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(trans_3_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(trans_3_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(trans_3_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(trans_3_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(trans_3_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(trans_3_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(trans_3_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(trans_3_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(trans_3_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(trans_3_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(trans_3_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(trans_3_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(trans_3_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(trans_3_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(trans_3_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(trans_3_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(trans_3_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(trans_3_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(trans_3_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(trans_3_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(trans_3_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(trans_3_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(trans_3_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(trans_3_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(trans_3_io_pipe_phv_out_is_valid_processor),
    .io_next_proc_exist(trans_3_io_next_proc_exist),
    .io_next_proc_id(trans_3_io_next_proc_id)
  );
  assign io_pipe_phv_out_data_0 = 2'h3 != last_proc_id ? _GEN_3096 : trans_3_io_pipe_phv_out_data_0; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_1 = 2'h3 != last_proc_id ? _GEN_3097 : trans_3_io_pipe_phv_out_data_1; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_2 = 2'h3 != last_proc_id ? _GEN_3098 : trans_3_io_pipe_phv_out_data_2; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_3 = 2'h3 != last_proc_id ? _GEN_3099 : trans_3_io_pipe_phv_out_data_3; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_4 = 2'h3 != last_proc_id ? _GEN_3100 : trans_3_io_pipe_phv_out_data_4; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_5 = 2'h3 != last_proc_id ? _GEN_3101 : trans_3_io_pipe_phv_out_data_5; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_6 = 2'h3 != last_proc_id ? _GEN_3102 : trans_3_io_pipe_phv_out_data_6; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_7 = 2'h3 != last_proc_id ? _GEN_3103 : trans_3_io_pipe_phv_out_data_7; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_8 = 2'h3 != last_proc_id ? _GEN_3104 : trans_3_io_pipe_phv_out_data_8; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_9 = 2'h3 != last_proc_id ? _GEN_3105 : trans_3_io_pipe_phv_out_data_9; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_10 = 2'h3 != last_proc_id ? _GEN_3106 : trans_3_io_pipe_phv_out_data_10; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_11 = 2'h3 != last_proc_id ? _GEN_3107 : trans_3_io_pipe_phv_out_data_11; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_12 = 2'h3 != last_proc_id ? _GEN_3108 : trans_3_io_pipe_phv_out_data_12; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_13 = 2'h3 != last_proc_id ? _GEN_3109 : trans_3_io_pipe_phv_out_data_13; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_14 = 2'h3 != last_proc_id ? _GEN_3110 : trans_3_io_pipe_phv_out_data_14; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_15 = 2'h3 != last_proc_id ? _GEN_3111 : trans_3_io_pipe_phv_out_data_15; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_16 = 2'h3 != last_proc_id ? _GEN_3112 : trans_3_io_pipe_phv_out_data_16; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_17 = 2'h3 != last_proc_id ? _GEN_3113 : trans_3_io_pipe_phv_out_data_17; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_18 = 2'h3 != last_proc_id ? _GEN_3114 : trans_3_io_pipe_phv_out_data_18; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_19 = 2'h3 != last_proc_id ? _GEN_3115 : trans_3_io_pipe_phv_out_data_19; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_20 = 2'h3 != last_proc_id ? _GEN_3116 : trans_3_io_pipe_phv_out_data_20; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_21 = 2'h3 != last_proc_id ? _GEN_3117 : trans_3_io_pipe_phv_out_data_21; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_22 = 2'h3 != last_proc_id ? _GEN_3118 : trans_3_io_pipe_phv_out_data_22; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_23 = 2'h3 != last_proc_id ? _GEN_3119 : trans_3_io_pipe_phv_out_data_23; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_24 = 2'h3 != last_proc_id ? _GEN_3120 : trans_3_io_pipe_phv_out_data_24; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_25 = 2'h3 != last_proc_id ? _GEN_3121 : trans_3_io_pipe_phv_out_data_25; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_26 = 2'h3 != last_proc_id ? _GEN_3122 : trans_3_io_pipe_phv_out_data_26; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_27 = 2'h3 != last_proc_id ? _GEN_3123 : trans_3_io_pipe_phv_out_data_27; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_28 = 2'h3 != last_proc_id ? _GEN_3124 : trans_3_io_pipe_phv_out_data_28; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_29 = 2'h3 != last_proc_id ? _GEN_3125 : trans_3_io_pipe_phv_out_data_29; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_30 = 2'h3 != last_proc_id ? _GEN_3126 : trans_3_io_pipe_phv_out_data_30; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_31 = 2'h3 != last_proc_id ? _GEN_3127 : trans_3_io_pipe_phv_out_data_31; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_32 = 2'h3 != last_proc_id ? _GEN_3128 : trans_3_io_pipe_phv_out_data_32; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_33 = 2'h3 != last_proc_id ? _GEN_3129 : trans_3_io_pipe_phv_out_data_33; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_34 = 2'h3 != last_proc_id ? _GEN_3130 : trans_3_io_pipe_phv_out_data_34; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_35 = 2'h3 != last_proc_id ? _GEN_3131 : trans_3_io_pipe_phv_out_data_35; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_36 = 2'h3 != last_proc_id ? _GEN_3132 : trans_3_io_pipe_phv_out_data_36; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_37 = 2'h3 != last_proc_id ? _GEN_3133 : trans_3_io_pipe_phv_out_data_37; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_38 = 2'h3 != last_proc_id ? _GEN_3134 : trans_3_io_pipe_phv_out_data_38; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_39 = 2'h3 != last_proc_id ? _GEN_3135 : trans_3_io_pipe_phv_out_data_39; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_40 = 2'h3 != last_proc_id ? _GEN_3136 : trans_3_io_pipe_phv_out_data_40; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_41 = 2'h3 != last_proc_id ? _GEN_3137 : trans_3_io_pipe_phv_out_data_41; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_42 = 2'h3 != last_proc_id ? _GEN_3138 : trans_3_io_pipe_phv_out_data_42; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_43 = 2'h3 != last_proc_id ? _GEN_3139 : trans_3_io_pipe_phv_out_data_43; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_44 = 2'h3 != last_proc_id ? _GEN_3140 : trans_3_io_pipe_phv_out_data_44; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_45 = 2'h3 != last_proc_id ? _GEN_3141 : trans_3_io_pipe_phv_out_data_45; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_46 = 2'h3 != last_proc_id ? _GEN_3142 : trans_3_io_pipe_phv_out_data_46; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_47 = 2'h3 != last_proc_id ? _GEN_3143 : trans_3_io_pipe_phv_out_data_47; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_48 = 2'h3 != last_proc_id ? _GEN_3144 : trans_3_io_pipe_phv_out_data_48; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_49 = 2'h3 != last_proc_id ? _GEN_3145 : trans_3_io_pipe_phv_out_data_49; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_50 = 2'h3 != last_proc_id ? _GEN_3146 : trans_3_io_pipe_phv_out_data_50; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_51 = 2'h3 != last_proc_id ? _GEN_3147 : trans_3_io_pipe_phv_out_data_51; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_52 = 2'h3 != last_proc_id ? _GEN_3148 : trans_3_io_pipe_phv_out_data_52; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_53 = 2'h3 != last_proc_id ? _GEN_3149 : trans_3_io_pipe_phv_out_data_53; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_54 = 2'h3 != last_proc_id ? _GEN_3150 : trans_3_io_pipe_phv_out_data_54; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_55 = 2'h3 != last_proc_id ? _GEN_3151 : trans_3_io_pipe_phv_out_data_55; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_56 = 2'h3 != last_proc_id ? _GEN_3152 : trans_3_io_pipe_phv_out_data_56; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_57 = 2'h3 != last_proc_id ? _GEN_3153 : trans_3_io_pipe_phv_out_data_57; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_58 = 2'h3 != last_proc_id ? _GEN_3154 : trans_3_io_pipe_phv_out_data_58; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_59 = 2'h3 != last_proc_id ? _GEN_3155 : trans_3_io_pipe_phv_out_data_59; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_60 = 2'h3 != last_proc_id ? _GEN_3156 : trans_3_io_pipe_phv_out_data_60; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_61 = 2'h3 != last_proc_id ? _GEN_3157 : trans_3_io_pipe_phv_out_data_61; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_62 = 2'h3 != last_proc_id ? _GEN_3158 : trans_3_io_pipe_phv_out_data_62; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_63 = 2'h3 != last_proc_id ? _GEN_3159 : trans_3_io_pipe_phv_out_data_63; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_64 = 2'h3 != last_proc_id ? _GEN_3160 : trans_3_io_pipe_phv_out_data_64; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_65 = 2'h3 != last_proc_id ? _GEN_3161 : trans_3_io_pipe_phv_out_data_65; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_66 = 2'h3 != last_proc_id ? _GEN_3162 : trans_3_io_pipe_phv_out_data_66; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_67 = 2'h3 != last_proc_id ? _GEN_3163 : trans_3_io_pipe_phv_out_data_67; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_68 = 2'h3 != last_proc_id ? _GEN_3164 : trans_3_io_pipe_phv_out_data_68; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_69 = 2'h3 != last_proc_id ? _GEN_3165 : trans_3_io_pipe_phv_out_data_69; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_70 = 2'h3 != last_proc_id ? _GEN_3166 : trans_3_io_pipe_phv_out_data_70; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_71 = 2'h3 != last_proc_id ? _GEN_3167 : trans_3_io_pipe_phv_out_data_71; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_72 = 2'h3 != last_proc_id ? _GEN_3168 : trans_3_io_pipe_phv_out_data_72; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_73 = 2'h3 != last_proc_id ? _GEN_3169 : trans_3_io_pipe_phv_out_data_73; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_74 = 2'h3 != last_proc_id ? _GEN_3170 : trans_3_io_pipe_phv_out_data_74; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_75 = 2'h3 != last_proc_id ? _GEN_3171 : trans_3_io_pipe_phv_out_data_75; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_76 = 2'h3 != last_proc_id ? _GEN_3172 : trans_3_io_pipe_phv_out_data_76; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_77 = 2'h3 != last_proc_id ? _GEN_3173 : trans_3_io_pipe_phv_out_data_77; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_78 = 2'h3 != last_proc_id ? _GEN_3174 : trans_3_io_pipe_phv_out_data_78; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_79 = 2'h3 != last_proc_id ? _GEN_3175 : trans_3_io_pipe_phv_out_data_79; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_80 = 2'h3 != last_proc_id ? _GEN_3176 : trans_3_io_pipe_phv_out_data_80; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_81 = 2'h3 != last_proc_id ? _GEN_3177 : trans_3_io_pipe_phv_out_data_81; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_82 = 2'h3 != last_proc_id ? _GEN_3178 : trans_3_io_pipe_phv_out_data_82; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_83 = 2'h3 != last_proc_id ? _GEN_3179 : trans_3_io_pipe_phv_out_data_83; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_84 = 2'h3 != last_proc_id ? _GEN_3180 : trans_3_io_pipe_phv_out_data_84; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_85 = 2'h3 != last_proc_id ? _GEN_3181 : trans_3_io_pipe_phv_out_data_85; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_86 = 2'h3 != last_proc_id ? _GEN_3182 : trans_3_io_pipe_phv_out_data_86; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_87 = 2'h3 != last_proc_id ? _GEN_3183 : trans_3_io_pipe_phv_out_data_87; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_88 = 2'h3 != last_proc_id ? _GEN_3184 : trans_3_io_pipe_phv_out_data_88; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_89 = 2'h3 != last_proc_id ? _GEN_3185 : trans_3_io_pipe_phv_out_data_89; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_90 = 2'h3 != last_proc_id ? _GEN_3186 : trans_3_io_pipe_phv_out_data_90; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_91 = 2'h3 != last_proc_id ? _GEN_3187 : trans_3_io_pipe_phv_out_data_91; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_92 = 2'h3 != last_proc_id ? _GEN_3188 : trans_3_io_pipe_phv_out_data_92; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_93 = 2'h3 != last_proc_id ? _GEN_3189 : trans_3_io_pipe_phv_out_data_93; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_94 = 2'h3 != last_proc_id ? _GEN_3190 : trans_3_io_pipe_phv_out_data_94; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_data_95 = 2'h3 != last_proc_id ? _GEN_3191 : trans_3_io_pipe_phv_out_data_95; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_header_0 = 2'h3 != last_proc_id ? _GEN_3080 : trans_3_io_pipe_phv_out_header_0; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_header_1 = 2'h3 != last_proc_id ? _GEN_3081 : trans_3_io_pipe_phv_out_header_1; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_header_2 = 2'h3 != last_proc_id ? _GEN_3082 : trans_3_io_pipe_phv_out_header_2; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_header_3 = 2'h3 != last_proc_id ? _GEN_3083 : trans_3_io_pipe_phv_out_header_3; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_header_4 = 2'h3 != last_proc_id ? _GEN_3084 : trans_3_io_pipe_phv_out_header_4; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_header_5 = 2'h3 != last_proc_id ? _GEN_3085 : trans_3_io_pipe_phv_out_header_5; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_header_6 = 2'h3 != last_proc_id ? _GEN_3086 : trans_3_io_pipe_phv_out_header_6; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_header_7 = 2'h3 != last_proc_id ? _GEN_3087 : trans_3_io_pipe_phv_out_header_7; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_header_8 = 2'h3 != last_proc_id ? _GEN_3088 : trans_3_io_pipe_phv_out_header_8; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_header_9 = 2'h3 != last_proc_id ? _GEN_3089 : trans_3_io_pipe_phv_out_header_9; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_header_10 = 2'h3 != last_proc_id ? _GEN_3090 : trans_3_io_pipe_phv_out_header_10; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_header_11 = 2'h3 != last_proc_id ? _GEN_3091 : trans_3_io_pipe_phv_out_header_11; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_header_12 = 2'h3 != last_proc_id ? _GEN_3092 : trans_3_io_pipe_phv_out_header_12; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_header_13 = 2'h3 != last_proc_id ? _GEN_3093 : trans_3_io_pipe_phv_out_header_13; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_header_14 = 2'h3 != last_proc_id ? _GEN_3094 : trans_3_io_pipe_phv_out_header_14; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_header_15 = 2'h3 != last_proc_id ? _GEN_3095 : trans_3_io_pipe_phv_out_header_15; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_parse_current_state = 2'h3 != last_proc_id ? _GEN_3079 :
    trans_3_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_parse_current_offset = 2'h3 != last_proc_id ? _GEN_3078 :
    trans_3_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_parse_transition_field = 2'h3 != last_proc_id ? _GEN_3077 :
    trans_3_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_next_processor_id = 2'h3 != last_proc_id ? _GEN_3076 :
    trans_3_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_next_config_id = 2'h3 != last_proc_id ? _GEN_3075 : trans_3_io_pipe_phv_out_next_config_id; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign io_pipe_phv_out_is_valid_processor = 2'h3 != last_proc_id ? _GEN_3074 :
    trans_3_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 94:65 ipsa.scala 101:29]
  assign proc_0_clock = clock;
  assign proc_0_io_pipe_phv_in_data_0 = 2'h3 != last_proc_id ? _GEN_3214 : _GEN_2624; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_1 = 2'h3 != last_proc_id ? _GEN_3215 : _GEN_2625; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_2 = 2'h3 != last_proc_id ? _GEN_3216 : _GEN_2626; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_3 = 2'h3 != last_proc_id ? _GEN_3217 : _GEN_2627; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_4 = 2'h3 != last_proc_id ? _GEN_3218 : _GEN_2628; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_5 = 2'h3 != last_proc_id ? _GEN_3219 : _GEN_2629; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_6 = 2'h3 != last_proc_id ? _GEN_3220 : _GEN_2630; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_7 = 2'h3 != last_proc_id ? _GEN_3221 : _GEN_2631; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_8 = 2'h3 != last_proc_id ? _GEN_3222 : _GEN_2632; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_9 = 2'h3 != last_proc_id ? _GEN_3223 : _GEN_2633; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_10 = 2'h3 != last_proc_id ? _GEN_3224 : _GEN_2634; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_11 = 2'h3 != last_proc_id ? _GEN_3225 : _GEN_2635; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_12 = 2'h3 != last_proc_id ? _GEN_3226 : _GEN_2636; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_13 = 2'h3 != last_proc_id ? _GEN_3227 : _GEN_2637; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_14 = 2'h3 != last_proc_id ? _GEN_3228 : _GEN_2638; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_15 = 2'h3 != last_proc_id ? _GEN_3229 : _GEN_2639; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_16 = 2'h3 != last_proc_id ? _GEN_3230 : _GEN_2640; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_17 = 2'h3 != last_proc_id ? _GEN_3231 : _GEN_2641; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_18 = 2'h3 != last_proc_id ? _GEN_3232 : _GEN_2642; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_19 = 2'h3 != last_proc_id ? _GEN_3233 : _GEN_2643; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_20 = 2'h3 != last_proc_id ? _GEN_3234 : _GEN_2644; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_21 = 2'h3 != last_proc_id ? _GEN_3235 : _GEN_2645; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_22 = 2'h3 != last_proc_id ? _GEN_3236 : _GEN_2646; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_23 = 2'h3 != last_proc_id ? _GEN_3237 : _GEN_2647; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_24 = 2'h3 != last_proc_id ? _GEN_3238 : _GEN_2648; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_25 = 2'h3 != last_proc_id ? _GEN_3239 : _GEN_2649; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_26 = 2'h3 != last_proc_id ? _GEN_3240 : _GEN_2650; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_27 = 2'h3 != last_proc_id ? _GEN_3241 : _GEN_2651; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_28 = 2'h3 != last_proc_id ? _GEN_3242 : _GEN_2652; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_29 = 2'h3 != last_proc_id ? _GEN_3243 : _GEN_2653; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_30 = 2'h3 != last_proc_id ? _GEN_3244 : _GEN_2654; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_31 = 2'h3 != last_proc_id ? _GEN_3245 : _GEN_2655; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_32 = 2'h3 != last_proc_id ? _GEN_3246 : _GEN_2656; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_33 = 2'h3 != last_proc_id ? _GEN_3247 : _GEN_2657; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_34 = 2'h3 != last_proc_id ? _GEN_3248 : _GEN_2658; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_35 = 2'h3 != last_proc_id ? _GEN_3249 : _GEN_2659; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_36 = 2'h3 != last_proc_id ? _GEN_3250 : _GEN_2660; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_37 = 2'h3 != last_proc_id ? _GEN_3251 : _GEN_2661; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_38 = 2'h3 != last_proc_id ? _GEN_3252 : _GEN_2662; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_39 = 2'h3 != last_proc_id ? _GEN_3253 : _GEN_2663; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_40 = 2'h3 != last_proc_id ? _GEN_3254 : _GEN_2664; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_41 = 2'h3 != last_proc_id ? _GEN_3255 : _GEN_2665; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_42 = 2'h3 != last_proc_id ? _GEN_3256 : _GEN_2666; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_43 = 2'h3 != last_proc_id ? _GEN_3257 : _GEN_2667; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_44 = 2'h3 != last_proc_id ? _GEN_3258 : _GEN_2668; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_45 = 2'h3 != last_proc_id ? _GEN_3259 : _GEN_2669; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_46 = 2'h3 != last_proc_id ? _GEN_3260 : _GEN_2670; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_47 = 2'h3 != last_proc_id ? _GEN_3261 : _GEN_2671; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_48 = 2'h3 != last_proc_id ? _GEN_3262 : _GEN_2672; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_49 = 2'h3 != last_proc_id ? _GEN_3263 : _GEN_2673; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_50 = 2'h3 != last_proc_id ? _GEN_3264 : _GEN_2674; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_51 = 2'h3 != last_proc_id ? _GEN_3265 : _GEN_2675; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_52 = 2'h3 != last_proc_id ? _GEN_3266 : _GEN_2676; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_53 = 2'h3 != last_proc_id ? _GEN_3267 : _GEN_2677; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_54 = 2'h3 != last_proc_id ? _GEN_3268 : _GEN_2678; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_55 = 2'h3 != last_proc_id ? _GEN_3269 : _GEN_2679; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_56 = 2'h3 != last_proc_id ? _GEN_3270 : _GEN_2680; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_57 = 2'h3 != last_proc_id ? _GEN_3271 : _GEN_2681; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_58 = 2'h3 != last_proc_id ? _GEN_3272 : _GEN_2682; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_59 = 2'h3 != last_proc_id ? _GEN_3273 : _GEN_2683; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_60 = 2'h3 != last_proc_id ? _GEN_3274 : _GEN_2684; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_61 = 2'h3 != last_proc_id ? _GEN_3275 : _GEN_2685; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_62 = 2'h3 != last_proc_id ? _GEN_3276 : _GEN_2686; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_63 = 2'h3 != last_proc_id ? _GEN_3277 : _GEN_2687; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_64 = 2'h3 != last_proc_id ? _GEN_3278 : _GEN_2688; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_65 = 2'h3 != last_proc_id ? _GEN_3279 : _GEN_2689; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_66 = 2'h3 != last_proc_id ? _GEN_3280 : _GEN_2690; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_67 = 2'h3 != last_proc_id ? _GEN_3281 : _GEN_2691; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_68 = 2'h3 != last_proc_id ? _GEN_3282 : _GEN_2692; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_69 = 2'h3 != last_proc_id ? _GEN_3283 : _GEN_2693; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_70 = 2'h3 != last_proc_id ? _GEN_3284 : _GEN_2694; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_71 = 2'h3 != last_proc_id ? _GEN_3285 : _GEN_2695; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_72 = 2'h3 != last_proc_id ? _GEN_3286 : _GEN_2696; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_73 = 2'h3 != last_proc_id ? _GEN_3287 : _GEN_2697; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_74 = 2'h3 != last_proc_id ? _GEN_3288 : _GEN_2698; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_75 = 2'h3 != last_proc_id ? _GEN_3289 : _GEN_2699; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_76 = 2'h3 != last_proc_id ? _GEN_3290 : _GEN_2700; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_77 = 2'h3 != last_proc_id ? _GEN_3291 : _GEN_2701; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_78 = 2'h3 != last_proc_id ? _GEN_3292 : _GEN_2702; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_79 = 2'h3 != last_proc_id ? _GEN_3293 : _GEN_2703; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_80 = 2'h3 != last_proc_id ? _GEN_3294 : _GEN_2704; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_81 = 2'h3 != last_proc_id ? _GEN_3295 : _GEN_2705; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_82 = 2'h3 != last_proc_id ? _GEN_3296 : _GEN_2706; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_83 = 2'h3 != last_proc_id ? _GEN_3297 : _GEN_2707; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_84 = 2'h3 != last_proc_id ? _GEN_3298 : _GEN_2708; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_85 = 2'h3 != last_proc_id ? _GEN_3299 : _GEN_2709; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_86 = 2'h3 != last_proc_id ? _GEN_3300 : _GEN_2710; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_87 = 2'h3 != last_proc_id ? _GEN_3301 : _GEN_2711; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_88 = 2'h3 != last_proc_id ? _GEN_3302 : _GEN_2712; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_89 = 2'h3 != last_proc_id ? _GEN_3303 : _GEN_2713; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_90 = 2'h3 != last_proc_id ? _GEN_3304 : _GEN_2714; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_91 = 2'h3 != last_proc_id ? _GEN_3305 : _GEN_2715; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_92 = 2'h3 != last_proc_id ? _GEN_3306 : _GEN_2716; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_93 = 2'h3 != last_proc_id ? _GEN_3307 : _GEN_2717; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_94 = 2'h3 != last_proc_id ? _GEN_3308 : _GEN_2718; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_data_95 = 2'h3 != last_proc_id ? _GEN_3309 : _GEN_2719; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_header_0 = 2'h3 != last_proc_id ? _GEN_3198 : _GEN_2608; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_header_1 = 2'h3 != last_proc_id ? _GEN_3199 : _GEN_2609; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_header_2 = 2'h3 != last_proc_id ? _GEN_3200 : _GEN_2610; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_header_3 = 2'h3 != last_proc_id ? _GEN_3201 : _GEN_2611; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_header_4 = 2'h3 != last_proc_id ? _GEN_3202 : _GEN_2612; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_header_5 = 2'h3 != last_proc_id ? _GEN_3203 : _GEN_2613; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_header_6 = 2'h3 != last_proc_id ? _GEN_3204 : _GEN_2614; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_header_7 = 2'h3 != last_proc_id ? _GEN_3205 : _GEN_2615; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_header_8 = 2'h3 != last_proc_id ? _GEN_3206 : _GEN_2616; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_header_9 = 2'h3 != last_proc_id ? _GEN_3207 : _GEN_2617; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_header_10 = 2'h3 != last_proc_id ? _GEN_3208 : _GEN_2618; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_header_11 = 2'h3 != last_proc_id ? _GEN_3209 : _GEN_2619; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_header_12 = 2'h3 != last_proc_id ? _GEN_3210 : _GEN_2620; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_header_13 = 2'h3 != last_proc_id ? _GEN_3211 : _GEN_2621; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_header_14 = 2'h3 != last_proc_id ? _GEN_3212 : _GEN_2622; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_header_15 = 2'h3 != last_proc_id ? _GEN_3213 : _GEN_2623; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_parse_current_state = 2'h3 != last_proc_id ? _GEN_3197 : _GEN_2607; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_parse_current_offset = 2'h3 != last_proc_id ? _GEN_3196 : _GEN_2606; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_parse_transition_field = 2'h3 != last_proc_id ? _GEN_3195 : _GEN_2605; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_next_processor_id = 2'h3 != last_proc_id ? _GEN_3194 : _GEN_2604; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_next_config_id = 2'h3 != last_proc_id ? _GEN_3193 : _GEN_2603; // @[ipsa.scala 94:65]
  assign proc_0_io_pipe_phv_in_is_valid_processor = 2'h3 != last_proc_id ? _GEN_3192 : _GEN_2602; // @[ipsa.scala 94:65]
  assign proc_0_io_mod_par_mod_en = io_mod_proc_mod_0_par_mod_en; // @[ipsa.scala 57:20]
  assign proc_0_io_mod_par_mod_last_mau_id_mod = io_mod_proc_mod_0_par_mod_last_mau_id_mod; // @[ipsa.scala 57:20]
  assign proc_0_io_mod_par_mod_last_mau_id = io_mod_proc_mod_0_par_mod_last_mau_id; // @[ipsa.scala 57:20]
  assign proc_0_io_mod_par_mod_cs = io_mod_proc_mod_0_par_mod_cs; // @[ipsa.scala 57:20]
  assign proc_0_io_mod_par_mod_module_mod_state_id_mod = io_mod_proc_mod_0_par_mod_module_mod_state_id_mod; // @[ipsa.scala 57:20]
  assign proc_0_io_mod_par_mod_module_mod_state_id = io_mod_proc_mod_0_par_mod_module_mod_state_id; // @[ipsa.scala 57:20]
  assign proc_0_io_mod_par_mod_module_mod_sram_w_cs = io_mod_proc_mod_0_par_mod_module_mod_sram_w_cs; // @[ipsa.scala 57:20]
  assign proc_0_io_mod_par_mod_module_mod_sram_w_addr = io_mod_proc_mod_0_par_mod_module_mod_sram_w_addr; // @[ipsa.scala 57:20]
  assign proc_0_io_mod_par_mod_module_mod_sram_w_data = io_mod_proc_mod_0_par_mod_module_mod_sram_w_data; // @[ipsa.scala 57:20]
  assign proc_0_io_mod_mat_mod_en = io_mod_proc_mod_0_mat_mod_en; // @[ipsa.scala 57:20]
  assign proc_0_io_mod_mat_mod_config_id = io_mod_proc_mod_0_mat_mod_config_id; // @[ipsa.scala 57:20]
  assign proc_0_io_mod_mat_mod_key_mod_header_id = io_mod_proc_mod_0_mat_mod_key_mod_header_id; // @[ipsa.scala 57:20]
  assign proc_0_io_mod_mat_mod_key_mod_internal_offset = io_mod_proc_mod_0_mat_mod_key_mod_internal_offset; // @[ipsa.scala 57:20]
  assign proc_0_io_mod_mat_mod_key_mod_key_length = io_mod_proc_mod_0_mat_mod_key_mod_key_length; // @[ipsa.scala 57:20]
  assign proc_0_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_0_mat_mod_table_mod_table_width; // @[ipsa.scala 57:20]
  assign proc_0_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_0_mat_mod_table_mod_table_depth; // @[ipsa.scala 57:20]
  assign proc_0_io_mod_act_mod_en = io_mod_proc_mod_0_act_mod_en; // @[ipsa.scala 57:20]
  assign proc_0_io_mod_act_mod_addr = io_mod_proc_mod_0_act_mod_addr; // @[ipsa.scala 57:20]
  assign proc_0_io_mod_act_mod_data_0 = io_mod_proc_mod_0_act_mod_data_0; // @[ipsa.scala 57:20]
  assign proc_0_io_mod_act_mod_data_1 = io_mod_proc_mod_0_act_mod_data_1; // @[ipsa.scala 57:20]
  assign proc_0_io_mem_cluster_0_data = sram_cluster_0_io_r_0_cluster_0_data; // @[ipsa.scala 70:37]
  assign proc_0_io_mem_cluster_1_data = sram_cluster_0_io_r_0_cluster_1_data; // @[ipsa.scala 70:37]
  assign proc_0_io_mem_cluster_2_data = sram_cluster_0_io_r_0_cluster_2_data; // @[ipsa.scala 70:37]
  assign proc_0_io_mem_cluster_3_data = sram_cluster_0_io_r_0_cluster_3_data; // @[ipsa.scala 70:37]
  assign proc_0_io_mem_cluster_4_data = sram_cluster_0_io_r_0_cluster_4_data; // @[ipsa.scala 70:37]
  assign proc_0_io_mem_cluster_5_data = sram_cluster_0_io_r_0_cluster_5_data; // @[ipsa.scala 70:37]
  assign proc_0_io_mem_cluster_6_data = sram_cluster_0_io_r_0_cluster_6_data; // @[ipsa.scala 70:37]
  assign proc_0_io_mem_cluster_7_data = sram_cluster_0_io_r_0_cluster_7_data; // @[ipsa.scala 70:37]
  assign proc_1_clock = clock;
  assign proc_1_io_pipe_phv_in_data_0 = 2'h3 != last_proc_id ? _GEN_3332 : _GEN_2742; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_1 = 2'h3 != last_proc_id ? _GEN_3333 : _GEN_2743; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_2 = 2'h3 != last_proc_id ? _GEN_3334 : _GEN_2744; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_3 = 2'h3 != last_proc_id ? _GEN_3335 : _GEN_2745; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_4 = 2'h3 != last_proc_id ? _GEN_3336 : _GEN_2746; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_5 = 2'h3 != last_proc_id ? _GEN_3337 : _GEN_2747; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_6 = 2'h3 != last_proc_id ? _GEN_3338 : _GEN_2748; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_7 = 2'h3 != last_proc_id ? _GEN_3339 : _GEN_2749; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_8 = 2'h3 != last_proc_id ? _GEN_3340 : _GEN_2750; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_9 = 2'h3 != last_proc_id ? _GEN_3341 : _GEN_2751; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_10 = 2'h3 != last_proc_id ? _GEN_3342 : _GEN_2752; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_11 = 2'h3 != last_proc_id ? _GEN_3343 : _GEN_2753; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_12 = 2'h3 != last_proc_id ? _GEN_3344 : _GEN_2754; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_13 = 2'h3 != last_proc_id ? _GEN_3345 : _GEN_2755; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_14 = 2'h3 != last_proc_id ? _GEN_3346 : _GEN_2756; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_15 = 2'h3 != last_proc_id ? _GEN_3347 : _GEN_2757; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_16 = 2'h3 != last_proc_id ? _GEN_3348 : _GEN_2758; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_17 = 2'h3 != last_proc_id ? _GEN_3349 : _GEN_2759; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_18 = 2'h3 != last_proc_id ? _GEN_3350 : _GEN_2760; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_19 = 2'h3 != last_proc_id ? _GEN_3351 : _GEN_2761; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_20 = 2'h3 != last_proc_id ? _GEN_3352 : _GEN_2762; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_21 = 2'h3 != last_proc_id ? _GEN_3353 : _GEN_2763; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_22 = 2'h3 != last_proc_id ? _GEN_3354 : _GEN_2764; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_23 = 2'h3 != last_proc_id ? _GEN_3355 : _GEN_2765; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_24 = 2'h3 != last_proc_id ? _GEN_3356 : _GEN_2766; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_25 = 2'h3 != last_proc_id ? _GEN_3357 : _GEN_2767; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_26 = 2'h3 != last_proc_id ? _GEN_3358 : _GEN_2768; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_27 = 2'h3 != last_proc_id ? _GEN_3359 : _GEN_2769; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_28 = 2'h3 != last_proc_id ? _GEN_3360 : _GEN_2770; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_29 = 2'h3 != last_proc_id ? _GEN_3361 : _GEN_2771; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_30 = 2'h3 != last_proc_id ? _GEN_3362 : _GEN_2772; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_31 = 2'h3 != last_proc_id ? _GEN_3363 : _GEN_2773; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_32 = 2'h3 != last_proc_id ? _GEN_3364 : _GEN_2774; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_33 = 2'h3 != last_proc_id ? _GEN_3365 : _GEN_2775; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_34 = 2'h3 != last_proc_id ? _GEN_3366 : _GEN_2776; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_35 = 2'h3 != last_proc_id ? _GEN_3367 : _GEN_2777; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_36 = 2'h3 != last_proc_id ? _GEN_3368 : _GEN_2778; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_37 = 2'h3 != last_proc_id ? _GEN_3369 : _GEN_2779; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_38 = 2'h3 != last_proc_id ? _GEN_3370 : _GEN_2780; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_39 = 2'h3 != last_proc_id ? _GEN_3371 : _GEN_2781; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_40 = 2'h3 != last_proc_id ? _GEN_3372 : _GEN_2782; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_41 = 2'h3 != last_proc_id ? _GEN_3373 : _GEN_2783; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_42 = 2'h3 != last_proc_id ? _GEN_3374 : _GEN_2784; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_43 = 2'h3 != last_proc_id ? _GEN_3375 : _GEN_2785; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_44 = 2'h3 != last_proc_id ? _GEN_3376 : _GEN_2786; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_45 = 2'h3 != last_proc_id ? _GEN_3377 : _GEN_2787; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_46 = 2'h3 != last_proc_id ? _GEN_3378 : _GEN_2788; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_47 = 2'h3 != last_proc_id ? _GEN_3379 : _GEN_2789; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_48 = 2'h3 != last_proc_id ? _GEN_3380 : _GEN_2790; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_49 = 2'h3 != last_proc_id ? _GEN_3381 : _GEN_2791; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_50 = 2'h3 != last_proc_id ? _GEN_3382 : _GEN_2792; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_51 = 2'h3 != last_proc_id ? _GEN_3383 : _GEN_2793; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_52 = 2'h3 != last_proc_id ? _GEN_3384 : _GEN_2794; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_53 = 2'h3 != last_proc_id ? _GEN_3385 : _GEN_2795; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_54 = 2'h3 != last_proc_id ? _GEN_3386 : _GEN_2796; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_55 = 2'h3 != last_proc_id ? _GEN_3387 : _GEN_2797; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_56 = 2'h3 != last_proc_id ? _GEN_3388 : _GEN_2798; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_57 = 2'h3 != last_proc_id ? _GEN_3389 : _GEN_2799; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_58 = 2'h3 != last_proc_id ? _GEN_3390 : _GEN_2800; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_59 = 2'h3 != last_proc_id ? _GEN_3391 : _GEN_2801; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_60 = 2'h3 != last_proc_id ? _GEN_3392 : _GEN_2802; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_61 = 2'h3 != last_proc_id ? _GEN_3393 : _GEN_2803; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_62 = 2'h3 != last_proc_id ? _GEN_3394 : _GEN_2804; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_63 = 2'h3 != last_proc_id ? _GEN_3395 : _GEN_2805; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_64 = 2'h3 != last_proc_id ? _GEN_3396 : _GEN_2806; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_65 = 2'h3 != last_proc_id ? _GEN_3397 : _GEN_2807; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_66 = 2'h3 != last_proc_id ? _GEN_3398 : _GEN_2808; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_67 = 2'h3 != last_proc_id ? _GEN_3399 : _GEN_2809; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_68 = 2'h3 != last_proc_id ? _GEN_3400 : _GEN_2810; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_69 = 2'h3 != last_proc_id ? _GEN_3401 : _GEN_2811; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_70 = 2'h3 != last_proc_id ? _GEN_3402 : _GEN_2812; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_71 = 2'h3 != last_proc_id ? _GEN_3403 : _GEN_2813; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_72 = 2'h3 != last_proc_id ? _GEN_3404 : _GEN_2814; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_73 = 2'h3 != last_proc_id ? _GEN_3405 : _GEN_2815; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_74 = 2'h3 != last_proc_id ? _GEN_3406 : _GEN_2816; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_75 = 2'h3 != last_proc_id ? _GEN_3407 : _GEN_2817; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_76 = 2'h3 != last_proc_id ? _GEN_3408 : _GEN_2818; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_77 = 2'h3 != last_proc_id ? _GEN_3409 : _GEN_2819; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_78 = 2'h3 != last_proc_id ? _GEN_3410 : _GEN_2820; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_79 = 2'h3 != last_proc_id ? _GEN_3411 : _GEN_2821; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_80 = 2'h3 != last_proc_id ? _GEN_3412 : _GEN_2822; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_81 = 2'h3 != last_proc_id ? _GEN_3413 : _GEN_2823; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_82 = 2'h3 != last_proc_id ? _GEN_3414 : _GEN_2824; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_83 = 2'h3 != last_proc_id ? _GEN_3415 : _GEN_2825; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_84 = 2'h3 != last_proc_id ? _GEN_3416 : _GEN_2826; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_85 = 2'h3 != last_proc_id ? _GEN_3417 : _GEN_2827; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_86 = 2'h3 != last_proc_id ? _GEN_3418 : _GEN_2828; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_87 = 2'h3 != last_proc_id ? _GEN_3419 : _GEN_2829; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_88 = 2'h3 != last_proc_id ? _GEN_3420 : _GEN_2830; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_89 = 2'h3 != last_proc_id ? _GEN_3421 : _GEN_2831; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_90 = 2'h3 != last_proc_id ? _GEN_3422 : _GEN_2832; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_91 = 2'h3 != last_proc_id ? _GEN_3423 : _GEN_2833; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_92 = 2'h3 != last_proc_id ? _GEN_3424 : _GEN_2834; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_93 = 2'h3 != last_proc_id ? _GEN_3425 : _GEN_2835; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_94 = 2'h3 != last_proc_id ? _GEN_3426 : _GEN_2836; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_data_95 = 2'h3 != last_proc_id ? _GEN_3427 : _GEN_2837; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_0 = 2'h3 != last_proc_id ? _GEN_3316 : _GEN_2726; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_1 = 2'h3 != last_proc_id ? _GEN_3317 : _GEN_2727; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_2 = 2'h3 != last_proc_id ? _GEN_3318 : _GEN_2728; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_3 = 2'h3 != last_proc_id ? _GEN_3319 : _GEN_2729; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_4 = 2'h3 != last_proc_id ? _GEN_3320 : _GEN_2730; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_5 = 2'h3 != last_proc_id ? _GEN_3321 : _GEN_2731; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_6 = 2'h3 != last_proc_id ? _GEN_3322 : _GEN_2732; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_7 = 2'h3 != last_proc_id ? _GEN_3323 : _GEN_2733; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_8 = 2'h3 != last_proc_id ? _GEN_3324 : _GEN_2734; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_9 = 2'h3 != last_proc_id ? _GEN_3325 : _GEN_2735; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_10 = 2'h3 != last_proc_id ? _GEN_3326 : _GEN_2736; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_11 = 2'h3 != last_proc_id ? _GEN_3327 : _GEN_2737; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_12 = 2'h3 != last_proc_id ? _GEN_3328 : _GEN_2738; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_13 = 2'h3 != last_proc_id ? _GEN_3329 : _GEN_2739; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_14 = 2'h3 != last_proc_id ? _GEN_3330 : _GEN_2740; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_header_15 = 2'h3 != last_proc_id ? _GEN_3331 : _GEN_2741; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_parse_current_state = 2'h3 != last_proc_id ? _GEN_3315 : _GEN_2725; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_parse_current_offset = 2'h3 != last_proc_id ? _GEN_3314 : _GEN_2724; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_parse_transition_field = 2'h3 != last_proc_id ? _GEN_3313 : _GEN_2723; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_next_processor_id = 2'h3 != last_proc_id ? _GEN_3312 : _GEN_2722; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_next_config_id = 2'h3 != last_proc_id ? _GEN_3311 : _GEN_2721; // @[ipsa.scala 94:65]
  assign proc_1_io_pipe_phv_in_is_valid_processor = 2'h3 != last_proc_id ? _GEN_3310 : _GEN_2720; // @[ipsa.scala 94:65]
  assign proc_1_io_mod_par_mod_en = io_mod_proc_mod_1_par_mod_en; // @[ipsa.scala 57:20]
  assign proc_1_io_mod_par_mod_last_mau_id_mod = io_mod_proc_mod_1_par_mod_last_mau_id_mod; // @[ipsa.scala 57:20]
  assign proc_1_io_mod_par_mod_last_mau_id = io_mod_proc_mod_1_par_mod_last_mau_id; // @[ipsa.scala 57:20]
  assign proc_1_io_mod_par_mod_cs = io_mod_proc_mod_1_par_mod_cs; // @[ipsa.scala 57:20]
  assign proc_1_io_mod_par_mod_module_mod_state_id_mod = io_mod_proc_mod_1_par_mod_module_mod_state_id_mod; // @[ipsa.scala 57:20]
  assign proc_1_io_mod_par_mod_module_mod_state_id = io_mod_proc_mod_1_par_mod_module_mod_state_id; // @[ipsa.scala 57:20]
  assign proc_1_io_mod_par_mod_module_mod_sram_w_cs = io_mod_proc_mod_1_par_mod_module_mod_sram_w_cs; // @[ipsa.scala 57:20]
  assign proc_1_io_mod_par_mod_module_mod_sram_w_addr = io_mod_proc_mod_1_par_mod_module_mod_sram_w_addr; // @[ipsa.scala 57:20]
  assign proc_1_io_mod_par_mod_module_mod_sram_w_data = io_mod_proc_mod_1_par_mod_module_mod_sram_w_data; // @[ipsa.scala 57:20]
  assign proc_1_io_mod_mat_mod_en = io_mod_proc_mod_1_mat_mod_en; // @[ipsa.scala 57:20]
  assign proc_1_io_mod_mat_mod_config_id = io_mod_proc_mod_1_mat_mod_config_id; // @[ipsa.scala 57:20]
  assign proc_1_io_mod_mat_mod_key_mod_header_id = io_mod_proc_mod_1_mat_mod_key_mod_header_id; // @[ipsa.scala 57:20]
  assign proc_1_io_mod_mat_mod_key_mod_internal_offset = io_mod_proc_mod_1_mat_mod_key_mod_internal_offset; // @[ipsa.scala 57:20]
  assign proc_1_io_mod_mat_mod_key_mod_key_length = io_mod_proc_mod_1_mat_mod_key_mod_key_length; // @[ipsa.scala 57:20]
  assign proc_1_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_1_mat_mod_table_mod_table_width; // @[ipsa.scala 57:20]
  assign proc_1_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_1_mat_mod_table_mod_table_depth; // @[ipsa.scala 57:20]
  assign proc_1_io_mod_act_mod_en = io_mod_proc_mod_1_act_mod_en; // @[ipsa.scala 57:20]
  assign proc_1_io_mod_act_mod_addr = io_mod_proc_mod_1_act_mod_addr; // @[ipsa.scala 57:20]
  assign proc_1_io_mod_act_mod_data_0 = io_mod_proc_mod_1_act_mod_data_0; // @[ipsa.scala 57:20]
  assign proc_1_io_mod_act_mod_data_1 = io_mod_proc_mod_1_act_mod_data_1; // @[ipsa.scala 57:20]
  assign proc_1_io_mem_cluster_0_data = sram_cluster_0_io_r_1_cluster_0_data; // @[ipsa.scala 70:37]
  assign proc_1_io_mem_cluster_1_data = sram_cluster_0_io_r_1_cluster_1_data; // @[ipsa.scala 70:37]
  assign proc_1_io_mem_cluster_2_data = sram_cluster_0_io_r_1_cluster_2_data; // @[ipsa.scala 70:37]
  assign proc_1_io_mem_cluster_3_data = sram_cluster_0_io_r_1_cluster_3_data; // @[ipsa.scala 70:37]
  assign proc_1_io_mem_cluster_4_data = sram_cluster_0_io_r_1_cluster_4_data; // @[ipsa.scala 70:37]
  assign proc_1_io_mem_cluster_5_data = sram_cluster_0_io_r_1_cluster_5_data; // @[ipsa.scala 70:37]
  assign proc_1_io_mem_cluster_6_data = sram_cluster_0_io_r_1_cluster_6_data; // @[ipsa.scala 70:37]
  assign proc_1_io_mem_cluster_7_data = sram_cluster_0_io_r_1_cluster_7_data; // @[ipsa.scala 70:37]
  assign proc_2_clock = clock;
  assign proc_2_io_pipe_phv_in_data_0 = 2'h3 != last_proc_id ? _GEN_3450 : _GEN_2860; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_1 = 2'h3 != last_proc_id ? _GEN_3451 : _GEN_2861; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_2 = 2'h3 != last_proc_id ? _GEN_3452 : _GEN_2862; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_3 = 2'h3 != last_proc_id ? _GEN_3453 : _GEN_2863; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_4 = 2'h3 != last_proc_id ? _GEN_3454 : _GEN_2864; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_5 = 2'h3 != last_proc_id ? _GEN_3455 : _GEN_2865; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_6 = 2'h3 != last_proc_id ? _GEN_3456 : _GEN_2866; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_7 = 2'h3 != last_proc_id ? _GEN_3457 : _GEN_2867; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_8 = 2'h3 != last_proc_id ? _GEN_3458 : _GEN_2868; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_9 = 2'h3 != last_proc_id ? _GEN_3459 : _GEN_2869; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_10 = 2'h3 != last_proc_id ? _GEN_3460 : _GEN_2870; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_11 = 2'h3 != last_proc_id ? _GEN_3461 : _GEN_2871; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_12 = 2'h3 != last_proc_id ? _GEN_3462 : _GEN_2872; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_13 = 2'h3 != last_proc_id ? _GEN_3463 : _GEN_2873; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_14 = 2'h3 != last_proc_id ? _GEN_3464 : _GEN_2874; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_15 = 2'h3 != last_proc_id ? _GEN_3465 : _GEN_2875; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_16 = 2'h3 != last_proc_id ? _GEN_3466 : _GEN_2876; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_17 = 2'h3 != last_proc_id ? _GEN_3467 : _GEN_2877; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_18 = 2'h3 != last_proc_id ? _GEN_3468 : _GEN_2878; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_19 = 2'h3 != last_proc_id ? _GEN_3469 : _GEN_2879; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_20 = 2'h3 != last_proc_id ? _GEN_3470 : _GEN_2880; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_21 = 2'h3 != last_proc_id ? _GEN_3471 : _GEN_2881; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_22 = 2'h3 != last_proc_id ? _GEN_3472 : _GEN_2882; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_23 = 2'h3 != last_proc_id ? _GEN_3473 : _GEN_2883; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_24 = 2'h3 != last_proc_id ? _GEN_3474 : _GEN_2884; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_25 = 2'h3 != last_proc_id ? _GEN_3475 : _GEN_2885; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_26 = 2'h3 != last_proc_id ? _GEN_3476 : _GEN_2886; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_27 = 2'h3 != last_proc_id ? _GEN_3477 : _GEN_2887; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_28 = 2'h3 != last_proc_id ? _GEN_3478 : _GEN_2888; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_29 = 2'h3 != last_proc_id ? _GEN_3479 : _GEN_2889; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_30 = 2'h3 != last_proc_id ? _GEN_3480 : _GEN_2890; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_31 = 2'h3 != last_proc_id ? _GEN_3481 : _GEN_2891; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_32 = 2'h3 != last_proc_id ? _GEN_3482 : _GEN_2892; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_33 = 2'h3 != last_proc_id ? _GEN_3483 : _GEN_2893; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_34 = 2'h3 != last_proc_id ? _GEN_3484 : _GEN_2894; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_35 = 2'h3 != last_proc_id ? _GEN_3485 : _GEN_2895; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_36 = 2'h3 != last_proc_id ? _GEN_3486 : _GEN_2896; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_37 = 2'h3 != last_proc_id ? _GEN_3487 : _GEN_2897; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_38 = 2'h3 != last_proc_id ? _GEN_3488 : _GEN_2898; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_39 = 2'h3 != last_proc_id ? _GEN_3489 : _GEN_2899; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_40 = 2'h3 != last_proc_id ? _GEN_3490 : _GEN_2900; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_41 = 2'h3 != last_proc_id ? _GEN_3491 : _GEN_2901; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_42 = 2'h3 != last_proc_id ? _GEN_3492 : _GEN_2902; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_43 = 2'h3 != last_proc_id ? _GEN_3493 : _GEN_2903; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_44 = 2'h3 != last_proc_id ? _GEN_3494 : _GEN_2904; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_45 = 2'h3 != last_proc_id ? _GEN_3495 : _GEN_2905; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_46 = 2'h3 != last_proc_id ? _GEN_3496 : _GEN_2906; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_47 = 2'h3 != last_proc_id ? _GEN_3497 : _GEN_2907; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_48 = 2'h3 != last_proc_id ? _GEN_3498 : _GEN_2908; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_49 = 2'h3 != last_proc_id ? _GEN_3499 : _GEN_2909; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_50 = 2'h3 != last_proc_id ? _GEN_3500 : _GEN_2910; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_51 = 2'h3 != last_proc_id ? _GEN_3501 : _GEN_2911; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_52 = 2'h3 != last_proc_id ? _GEN_3502 : _GEN_2912; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_53 = 2'h3 != last_proc_id ? _GEN_3503 : _GEN_2913; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_54 = 2'h3 != last_proc_id ? _GEN_3504 : _GEN_2914; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_55 = 2'h3 != last_proc_id ? _GEN_3505 : _GEN_2915; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_56 = 2'h3 != last_proc_id ? _GEN_3506 : _GEN_2916; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_57 = 2'h3 != last_proc_id ? _GEN_3507 : _GEN_2917; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_58 = 2'h3 != last_proc_id ? _GEN_3508 : _GEN_2918; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_59 = 2'h3 != last_proc_id ? _GEN_3509 : _GEN_2919; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_60 = 2'h3 != last_proc_id ? _GEN_3510 : _GEN_2920; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_61 = 2'h3 != last_proc_id ? _GEN_3511 : _GEN_2921; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_62 = 2'h3 != last_proc_id ? _GEN_3512 : _GEN_2922; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_63 = 2'h3 != last_proc_id ? _GEN_3513 : _GEN_2923; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_64 = 2'h3 != last_proc_id ? _GEN_3514 : _GEN_2924; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_65 = 2'h3 != last_proc_id ? _GEN_3515 : _GEN_2925; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_66 = 2'h3 != last_proc_id ? _GEN_3516 : _GEN_2926; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_67 = 2'h3 != last_proc_id ? _GEN_3517 : _GEN_2927; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_68 = 2'h3 != last_proc_id ? _GEN_3518 : _GEN_2928; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_69 = 2'h3 != last_proc_id ? _GEN_3519 : _GEN_2929; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_70 = 2'h3 != last_proc_id ? _GEN_3520 : _GEN_2930; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_71 = 2'h3 != last_proc_id ? _GEN_3521 : _GEN_2931; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_72 = 2'h3 != last_proc_id ? _GEN_3522 : _GEN_2932; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_73 = 2'h3 != last_proc_id ? _GEN_3523 : _GEN_2933; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_74 = 2'h3 != last_proc_id ? _GEN_3524 : _GEN_2934; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_75 = 2'h3 != last_proc_id ? _GEN_3525 : _GEN_2935; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_76 = 2'h3 != last_proc_id ? _GEN_3526 : _GEN_2936; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_77 = 2'h3 != last_proc_id ? _GEN_3527 : _GEN_2937; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_78 = 2'h3 != last_proc_id ? _GEN_3528 : _GEN_2938; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_79 = 2'h3 != last_proc_id ? _GEN_3529 : _GEN_2939; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_80 = 2'h3 != last_proc_id ? _GEN_3530 : _GEN_2940; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_81 = 2'h3 != last_proc_id ? _GEN_3531 : _GEN_2941; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_82 = 2'h3 != last_proc_id ? _GEN_3532 : _GEN_2942; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_83 = 2'h3 != last_proc_id ? _GEN_3533 : _GEN_2943; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_84 = 2'h3 != last_proc_id ? _GEN_3534 : _GEN_2944; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_85 = 2'h3 != last_proc_id ? _GEN_3535 : _GEN_2945; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_86 = 2'h3 != last_proc_id ? _GEN_3536 : _GEN_2946; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_87 = 2'h3 != last_proc_id ? _GEN_3537 : _GEN_2947; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_88 = 2'h3 != last_proc_id ? _GEN_3538 : _GEN_2948; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_89 = 2'h3 != last_proc_id ? _GEN_3539 : _GEN_2949; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_90 = 2'h3 != last_proc_id ? _GEN_3540 : _GEN_2950; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_91 = 2'h3 != last_proc_id ? _GEN_3541 : _GEN_2951; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_92 = 2'h3 != last_proc_id ? _GEN_3542 : _GEN_2952; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_93 = 2'h3 != last_proc_id ? _GEN_3543 : _GEN_2953; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_94 = 2'h3 != last_proc_id ? _GEN_3544 : _GEN_2954; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_data_95 = 2'h3 != last_proc_id ? _GEN_3545 : _GEN_2955; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_0 = 2'h3 != last_proc_id ? _GEN_3434 : _GEN_2844; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_1 = 2'h3 != last_proc_id ? _GEN_3435 : _GEN_2845; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_2 = 2'h3 != last_proc_id ? _GEN_3436 : _GEN_2846; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_3 = 2'h3 != last_proc_id ? _GEN_3437 : _GEN_2847; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_4 = 2'h3 != last_proc_id ? _GEN_3438 : _GEN_2848; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_5 = 2'h3 != last_proc_id ? _GEN_3439 : _GEN_2849; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_6 = 2'h3 != last_proc_id ? _GEN_3440 : _GEN_2850; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_7 = 2'h3 != last_proc_id ? _GEN_3441 : _GEN_2851; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_8 = 2'h3 != last_proc_id ? _GEN_3442 : _GEN_2852; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_9 = 2'h3 != last_proc_id ? _GEN_3443 : _GEN_2853; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_10 = 2'h3 != last_proc_id ? _GEN_3444 : _GEN_2854; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_11 = 2'h3 != last_proc_id ? _GEN_3445 : _GEN_2855; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_12 = 2'h3 != last_proc_id ? _GEN_3446 : _GEN_2856; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_13 = 2'h3 != last_proc_id ? _GEN_3447 : _GEN_2857; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_14 = 2'h3 != last_proc_id ? _GEN_3448 : _GEN_2858; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_header_15 = 2'h3 != last_proc_id ? _GEN_3449 : _GEN_2859; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_parse_current_state = 2'h3 != last_proc_id ? _GEN_3433 : _GEN_2843; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_parse_current_offset = 2'h3 != last_proc_id ? _GEN_3432 : _GEN_2842; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_parse_transition_field = 2'h3 != last_proc_id ? _GEN_3431 : _GEN_2841; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_next_processor_id = 2'h3 != last_proc_id ? _GEN_3430 : _GEN_2840; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_next_config_id = 2'h3 != last_proc_id ? _GEN_3429 : _GEN_2839; // @[ipsa.scala 94:65]
  assign proc_2_io_pipe_phv_in_is_valid_processor = 2'h3 != last_proc_id ? _GEN_3428 : _GEN_2838; // @[ipsa.scala 94:65]
  assign proc_2_io_mod_par_mod_en = io_mod_proc_mod_2_par_mod_en; // @[ipsa.scala 57:20]
  assign proc_2_io_mod_par_mod_last_mau_id_mod = io_mod_proc_mod_2_par_mod_last_mau_id_mod; // @[ipsa.scala 57:20]
  assign proc_2_io_mod_par_mod_last_mau_id = io_mod_proc_mod_2_par_mod_last_mau_id; // @[ipsa.scala 57:20]
  assign proc_2_io_mod_par_mod_cs = io_mod_proc_mod_2_par_mod_cs; // @[ipsa.scala 57:20]
  assign proc_2_io_mod_par_mod_module_mod_state_id_mod = io_mod_proc_mod_2_par_mod_module_mod_state_id_mod; // @[ipsa.scala 57:20]
  assign proc_2_io_mod_par_mod_module_mod_state_id = io_mod_proc_mod_2_par_mod_module_mod_state_id; // @[ipsa.scala 57:20]
  assign proc_2_io_mod_par_mod_module_mod_sram_w_cs = io_mod_proc_mod_2_par_mod_module_mod_sram_w_cs; // @[ipsa.scala 57:20]
  assign proc_2_io_mod_par_mod_module_mod_sram_w_addr = io_mod_proc_mod_2_par_mod_module_mod_sram_w_addr; // @[ipsa.scala 57:20]
  assign proc_2_io_mod_par_mod_module_mod_sram_w_data = io_mod_proc_mod_2_par_mod_module_mod_sram_w_data; // @[ipsa.scala 57:20]
  assign proc_2_io_mod_mat_mod_en = io_mod_proc_mod_2_mat_mod_en; // @[ipsa.scala 57:20]
  assign proc_2_io_mod_mat_mod_config_id = io_mod_proc_mod_2_mat_mod_config_id; // @[ipsa.scala 57:20]
  assign proc_2_io_mod_mat_mod_key_mod_header_id = io_mod_proc_mod_2_mat_mod_key_mod_header_id; // @[ipsa.scala 57:20]
  assign proc_2_io_mod_mat_mod_key_mod_internal_offset = io_mod_proc_mod_2_mat_mod_key_mod_internal_offset; // @[ipsa.scala 57:20]
  assign proc_2_io_mod_mat_mod_key_mod_key_length = io_mod_proc_mod_2_mat_mod_key_mod_key_length; // @[ipsa.scala 57:20]
  assign proc_2_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_2_mat_mod_table_mod_table_width; // @[ipsa.scala 57:20]
  assign proc_2_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_2_mat_mod_table_mod_table_depth; // @[ipsa.scala 57:20]
  assign proc_2_io_mod_act_mod_en = io_mod_proc_mod_2_act_mod_en; // @[ipsa.scala 57:20]
  assign proc_2_io_mod_act_mod_addr = io_mod_proc_mod_2_act_mod_addr; // @[ipsa.scala 57:20]
  assign proc_2_io_mod_act_mod_data_0 = io_mod_proc_mod_2_act_mod_data_0; // @[ipsa.scala 57:20]
  assign proc_2_io_mod_act_mod_data_1 = io_mod_proc_mod_2_act_mod_data_1; // @[ipsa.scala 57:20]
  assign proc_2_io_mem_cluster_0_data = sram_cluster_0_io_r_2_cluster_0_data; // @[ipsa.scala 70:37]
  assign proc_2_io_mem_cluster_1_data = sram_cluster_0_io_r_2_cluster_1_data; // @[ipsa.scala 70:37]
  assign proc_2_io_mem_cluster_2_data = sram_cluster_0_io_r_2_cluster_2_data; // @[ipsa.scala 70:37]
  assign proc_2_io_mem_cluster_3_data = sram_cluster_0_io_r_2_cluster_3_data; // @[ipsa.scala 70:37]
  assign proc_2_io_mem_cluster_4_data = sram_cluster_0_io_r_2_cluster_4_data; // @[ipsa.scala 70:37]
  assign proc_2_io_mem_cluster_5_data = sram_cluster_0_io_r_2_cluster_5_data; // @[ipsa.scala 70:37]
  assign proc_2_io_mem_cluster_6_data = sram_cluster_0_io_r_2_cluster_6_data; // @[ipsa.scala 70:37]
  assign proc_2_io_mem_cluster_7_data = sram_cluster_0_io_r_2_cluster_7_data; // @[ipsa.scala 70:37]
  assign proc_3_clock = clock;
  assign proc_3_io_pipe_phv_in_data_0 = 2'h3 != last_proc_id ? _GEN_3568 : _GEN_2978; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_1 = 2'h3 != last_proc_id ? _GEN_3569 : _GEN_2979; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_2 = 2'h3 != last_proc_id ? _GEN_3570 : _GEN_2980; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_3 = 2'h3 != last_proc_id ? _GEN_3571 : _GEN_2981; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_4 = 2'h3 != last_proc_id ? _GEN_3572 : _GEN_2982; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_5 = 2'h3 != last_proc_id ? _GEN_3573 : _GEN_2983; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_6 = 2'h3 != last_proc_id ? _GEN_3574 : _GEN_2984; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_7 = 2'h3 != last_proc_id ? _GEN_3575 : _GEN_2985; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_8 = 2'h3 != last_proc_id ? _GEN_3576 : _GEN_2986; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_9 = 2'h3 != last_proc_id ? _GEN_3577 : _GEN_2987; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_10 = 2'h3 != last_proc_id ? _GEN_3578 : _GEN_2988; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_11 = 2'h3 != last_proc_id ? _GEN_3579 : _GEN_2989; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_12 = 2'h3 != last_proc_id ? _GEN_3580 : _GEN_2990; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_13 = 2'h3 != last_proc_id ? _GEN_3581 : _GEN_2991; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_14 = 2'h3 != last_proc_id ? _GEN_3582 : _GEN_2992; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_15 = 2'h3 != last_proc_id ? _GEN_3583 : _GEN_2993; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_16 = 2'h3 != last_proc_id ? _GEN_3584 : _GEN_2994; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_17 = 2'h3 != last_proc_id ? _GEN_3585 : _GEN_2995; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_18 = 2'h3 != last_proc_id ? _GEN_3586 : _GEN_2996; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_19 = 2'h3 != last_proc_id ? _GEN_3587 : _GEN_2997; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_20 = 2'h3 != last_proc_id ? _GEN_3588 : _GEN_2998; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_21 = 2'h3 != last_proc_id ? _GEN_3589 : _GEN_2999; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_22 = 2'h3 != last_proc_id ? _GEN_3590 : _GEN_3000; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_23 = 2'h3 != last_proc_id ? _GEN_3591 : _GEN_3001; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_24 = 2'h3 != last_proc_id ? _GEN_3592 : _GEN_3002; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_25 = 2'h3 != last_proc_id ? _GEN_3593 : _GEN_3003; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_26 = 2'h3 != last_proc_id ? _GEN_3594 : _GEN_3004; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_27 = 2'h3 != last_proc_id ? _GEN_3595 : _GEN_3005; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_28 = 2'h3 != last_proc_id ? _GEN_3596 : _GEN_3006; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_29 = 2'h3 != last_proc_id ? _GEN_3597 : _GEN_3007; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_30 = 2'h3 != last_proc_id ? _GEN_3598 : _GEN_3008; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_31 = 2'h3 != last_proc_id ? _GEN_3599 : _GEN_3009; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_32 = 2'h3 != last_proc_id ? _GEN_3600 : _GEN_3010; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_33 = 2'h3 != last_proc_id ? _GEN_3601 : _GEN_3011; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_34 = 2'h3 != last_proc_id ? _GEN_3602 : _GEN_3012; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_35 = 2'h3 != last_proc_id ? _GEN_3603 : _GEN_3013; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_36 = 2'h3 != last_proc_id ? _GEN_3604 : _GEN_3014; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_37 = 2'h3 != last_proc_id ? _GEN_3605 : _GEN_3015; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_38 = 2'h3 != last_proc_id ? _GEN_3606 : _GEN_3016; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_39 = 2'h3 != last_proc_id ? _GEN_3607 : _GEN_3017; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_40 = 2'h3 != last_proc_id ? _GEN_3608 : _GEN_3018; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_41 = 2'h3 != last_proc_id ? _GEN_3609 : _GEN_3019; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_42 = 2'h3 != last_proc_id ? _GEN_3610 : _GEN_3020; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_43 = 2'h3 != last_proc_id ? _GEN_3611 : _GEN_3021; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_44 = 2'h3 != last_proc_id ? _GEN_3612 : _GEN_3022; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_45 = 2'h3 != last_proc_id ? _GEN_3613 : _GEN_3023; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_46 = 2'h3 != last_proc_id ? _GEN_3614 : _GEN_3024; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_47 = 2'h3 != last_proc_id ? _GEN_3615 : _GEN_3025; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_48 = 2'h3 != last_proc_id ? _GEN_3616 : _GEN_3026; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_49 = 2'h3 != last_proc_id ? _GEN_3617 : _GEN_3027; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_50 = 2'h3 != last_proc_id ? _GEN_3618 : _GEN_3028; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_51 = 2'h3 != last_proc_id ? _GEN_3619 : _GEN_3029; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_52 = 2'h3 != last_proc_id ? _GEN_3620 : _GEN_3030; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_53 = 2'h3 != last_proc_id ? _GEN_3621 : _GEN_3031; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_54 = 2'h3 != last_proc_id ? _GEN_3622 : _GEN_3032; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_55 = 2'h3 != last_proc_id ? _GEN_3623 : _GEN_3033; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_56 = 2'h3 != last_proc_id ? _GEN_3624 : _GEN_3034; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_57 = 2'h3 != last_proc_id ? _GEN_3625 : _GEN_3035; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_58 = 2'h3 != last_proc_id ? _GEN_3626 : _GEN_3036; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_59 = 2'h3 != last_proc_id ? _GEN_3627 : _GEN_3037; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_60 = 2'h3 != last_proc_id ? _GEN_3628 : _GEN_3038; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_61 = 2'h3 != last_proc_id ? _GEN_3629 : _GEN_3039; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_62 = 2'h3 != last_proc_id ? _GEN_3630 : _GEN_3040; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_63 = 2'h3 != last_proc_id ? _GEN_3631 : _GEN_3041; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_64 = 2'h3 != last_proc_id ? _GEN_3632 : _GEN_3042; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_65 = 2'h3 != last_proc_id ? _GEN_3633 : _GEN_3043; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_66 = 2'h3 != last_proc_id ? _GEN_3634 : _GEN_3044; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_67 = 2'h3 != last_proc_id ? _GEN_3635 : _GEN_3045; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_68 = 2'h3 != last_proc_id ? _GEN_3636 : _GEN_3046; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_69 = 2'h3 != last_proc_id ? _GEN_3637 : _GEN_3047; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_70 = 2'h3 != last_proc_id ? _GEN_3638 : _GEN_3048; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_71 = 2'h3 != last_proc_id ? _GEN_3639 : _GEN_3049; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_72 = 2'h3 != last_proc_id ? _GEN_3640 : _GEN_3050; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_73 = 2'h3 != last_proc_id ? _GEN_3641 : _GEN_3051; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_74 = 2'h3 != last_proc_id ? _GEN_3642 : _GEN_3052; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_75 = 2'h3 != last_proc_id ? _GEN_3643 : _GEN_3053; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_76 = 2'h3 != last_proc_id ? _GEN_3644 : _GEN_3054; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_77 = 2'h3 != last_proc_id ? _GEN_3645 : _GEN_3055; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_78 = 2'h3 != last_proc_id ? _GEN_3646 : _GEN_3056; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_79 = 2'h3 != last_proc_id ? _GEN_3647 : _GEN_3057; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_80 = 2'h3 != last_proc_id ? _GEN_3648 : _GEN_3058; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_81 = 2'h3 != last_proc_id ? _GEN_3649 : _GEN_3059; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_82 = 2'h3 != last_proc_id ? _GEN_3650 : _GEN_3060; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_83 = 2'h3 != last_proc_id ? _GEN_3651 : _GEN_3061; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_84 = 2'h3 != last_proc_id ? _GEN_3652 : _GEN_3062; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_85 = 2'h3 != last_proc_id ? _GEN_3653 : _GEN_3063; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_86 = 2'h3 != last_proc_id ? _GEN_3654 : _GEN_3064; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_87 = 2'h3 != last_proc_id ? _GEN_3655 : _GEN_3065; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_88 = 2'h3 != last_proc_id ? _GEN_3656 : _GEN_3066; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_89 = 2'h3 != last_proc_id ? _GEN_3657 : _GEN_3067; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_90 = 2'h3 != last_proc_id ? _GEN_3658 : _GEN_3068; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_91 = 2'h3 != last_proc_id ? _GEN_3659 : _GEN_3069; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_92 = 2'h3 != last_proc_id ? _GEN_3660 : _GEN_3070; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_93 = 2'h3 != last_proc_id ? _GEN_3661 : _GEN_3071; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_94 = 2'h3 != last_proc_id ? _GEN_3662 : _GEN_3072; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_data_95 = 2'h3 != last_proc_id ? _GEN_3663 : _GEN_3073; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_0 = 2'h3 != last_proc_id ? _GEN_3552 : _GEN_2962; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_1 = 2'h3 != last_proc_id ? _GEN_3553 : _GEN_2963; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_2 = 2'h3 != last_proc_id ? _GEN_3554 : _GEN_2964; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_3 = 2'h3 != last_proc_id ? _GEN_3555 : _GEN_2965; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_4 = 2'h3 != last_proc_id ? _GEN_3556 : _GEN_2966; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_5 = 2'h3 != last_proc_id ? _GEN_3557 : _GEN_2967; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_6 = 2'h3 != last_proc_id ? _GEN_3558 : _GEN_2968; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_7 = 2'h3 != last_proc_id ? _GEN_3559 : _GEN_2969; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_8 = 2'h3 != last_proc_id ? _GEN_3560 : _GEN_2970; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_9 = 2'h3 != last_proc_id ? _GEN_3561 : _GEN_2971; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_10 = 2'h3 != last_proc_id ? _GEN_3562 : _GEN_2972; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_11 = 2'h3 != last_proc_id ? _GEN_3563 : _GEN_2973; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_12 = 2'h3 != last_proc_id ? _GEN_3564 : _GEN_2974; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_13 = 2'h3 != last_proc_id ? _GEN_3565 : _GEN_2975; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_14 = 2'h3 != last_proc_id ? _GEN_3566 : _GEN_2976; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_header_15 = 2'h3 != last_proc_id ? _GEN_3567 : _GEN_2977; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_parse_current_state = 2'h3 != last_proc_id ? _GEN_3551 : _GEN_2961; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_parse_current_offset = 2'h3 != last_proc_id ? _GEN_3550 : _GEN_2960; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_parse_transition_field = 2'h3 != last_proc_id ? _GEN_3549 : _GEN_2959; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_next_processor_id = 2'h3 != last_proc_id ? _GEN_3548 : _GEN_2958; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_next_config_id = 2'h3 != last_proc_id ? _GEN_3547 : _GEN_2957; // @[ipsa.scala 94:65]
  assign proc_3_io_pipe_phv_in_is_valid_processor = 2'h3 != last_proc_id ? _GEN_3546 : _GEN_2956; // @[ipsa.scala 94:65]
  assign proc_3_io_mod_par_mod_en = io_mod_proc_mod_3_par_mod_en; // @[ipsa.scala 57:20]
  assign proc_3_io_mod_par_mod_last_mau_id_mod = io_mod_proc_mod_3_par_mod_last_mau_id_mod; // @[ipsa.scala 57:20]
  assign proc_3_io_mod_par_mod_last_mau_id = io_mod_proc_mod_3_par_mod_last_mau_id; // @[ipsa.scala 57:20]
  assign proc_3_io_mod_par_mod_cs = io_mod_proc_mod_3_par_mod_cs; // @[ipsa.scala 57:20]
  assign proc_3_io_mod_par_mod_module_mod_state_id_mod = io_mod_proc_mod_3_par_mod_module_mod_state_id_mod; // @[ipsa.scala 57:20]
  assign proc_3_io_mod_par_mod_module_mod_state_id = io_mod_proc_mod_3_par_mod_module_mod_state_id; // @[ipsa.scala 57:20]
  assign proc_3_io_mod_par_mod_module_mod_sram_w_cs = io_mod_proc_mod_3_par_mod_module_mod_sram_w_cs; // @[ipsa.scala 57:20]
  assign proc_3_io_mod_par_mod_module_mod_sram_w_addr = io_mod_proc_mod_3_par_mod_module_mod_sram_w_addr; // @[ipsa.scala 57:20]
  assign proc_3_io_mod_par_mod_module_mod_sram_w_data = io_mod_proc_mod_3_par_mod_module_mod_sram_w_data; // @[ipsa.scala 57:20]
  assign proc_3_io_mod_mat_mod_en = io_mod_proc_mod_3_mat_mod_en; // @[ipsa.scala 57:20]
  assign proc_3_io_mod_mat_mod_config_id = io_mod_proc_mod_3_mat_mod_config_id; // @[ipsa.scala 57:20]
  assign proc_3_io_mod_mat_mod_key_mod_header_id = io_mod_proc_mod_3_mat_mod_key_mod_header_id; // @[ipsa.scala 57:20]
  assign proc_3_io_mod_mat_mod_key_mod_internal_offset = io_mod_proc_mod_3_mat_mod_key_mod_internal_offset; // @[ipsa.scala 57:20]
  assign proc_3_io_mod_mat_mod_key_mod_key_length = io_mod_proc_mod_3_mat_mod_key_mod_key_length; // @[ipsa.scala 57:20]
  assign proc_3_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_3_mat_mod_table_mod_table_width; // @[ipsa.scala 57:20]
  assign proc_3_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_3_mat_mod_table_mod_table_depth; // @[ipsa.scala 57:20]
  assign proc_3_io_mod_act_mod_en = io_mod_proc_mod_3_act_mod_en; // @[ipsa.scala 57:20]
  assign proc_3_io_mod_act_mod_addr = io_mod_proc_mod_3_act_mod_addr; // @[ipsa.scala 57:20]
  assign proc_3_io_mod_act_mod_data_0 = io_mod_proc_mod_3_act_mod_data_0; // @[ipsa.scala 57:20]
  assign proc_3_io_mod_act_mod_data_1 = io_mod_proc_mod_3_act_mod_data_1; // @[ipsa.scala 57:20]
  assign proc_3_io_mem_cluster_0_data = sram_cluster_0_io_r_3_cluster_0_data; // @[ipsa.scala 70:37]
  assign proc_3_io_mem_cluster_1_data = sram_cluster_0_io_r_3_cluster_1_data; // @[ipsa.scala 70:37]
  assign proc_3_io_mem_cluster_2_data = sram_cluster_0_io_r_3_cluster_2_data; // @[ipsa.scala 70:37]
  assign proc_3_io_mem_cluster_3_data = sram_cluster_0_io_r_3_cluster_3_data; // @[ipsa.scala 70:37]
  assign proc_3_io_mem_cluster_4_data = sram_cluster_0_io_r_3_cluster_4_data; // @[ipsa.scala 70:37]
  assign proc_3_io_mem_cluster_5_data = sram_cluster_0_io_r_3_cluster_5_data; // @[ipsa.scala 70:37]
  assign proc_3_io_mem_cluster_6_data = sram_cluster_0_io_r_3_cluster_6_data; // @[ipsa.scala 70:37]
  assign proc_3_io_mem_cluster_7_data = sram_cluster_0_io_r_3_cluster_7_data; // @[ipsa.scala 70:37]
  assign sram_cluster_0_clock = clock;
  assign sram_cluster_0_io_w_wcs = io_w_0_wcs; // @[ipsa.scala 63:18]
  assign sram_cluster_0_io_w_w_en = io_w_0_w_en; // @[ipsa.scala 63:18]
  assign sram_cluster_0_io_w_w_addr = io_w_0_w_addr; // @[ipsa.scala 63:18]
  assign sram_cluster_0_io_w_w_data = io_w_0_w_data; // @[ipsa.scala 63:18]
  assign sram_cluster_0_io_r_0_cluster_0_en = proc_0_io_mem_cluster_0_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_0_cluster_0_addr = proc_0_io_mem_cluster_0_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_0_cluster_1_en = proc_0_io_mem_cluster_1_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_0_cluster_1_addr = proc_0_io_mem_cluster_1_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_0_cluster_2_en = proc_0_io_mem_cluster_2_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_0_cluster_2_addr = proc_0_io_mem_cluster_2_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_0_cluster_3_en = proc_0_io_mem_cluster_3_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_0_cluster_3_addr = proc_0_io_mem_cluster_3_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_0_cluster_4_en = proc_0_io_mem_cluster_4_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_0_cluster_4_addr = proc_0_io_mem_cluster_4_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_0_cluster_5_en = proc_0_io_mem_cluster_5_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_0_cluster_5_addr = proc_0_io_mem_cluster_5_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_0_cluster_6_en = proc_0_io_mem_cluster_6_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_0_cluster_6_addr = proc_0_io_mem_cluster_6_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_0_cluster_7_en = proc_0_io_mem_cluster_7_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_0_cluster_7_addr = proc_0_io_mem_cluster_7_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_1_cluster_0_en = proc_1_io_mem_cluster_0_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_1_cluster_0_addr = proc_1_io_mem_cluster_0_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_1_cluster_1_en = proc_1_io_mem_cluster_1_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_1_cluster_1_addr = proc_1_io_mem_cluster_1_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_1_cluster_2_en = proc_1_io_mem_cluster_2_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_1_cluster_2_addr = proc_1_io_mem_cluster_2_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_1_cluster_3_en = proc_1_io_mem_cluster_3_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_1_cluster_3_addr = proc_1_io_mem_cluster_3_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_1_cluster_4_en = proc_1_io_mem_cluster_4_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_1_cluster_4_addr = proc_1_io_mem_cluster_4_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_1_cluster_5_en = proc_1_io_mem_cluster_5_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_1_cluster_5_addr = proc_1_io_mem_cluster_5_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_1_cluster_6_en = proc_1_io_mem_cluster_6_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_1_cluster_6_addr = proc_1_io_mem_cluster_6_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_1_cluster_7_en = proc_1_io_mem_cluster_7_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_1_cluster_7_addr = proc_1_io_mem_cluster_7_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_2_cluster_0_en = proc_2_io_mem_cluster_0_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_2_cluster_0_addr = proc_2_io_mem_cluster_0_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_2_cluster_1_en = proc_2_io_mem_cluster_1_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_2_cluster_1_addr = proc_2_io_mem_cluster_1_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_2_cluster_2_en = proc_2_io_mem_cluster_2_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_2_cluster_2_addr = proc_2_io_mem_cluster_2_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_2_cluster_3_en = proc_2_io_mem_cluster_3_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_2_cluster_3_addr = proc_2_io_mem_cluster_3_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_2_cluster_4_en = proc_2_io_mem_cluster_4_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_2_cluster_4_addr = proc_2_io_mem_cluster_4_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_2_cluster_5_en = proc_2_io_mem_cluster_5_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_2_cluster_5_addr = proc_2_io_mem_cluster_5_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_2_cluster_6_en = proc_2_io_mem_cluster_6_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_2_cluster_6_addr = proc_2_io_mem_cluster_6_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_2_cluster_7_en = proc_2_io_mem_cluster_7_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_2_cluster_7_addr = proc_2_io_mem_cluster_7_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_3_cluster_0_en = proc_3_io_mem_cluster_0_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_3_cluster_0_addr = proc_3_io_mem_cluster_0_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_3_cluster_1_en = proc_3_io_mem_cluster_1_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_3_cluster_1_addr = proc_3_io_mem_cluster_1_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_3_cluster_2_en = proc_3_io_mem_cluster_2_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_3_cluster_2_addr = proc_3_io_mem_cluster_2_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_3_cluster_3_en = proc_3_io_mem_cluster_3_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_3_cluster_3_addr = proc_3_io_mem_cluster_3_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_3_cluster_4_en = proc_3_io_mem_cluster_4_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_3_cluster_4_addr = proc_3_io_mem_cluster_4_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_3_cluster_5_en = proc_3_io_mem_cluster_5_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_3_cluster_5_addr = proc_3_io_mem_cluster_5_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_3_cluster_6_en = proc_3_io_mem_cluster_6_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_3_cluster_6_addr = proc_3_io_mem_cluster_6_addr; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_3_cluster_7_en = proc_3_io_mem_cluster_7_en; // @[ipsa.scala 70:37]
  assign sram_cluster_0_io_r_3_cluster_7_addr = proc_3_io_mem_cluster_7_addr; // @[ipsa.scala 70:37]
  assign init_clock = clock;
  assign init_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_header_0 = io_pipe_phv_in_header_0; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_header_1 = io_pipe_phv_in_header_1; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_header_2 = io_pipe_phv_in_header_2; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_header_3 = io_pipe_phv_in_header_3; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_header_4 = io_pipe_phv_in_header_4; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_header_5 = io_pipe_phv_in_header_5; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_header_6 = io_pipe_phv_in_header_6; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_header_7 = io_pipe_phv_in_header_7; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_header_8 = io_pipe_phv_in_header_8; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_header_9 = io_pipe_phv_in_header_9; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_header_10 = io_pipe_phv_in_header_10; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_header_11 = io_pipe_phv_in_header_11; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_header_12 = io_pipe_phv_in_header_12; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_header_13 = io_pipe_phv_in_header_13; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_header_14 = io_pipe_phv_in_header_14; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_header_15 = io_pipe_phv_in_header_15; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_parse_current_state = io_pipe_phv_in_parse_current_state; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_parse_current_offset = io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 75:25]
  assign init_io_pipe_phv_in_parse_transition_field = io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 75:25]
  assign init_io_first_proc_id = first_proc_id; // @[ipsa.scala 76:27]
  assign trans_0_clock = clock;
  assign trans_0_io_pipe_phv_in_data_0 = proc_0_io_pipe_phv_out_data_0; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_1 = proc_0_io_pipe_phv_out_data_1; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_2 = proc_0_io_pipe_phv_out_data_2; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_3 = proc_0_io_pipe_phv_out_data_3; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_4 = proc_0_io_pipe_phv_out_data_4; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_5 = proc_0_io_pipe_phv_out_data_5; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_6 = proc_0_io_pipe_phv_out_data_6; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_7 = proc_0_io_pipe_phv_out_data_7; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_8 = proc_0_io_pipe_phv_out_data_8; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_9 = proc_0_io_pipe_phv_out_data_9; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_10 = proc_0_io_pipe_phv_out_data_10; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_11 = proc_0_io_pipe_phv_out_data_11; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_12 = proc_0_io_pipe_phv_out_data_12; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_13 = proc_0_io_pipe_phv_out_data_13; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_14 = proc_0_io_pipe_phv_out_data_14; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_15 = proc_0_io_pipe_phv_out_data_15; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_16 = proc_0_io_pipe_phv_out_data_16; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_17 = proc_0_io_pipe_phv_out_data_17; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_18 = proc_0_io_pipe_phv_out_data_18; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_19 = proc_0_io_pipe_phv_out_data_19; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_20 = proc_0_io_pipe_phv_out_data_20; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_21 = proc_0_io_pipe_phv_out_data_21; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_22 = proc_0_io_pipe_phv_out_data_22; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_23 = proc_0_io_pipe_phv_out_data_23; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_24 = proc_0_io_pipe_phv_out_data_24; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_25 = proc_0_io_pipe_phv_out_data_25; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_26 = proc_0_io_pipe_phv_out_data_26; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_27 = proc_0_io_pipe_phv_out_data_27; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_28 = proc_0_io_pipe_phv_out_data_28; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_29 = proc_0_io_pipe_phv_out_data_29; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_30 = proc_0_io_pipe_phv_out_data_30; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_31 = proc_0_io_pipe_phv_out_data_31; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_32 = proc_0_io_pipe_phv_out_data_32; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_33 = proc_0_io_pipe_phv_out_data_33; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_34 = proc_0_io_pipe_phv_out_data_34; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_35 = proc_0_io_pipe_phv_out_data_35; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_36 = proc_0_io_pipe_phv_out_data_36; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_37 = proc_0_io_pipe_phv_out_data_37; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_38 = proc_0_io_pipe_phv_out_data_38; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_39 = proc_0_io_pipe_phv_out_data_39; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_40 = proc_0_io_pipe_phv_out_data_40; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_41 = proc_0_io_pipe_phv_out_data_41; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_42 = proc_0_io_pipe_phv_out_data_42; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_43 = proc_0_io_pipe_phv_out_data_43; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_44 = proc_0_io_pipe_phv_out_data_44; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_45 = proc_0_io_pipe_phv_out_data_45; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_46 = proc_0_io_pipe_phv_out_data_46; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_47 = proc_0_io_pipe_phv_out_data_47; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_48 = proc_0_io_pipe_phv_out_data_48; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_49 = proc_0_io_pipe_phv_out_data_49; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_50 = proc_0_io_pipe_phv_out_data_50; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_51 = proc_0_io_pipe_phv_out_data_51; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_52 = proc_0_io_pipe_phv_out_data_52; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_53 = proc_0_io_pipe_phv_out_data_53; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_54 = proc_0_io_pipe_phv_out_data_54; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_55 = proc_0_io_pipe_phv_out_data_55; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_56 = proc_0_io_pipe_phv_out_data_56; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_57 = proc_0_io_pipe_phv_out_data_57; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_58 = proc_0_io_pipe_phv_out_data_58; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_59 = proc_0_io_pipe_phv_out_data_59; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_60 = proc_0_io_pipe_phv_out_data_60; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_61 = proc_0_io_pipe_phv_out_data_61; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_62 = proc_0_io_pipe_phv_out_data_62; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_63 = proc_0_io_pipe_phv_out_data_63; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_64 = proc_0_io_pipe_phv_out_data_64; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_65 = proc_0_io_pipe_phv_out_data_65; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_66 = proc_0_io_pipe_phv_out_data_66; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_67 = proc_0_io_pipe_phv_out_data_67; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_68 = proc_0_io_pipe_phv_out_data_68; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_69 = proc_0_io_pipe_phv_out_data_69; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_70 = proc_0_io_pipe_phv_out_data_70; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_71 = proc_0_io_pipe_phv_out_data_71; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_72 = proc_0_io_pipe_phv_out_data_72; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_73 = proc_0_io_pipe_phv_out_data_73; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_74 = proc_0_io_pipe_phv_out_data_74; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_75 = proc_0_io_pipe_phv_out_data_75; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_76 = proc_0_io_pipe_phv_out_data_76; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_77 = proc_0_io_pipe_phv_out_data_77; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_78 = proc_0_io_pipe_phv_out_data_78; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_79 = proc_0_io_pipe_phv_out_data_79; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_80 = proc_0_io_pipe_phv_out_data_80; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_81 = proc_0_io_pipe_phv_out_data_81; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_82 = proc_0_io_pipe_phv_out_data_82; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_83 = proc_0_io_pipe_phv_out_data_83; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_84 = proc_0_io_pipe_phv_out_data_84; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_85 = proc_0_io_pipe_phv_out_data_85; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_86 = proc_0_io_pipe_phv_out_data_86; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_87 = proc_0_io_pipe_phv_out_data_87; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_88 = proc_0_io_pipe_phv_out_data_88; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_89 = proc_0_io_pipe_phv_out_data_89; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_90 = proc_0_io_pipe_phv_out_data_90; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_91 = proc_0_io_pipe_phv_out_data_91; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_92 = proc_0_io_pipe_phv_out_data_92; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_93 = proc_0_io_pipe_phv_out_data_93; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_94 = proc_0_io_pipe_phv_out_data_94; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_data_95 = proc_0_io_pipe_phv_out_data_95; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_0 = proc_0_io_pipe_phv_out_header_0; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_1 = proc_0_io_pipe_phv_out_header_1; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_2 = proc_0_io_pipe_phv_out_header_2; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_3 = proc_0_io_pipe_phv_out_header_3; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_4 = proc_0_io_pipe_phv_out_header_4; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_5 = proc_0_io_pipe_phv_out_header_5; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_6 = proc_0_io_pipe_phv_out_header_6; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_7 = proc_0_io_pipe_phv_out_header_7; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_8 = proc_0_io_pipe_phv_out_header_8; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_9 = proc_0_io_pipe_phv_out_header_9; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_10 = proc_0_io_pipe_phv_out_header_10; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_11 = proc_0_io_pipe_phv_out_header_11; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_12 = proc_0_io_pipe_phv_out_header_12; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_13 = proc_0_io_pipe_phv_out_header_13; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_14 = proc_0_io_pipe_phv_out_header_14; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_header_15 = proc_0_io_pipe_phv_out_header_15; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_parse_current_state = proc_0_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_parse_current_offset = proc_0_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_parse_transition_field = proc_0_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_next_processor_id = proc_0_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 82:32]
  assign trans_0_io_pipe_phv_in_next_config_id = proc_0_io_pipe_phv_out_next_config_id; // @[ipsa.scala 82:32]
  assign trans_0_io_next_proc_exist = last_proc_id != 2'h0; // @[ipsa.scala 80:48]
  assign trans_0_io_next_proc_id = next_proc_id_0; // @[ipsa.scala 81:32]
  assign trans_1_clock = clock;
  assign trans_1_io_pipe_phv_in_data_0 = proc_1_io_pipe_phv_out_data_0; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_1 = proc_1_io_pipe_phv_out_data_1; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_2 = proc_1_io_pipe_phv_out_data_2; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_3 = proc_1_io_pipe_phv_out_data_3; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_4 = proc_1_io_pipe_phv_out_data_4; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_5 = proc_1_io_pipe_phv_out_data_5; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_6 = proc_1_io_pipe_phv_out_data_6; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_7 = proc_1_io_pipe_phv_out_data_7; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_8 = proc_1_io_pipe_phv_out_data_8; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_9 = proc_1_io_pipe_phv_out_data_9; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_10 = proc_1_io_pipe_phv_out_data_10; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_11 = proc_1_io_pipe_phv_out_data_11; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_12 = proc_1_io_pipe_phv_out_data_12; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_13 = proc_1_io_pipe_phv_out_data_13; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_14 = proc_1_io_pipe_phv_out_data_14; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_15 = proc_1_io_pipe_phv_out_data_15; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_16 = proc_1_io_pipe_phv_out_data_16; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_17 = proc_1_io_pipe_phv_out_data_17; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_18 = proc_1_io_pipe_phv_out_data_18; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_19 = proc_1_io_pipe_phv_out_data_19; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_20 = proc_1_io_pipe_phv_out_data_20; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_21 = proc_1_io_pipe_phv_out_data_21; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_22 = proc_1_io_pipe_phv_out_data_22; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_23 = proc_1_io_pipe_phv_out_data_23; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_24 = proc_1_io_pipe_phv_out_data_24; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_25 = proc_1_io_pipe_phv_out_data_25; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_26 = proc_1_io_pipe_phv_out_data_26; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_27 = proc_1_io_pipe_phv_out_data_27; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_28 = proc_1_io_pipe_phv_out_data_28; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_29 = proc_1_io_pipe_phv_out_data_29; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_30 = proc_1_io_pipe_phv_out_data_30; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_31 = proc_1_io_pipe_phv_out_data_31; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_32 = proc_1_io_pipe_phv_out_data_32; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_33 = proc_1_io_pipe_phv_out_data_33; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_34 = proc_1_io_pipe_phv_out_data_34; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_35 = proc_1_io_pipe_phv_out_data_35; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_36 = proc_1_io_pipe_phv_out_data_36; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_37 = proc_1_io_pipe_phv_out_data_37; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_38 = proc_1_io_pipe_phv_out_data_38; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_39 = proc_1_io_pipe_phv_out_data_39; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_40 = proc_1_io_pipe_phv_out_data_40; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_41 = proc_1_io_pipe_phv_out_data_41; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_42 = proc_1_io_pipe_phv_out_data_42; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_43 = proc_1_io_pipe_phv_out_data_43; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_44 = proc_1_io_pipe_phv_out_data_44; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_45 = proc_1_io_pipe_phv_out_data_45; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_46 = proc_1_io_pipe_phv_out_data_46; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_47 = proc_1_io_pipe_phv_out_data_47; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_48 = proc_1_io_pipe_phv_out_data_48; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_49 = proc_1_io_pipe_phv_out_data_49; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_50 = proc_1_io_pipe_phv_out_data_50; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_51 = proc_1_io_pipe_phv_out_data_51; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_52 = proc_1_io_pipe_phv_out_data_52; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_53 = proc_1_io_pipe_phv_out_data_53; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_54 = proc_1_io_pipe_phv_out_data_54; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_55 = proc_1_io_pipe_phv_out_data_55; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_56 = proc_1_io_pipe_phv_out_data_56; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_57 = proc_1_io_pipe_phv_out_data_57; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_58 = proc_1_io_pipe_phv_out_data_58; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_59 = proc_1_io_pipe_phv_out_data_59; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_60 = proc_1_io_pipe_phv_out_data_60; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_61 = proc_1_io_pipe_phv_out_data_61; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_62 = proc_1_io_pipe_phv_out_data_62; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_63 = proc_1_io_pipe_phv_out_data_63; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_64 = proc_1_io_pipe_phv_out_data_64; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_65 = proc_1_io_pipe_phv_out_data_65; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_66 = proc_1_io_pipe_phv_out_data_66; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_67 = proc_1_io_pipe_phv_out_data_67; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_68 = proc_1_io_pipe_phv_out_data_68; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_69 = proc_1_io_pipe_phv_out_data_69; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_70 = proc_1_io_pipe_phv_out_data_70; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_71 = proc_1_io_pipe_phv_out_data_71; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_72 = proc_1_io_pipe_phv_out_data_72; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_73 = proc_1_io_pipe_phv_out_data_73; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_74 = proc_1_io_pipe_phv_out_data_74; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_75 = proc_1_io_pipe_phv_out_data_75; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_76 = proc_1_io_pipe_phv_out_data_76; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_77 = proc_1_io_pipe_phv_out_data_77; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_78 = proc_1_io_pipe_phv_out_data_78; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_79 = proc_1_io_pipe_phv_out_data_79; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_80 = proc_1_io_pipe_phv_out_data_80; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_81 = proc_1_io_pipe_phv_out_data_81; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_82 = proc_1_io_pipe_phv_out_data_82; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_83 = proc_1_io_pipe_phv_out_data_83; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_84 = proc_1_io_pipe_phv_out_data_84; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_85 = proc_1_io_pipe_phv_out_data_85; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_86 = proc_1_io_pipe_phv_out_data_86; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_87 = proc_1_io_pipe_phv_out_data_87; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_88 = proc_1_io_pipe_phv_out_data_88; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_89 = proc_1_io_pipe_phv_out_data_89; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_90 = proc_1_io_pipe_phv_out_data_90; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_91 = proc_1_io_pipe_phv_out_data_91; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_92 = proc_1_io_pipe_phv_out_data_92; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_93 = proc_1_io_pipe_phv_out_data_93; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_94 = proc_1_io_pipe_phv_out_data_94; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_data_95 = proc_1_io_pipe_phv_out_data_95; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_0 = proc_1_io_pipe_phv_out_header_0; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_1 = proc_1_io_pipe_phv_out_header_1; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_2 = proc_1_io_pipe_phv_out_header_2; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_3 = proc_1_io_pipe_phv_out_header_3; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_4 = proc_1_io_pipe_phv_out_header_4; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_5 = proc_1_io_pipe_phv_out_header_5; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_6 = proc_1_io_pipe_phv_out_header_6; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_7 = proc_1_io_pipe_phv_out_header_7; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_8 = proc_1_io_pipe_phv_out_header_8; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_9 = proc_1_io_pipe_phv_out_header_9; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_10 = proc_1_io_pipe_phv_out_header_10; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_11 = proc_1_io_pipe_phv_out_header_11; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_12 = proc_1_io_pipe_phv_out_header_12; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_13 = proc_1_io_pipe_phv_out_header_13; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_14 = proc_1_io_pipe_phv_out_header_14; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_header_15 = proc_1_io_pipe_phv_out_header_15; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_parse_current_state = proc_1_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_parse_current_offset = proc_1_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_parse_transition_field = proc_1_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_next_processor_id = proc_1_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 82:32]
  assign trans_1_io_pipe_phv_in_next_config_id = proc_1_io_pipe_phv_out_next_config_id; // @[ipsa.scala 82:32]
  assign trans_1_io_next_proc_exist = last_proc_id != 2'h1; // @[ipsa.scala 80:48]
  assign trans_1_io_next_proc_id = next_proc_id_1; // @[ipsa.scala 81:32]
  assign trans_2_clock = clock;
  assign trans_2_io_pipe_phv_in_data_0 = proc_2_io_pipe_phv_out_data_0; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_1 = proc_2_io_pipe_phv_out_data_1; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_2 = proc_2_io_pipe_phv_out_data_2; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_3 = proc_2_io_pipe_phv_out_data_3; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_4 = proc_2_io_pipe_phv_out_data_4; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_5 = proc_2_io_pipe_phv_out_data_5; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_6 = proc_2_io_pipe_phv_out_data_6; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_7 = proc_2_io_pipe_phv_out_data_7; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_8 = proc_2_io_pipe_phv_out_data_8; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_9 = proc_2_io_pipe_phv_out_data_9; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_10 = proc_2_io_pipe_phv_out_data_10; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_11 = proc_2_io_pipe_phv_out_data_11; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_12 = proc_2_io_pipe_phv_out_data_12; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_13 = proc_2_io_pipe_phv_out_data_13; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_14 = proc_2_io_pipe_phv_out_data_14; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_15 = proc_2_io_pipe_phv_out_data_15; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_16 = proc_2_io_pipe_phv_out_data_16; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_17 = proc_2_io_pipe_phv_out_data_17; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_18 = proc_2_io_pipe_phv_out_data_18; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_19 = proc_2_io_pipe_phv_out_data_19; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_20 = proc_2_io_pipe_phv_out_data_20; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_21 = proc_2_io_pipe_phv_out_data_21; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_22 = proc_2_io_pipe_phv_out_data_22; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_23 = proc_2_io_pipe_phv_out_data_23; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_24 = proc_2_io_pipe_phv_out_data_24; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_25 = proc_2_io_pipe_phv_out_data_25; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_26 = proc_2_io_pipe_phv_out_data_26; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_27 = proc_2_io_pipe_phv_out_data_27; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_28 = proc_2_io_pipe_phv_out_data_28; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_29 = proc_2_io_pipe_phv_out_data_29; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_30 = proc_2_io_pipe_phv_out_data_30; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_31 = proc_2_io_pipe_phv_out_data_31; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_32 = proc_2_io_pipe_phv_out_data_32; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_33 = proc_2_io_pipe_phv_out_data_33; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_34 = proc_2_io_pipe_phv_out_data_34; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_35 = proc_2_io_pipe_phv_out_data_35; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_36 = proc_2_io_pipe_phv_out_data_36; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_37 = proc_2_io_pipe_phv_out_data_37; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_38 = proc_2_io_pipe_phv_out_data_38; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_39 = proc_2_io_pipe_phv_out_data_39; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_40 = proc_2_io_pipe_phv_out_data_40; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_41 = proc_2_io_pipe_phv_out_data_41; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_42 = proc_2_io_pipe_phv_out_data_42; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_43 = proc_2_io_pipe_phv_out_data_43; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_44 = proc_2_io_pipe_phv_out_data_44; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_45 = proc_2_io_pipe_phv_out_data_45; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_46 = proc_2_io_pipe_phv_out_data_46; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_47 = proc_2_io_pipe_phv_out_data_47; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_48 = proc_2_io_pipe_phv_out_data_48; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_49 = proc_2_io_pipe_phv_out_data_49; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_50 = proc_2_io_pipe_phv_out_data_50; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_51 = proc_2_io_pipe_phv_out_data_51; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_52 = proc_2_io_pipe_phv_out_data_52; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_53 = proc_2_io_pipe_phv_out_data_53; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_54 = proc_2_io_pipe_phv_out_data_54; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_55 = proc_2_io_pipe_phv_out_data_55; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_56 = proc_2_io_pipe_phv_out_data_56; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_57 = proc_2_io_pipe_phv_out_data_57; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_58 = proc_2_io_pipe_phv_out_data_58; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_59 = proc_2_io_pipe_phv_out_data_59; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_60 = proc_2_io_pipe_phv_out_data_60; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_61 = proc_2_io_pipe_phv_out_data_61; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_62 = proc_2_io_pipe_phv_out_data_62; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_63 = proc_2_io_pipe_phv_out_data_63; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_64 = proc_2_io_pipe_phv_out_data_64; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_65 = proc_2_io_pipe_phv_out_data_65; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_66 = proc_2_io_pipe_phv_out_data_66; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_67 = proc_2_io_pipe_phv_out_data_67; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_68 = proc_2_io_pipe_phv_out_data_68; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_69 = proc_2_io_pipe_phv_out_data_69; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_70 = proc_2_io_pipe_phv_out_data_70; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_71 = proc_2_io_pipe_phv_out_data_71; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_72 = proc_2_io_pipe_phv_out_data_72; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_73 = proc_2_io_pipe_phv_out_data_73; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_74 = proc_2_io_pipe_phv_out_data_74; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_75 = proc_2_io_pipe_phv_out_data_75; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_76 = proc_2_io_pipe_phv_out_data_76; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_77 = proc_2_io_pipe_phv_out_data_77; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_78 = proc_2_io_pipe_phv_out_data_78; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_79 = proc_2_io_pipe_phv_out_data_79; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_80 = proc_2_io_pipe_phv_out_data_80; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_81 = proc_2_io_pipe_phv_out_data_81; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_82 = proc_2_io_pipe_phv_out_data_82; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_83 = proc_2_io_pipe_phv_out_data_83; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_84 = proc_2_io_pipe_phv_out_data_84; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_85 = proc_2_io_pipe_phv_out_data_85; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_86 = proc_2_io_pipe_phv_out_data_86; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_87 = proc_2_io_pipe_phv_out_data_87; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_88 = proc_2_io_pipe_phv_out_data_88; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_89 = proc_2_io_pipe_phv_out_data_89; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_90 = proc_2_io_pipe_phv_out_data_90; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_91 = proc_2_io_pipe_phv_out_data_91; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_92 = proc_2_io_pipe_phv_out_data_92; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_93 = proc_2_io_pipe_phv_out_data_93; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_94 = proc_2_io_pipe_phv_out_data_94; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_data_95 = proc_2_io_pipe_phv_out_data_95; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_0 = proc_2_io_pipe_phv_out_header_0; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_1 = proc_2_io_pipe_phv_out_header_1; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_2 = proc_2_io_pipe_phv_out_header_2; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_3 = proc_2_io_pipe_phv_out_header_3; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_4 = proc_2_io_pipe_phv_out_header_4; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_5 = proc_2_io_pipe_phv_out_header_5; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_6 = proc_2_io_pipe_phv_out_header_6; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_7 = proc_2_io_pipe_phv_out_header_7; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_8 = proc_2_io_pipe_phv_out_header_8; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_9 = proc_2_io_pipe_phv_out_header_9; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_10 = proc_2_io_pipe_phv_out_header_10; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_11 = proc_2_io_pipe_phv_out_header_11; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_12 = proc_2_io_pipe_phv_out_header_12; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_13 = proc_2_io_pipe_phv_out_header_13; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_14 = proc_2_io_pipe_phv_out_header_14; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_header_15 = proc_2_io_pipe_phv_out_header_15; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_parse_current_state = proc_2_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_parse_current_offset = proc_2_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_parse_transition_field = proc_2_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_next_processor_id = proc_2_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 82:32]
  assign trans_2_io_pipe_phv_in_next_config_id = proc_2_io_pipe_phv_out_next_config_id; // @[ipsa.scala 82:32]
  assign trans_2_io_next_proc_exist = last_proc_id != 2'h2; // @[ipsa.scala 80:48]
  assign trans_2_io_next_proc_id = next_proc_id_2; // @[ipsa.scala 81:32]
  assign trans_3_clock = clock;
  assign trans_3_io_pipe_phv_in_data_0 = proc_3_io_pipe_phv_out_data_0; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_1 = proc_3_io_pipe_phv_out_data_1; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_2 = proc_3_io_pipe_phv_out_data_2; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_3 = proc_3_io_pipe_phv_out_data_3; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_4 = proc_3_io_pipe_phv_out_data_4; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_5 = proc_3_io_pipe_phv_out_data_5; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_6 = proc_3_io_pipe_phv_out_data_6; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_7 = proc_3_io_pipe_phv_out_data_7; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_8 = proc_3_io_pipe_phv_out_data_8; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_9 = proc_3_io_pipe_phv_out_data_9; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_10 = proc_3_io_pipe_phv_out_data_10; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_11 = proc_3_io_pipe_phv_out_data_11; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_12 = proc_3_io_pipe_phv_out_data_12; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_13 = proc_3_io_pipe_phv_out_data_13; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_14 = proc_3_io_pipe_phv_out_data_14; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_15 = proc_3_io_pipe_phv_out_data_15; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_16 = proc_3_io_pipe_phv_out_data_16; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_17 = proc_3_io_pipe_phv_out_data_17; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_18 = proc_3_io_pipe_phv_out_data_18; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_19 = proc_3_io_pipe_phv_out_data_19; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_20 = proc_3_io_pipe_phv_out_data_20; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_21 = proc_3_io_pipe_phv_out_data_21; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_22 = proc_3_io_pipe_phv_out_data_22; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_23 = proc_3_io_pipe_phv_out_data_23; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_24 = proc_3_io_pipe_phv_out_data_24; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_25 = proc_3_io_pipe_phv_out_data_25; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_26 = proc_3_io_pipe_phv_out_data_26; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_27 = proc_3_io_pipe_phv_out_data_27; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_28 = proc_3_io_pipe_phv_out_data_28; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_29 = proc_3_io_pipe_phv_out_data_29; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_30 = proc_3_io_pipe_phv_out_data_30; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_31 = proc_3_io_pipe_phv_out_data_31; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_32 = proc_3_io_pipe_phv_out_data_32; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_33 = proc_3_io_pipe_phv_out_data_33; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_34 = proc_3_io_pipe_phv_out_data_34; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_35 = proc_3_io_pipe_phv_out_data_35; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_36 = proc_3_io_pipe_phv_out_data_36; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_37 = proc_3_io_pipe_phv_out_data_37; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_38 = proc_3_io_pipe_phv_out_data_38; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_39 = proc_3_io_pipe_phv_out_data_39; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_40 = proc_3_io_pipe_phv_out_data_40; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_41 = proc_3_io_pipe_phv_out_data_41; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_42 = proc_3_io_pipe_phv_out_data_42; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_43 = proc_3_io_pipe_phv_out_data_43; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_44 = proc_3_io_pipe_phv_out_data_44; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_45 = proc_3_io_pipe_phv_out_data_45; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_46 = proc_3_io_pipe_phv_out_data_46; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_47 = proc_3_io_pipe_phv_out_data_47; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_48 = proc_3_io_pipe_phv_out_data_48; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_49 = proc_3_io_pipe_phv_out_data_49; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_50 = proc_3_io_pipe_phv_out_data_50; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_51 = proc_3_io_pipe_phv_out_data_51; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_52 = proc_3_io_pipe_phv_out_data_52; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_53 = proc_3_io_pipe_phv_out_data_53; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_54 = proc_3_io_pipe_phv_out_data_54; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_55 = proc_3_io_pipe_phv_out_data_55; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_56 = proc_3_io_pipe_phv_out_data_56; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_57 = proc_3_io_pipe_phv_out_data_57; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_58 = proc_3_io_pipe_phv_out_data_58; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_59 = proc_3_io_pipe_phv_out_data_59; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_60 = proc_3_io_pipe_phv_out_data_60; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_61 = proc_3_io_pipe_phv_out_data_61; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_62 = proc_3_io_pipe_phv_out_data_62; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_63 = proc_3_io_pipe_phv_out_data_63; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_64 = proc_3_io_pipe_phv_out_data_64; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_65 = proc_3_io_pipe_phv_out_data_65; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_66 = proc_3_io_pipe_phv_out_data_66; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_67 = proc_3_io_pipe_phv_out_data_67; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_68 = proc_3_io_pipe_phv_out_data_68; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_69 = proc_3_io_pipe_phv_out_data_69; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_70 = proc_3_io_pipe_phv_out_data_70; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_71 = proc_3_io_pipe_phv_out_data_71; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_72 = proc_3_io_pipe_phv_out_data_72; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_73 = proc_3_io_pipe_phv_out_data_73; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_74 = proc_3_io_pipe_phv_out_data_74; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_75 = proc_3_io_pipe_phv_out_data_75; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_76 = proc_3_io_pipe_phv_out_data_76; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_77 = proc_3_io_pipe_phv_out_data_77; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_78 = proc_3_io_pipe_phv_out_data_78; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_79 = proc_3_io_pipe_phv_out_data_79; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_80 = proc_3_io_pipe_phv_out_data_80; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_81 = proc_3_io_pipe_phv_out_data_81; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_82 = proc_3_io_pipe_phv_out_data_82; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_83 = proc_3_io_pipe_phv_out_data_83; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_84 = proc_3_io_pipe_phv_out_data_84; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_85 = proc_3_io_pipe_phv_out_data_85; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_86 = proc_3_io_pipe_phv_out_data_86; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_87 = proc_3_io_pipe_phv_out_data_87; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_88 = proc_3_io_pipe_phv_out_data_88; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_89 = proc_3_io_pipe_phv_out_data_89; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_90 = proc_3_io_pipe_phv_out_data_90; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_91 = proc_3_io_pipe_phv_out_data_91; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_92 = proc_3_io_pipe_phv_out_data_92; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_93 = proc_3_io_pipe_phv_out_data_93; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_94 = proc_3_io_pipe_phv_out_data_94; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_data_95 = proc_3_io_pipe_phv_out_data_95; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_0 = proc_3_io_pipe_phv_out_header_0; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_1 = proc_3_io_pipe_phv_out_header_1; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_2 = proc_3_io_pipe_phv_out_header_2; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_3 = proc_3_io_pipe_phv_out_header_3; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_4 = proc_3_io_pipe_phv_out_header_4; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_5 = proc_3_io_pipe_phv_out_header_5; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_6 = proc_3_io_pipe_phv_out_header_6; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_7 = proc_3_io_pipe_phv_out_header_7; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_8 = proc_3_io_pipe_phv_out_header_8; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_9 = proc_3_io_pipe_phv_out_header_9; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_10 = proc_3_io_pipe_phv_out_header_10; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_11 = proc_3_io_pipe_phv_out_header_11; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_12 = proc_3_io_pipe_phv_out_header_12; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_13 = proc_3_io_pipe_phv_out_header_13; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_14 = proc_3_io_pipe_phv_out_header_14; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_header_15 = proc_3_io_pipe_phv_out_header_15; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_parse_current_state = proc_3_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_parse_current_offset = proc_3_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_parse_transition_field = proc_3_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_next_processor_id = proc_3_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 82:32]
  assign trans_3_io_pipe_phv_in_next_config_id = proc_3_io_pipe_phv_out_next_config_id; // @[ipsa.scala 82:32]
  assign trans_3_io_next_proc_exist = last_proc_id != 2'h3; // @[ipsa.scala 80:48]
  assign trans_3_io_next_proc_id = next_proc_id_3; // @[ipsa.scala 81:32]
  always @(posedge clock) begin
    if (io_mod_xbar_mod_en) begin // @[ipsa.scala 47:31]
      first_proc_id <= io_mod_xbar_mod_first_proc_id; // @[ipsa.scala 48:23]
    end
    if (io_mod_xbar_mod_en) begin // @[ipsa.scala 47:31]
      last_proc_id <= io_mod_xbar_mod_last_proc_id; // @[ipsa.scala 49:23]
    end
    if (io_mod_xbar_mod_en) begin // @[ipsa.scala 47:31]
      next_proc_id_0 <= io_mod_xbar_mod_next_proc_id_0; // @[ipsa.scala 51:29]
    end
    if (io_mod_xbar_mod_en) begin // @[ipsa.scala 47:31]
      next_proc_id_1 <= io_mod_xbar_mod_next_proc_id_1; // @[ipsa.scala 51:29]
    end
    if (io_mod_xbar_mod_en) begin // @[ipsa.scala 47:31]
      next_proc_id_2 <= io_mod_xbar_mod_next_proc_id_2; // @[ipsa.scala 51:29]
    end
    if (io_mod_xbar_mod_en) begin // @[ipsa.scala 47:31]
      next_proc_id_3 <= io_mod_xbar_mod_next_proc_id_3; // @[ipsa.scala 51:29]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  first_proc_id = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  last_proc_id = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  next_proc_id_0 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  next_proc_id_1 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  next_proc_id_2 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  next_proc_id_3 = _RAND_5[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
