module MatchGetKeyPISA(
  input          clock,
  input  [7:0]   io_pipe_phv_in_data_0,
  input  [7:0]   io_pipe_phv_in_data_1,
  input  [7:0]   io_pipe_phv_in_data_2,
  input  [7:0]   io_pipe_phv_in_data_3,
  input  [7:0]   io_pipe_phv_in_data_4,
  input  [7:0]   io_pipe_phv_in_data_5,
  input  [7:0]   io_pipe_phv_in_data_6,
  input  [7:0]   io_pipe_phv_in_data_7,
  input  [7:0]   io_pipe_phv_in_data_8,
  input  [7:0]   io_pipe_phv_in_data_9,
  input  [7:0]   io_pipe_phv_in_data_10,
  input  [7:0]   io_pipe_phv_in_data_11,
  input  [7:0]   io_pipe_phv_in_data_12,
  input  [7:0]   io_pipe_phv_in_data_13,
  input  [7:0]   io_pipe_phv_in_data_14,
  input  [7:0]   io_pipe_phv_in_data_15,
  input  [7:0]   io_pipe_phv_in_data_16,
  input  [7:0]   io_pipe_phv_in_data_17,
  input  [7:0]   io_pipe_phv_in_data_18,
  input  [7:0]   io_pipe_phv_in_data_19,
  input  [7:0]   io_pipe_phv_in_data_20,
  input  [7:0]   io_pipe_phv_in_data_21,
  input  [7:0]   io_pipe_phv_in_data_22,
  input  [7:0]   io_pipe_phv_in_data_23,
  input  [7:0]   io_pipe_phv_in_data_24,
  input  [7:0]   io_pipe_phv_in_data_25,
  input  [7:0]   io_pipe_phv_in_data_26,
  input  [7:0]   io_pipe_phv_in_data_27,
  input  [7:0]   io_pipe_phv_in_data_28,
  input  [7:0]   io_pipe_phv_in_data_29,
  input  [7:0]   io_pipe_phv_in_data_30,
  input  [7:0]   io_pipe_phv_in_data_31,
  input  [7:0]   io_pipe_phv_in_data_32,
  input  [7:0]   io_pipe_phv_in_data_33,
  input  [7:0]   io_pipe_phv_in_data_34,
  input  [7:0]   io_pipe_phv_in_data_35,
  input  [7:0]   io_pipe_phv_in_data_36,
  input  [7:0]   io_pipe_phv_in_data_37,
  input  [7:0]   io_pipe_phv_in_data_38,
  input  [7:0]   io_pipe_phv_in_data_39,
  input  [7:0]   io_pipe_phv_in_data_40,
  input  [7:0]   io_pipe_phv_in_data_41,
  input  [7:0]   io_pipe_phv_in_data_42,
  input  [7:0]   io_pipe_phv_in_data_43,
  input  [7:0]   io_pipe_phv_in_data_44,
  input  [7:0]   io_pipe_phv_in_data_45,
  input  [7:0]   io_pipe_phv_in_data_46,
  input  [7:0]   io_pipe_phv_in_data_47,
  input  [7:0]   io_pipe_phv_in_data_48,
  input  [7:0]   io_pipe_phv_in_data_49,
  input  [7:0]   io_pipe_phv_in_data_50,
  input  [7:0]   io_pipe_phv_in_data_51,
  input  [7:0]   io_pipe_phv_in_data_52,
  input  [7:0]   io_pipe_phv_in_data_53,
  input  [7:0]   io_pipe_phv_in_data_54,
  input  [7:0]   io_pipe_phv_in_data_55,
  input  [7:0]   io_pipe_phv_in_data_56,
  input  [7:0]   io_pipe_phv_in_data_57,
  input  [7:0]   io_pipe_phv_in_data_58,
  input  [7:0]   io_pipe_phv_in_data_59,
  input  [7:0]   io_pipe_phv_in_data_60,
  input  [7:0]   io_pipe_phv_in_data_61,
  input  [7:0]   io_pipe_phv_in_data_62,
  input  [7:0]   io_pipe_phv_in_data_63,
  input  [7:0]   io_pipe_phv_in_data_64,
  input  [7:0]   io_pipe_phv_in_data_65,
  input  [7:0]   io_pipe_phv_in_data_66,
  input  [7:0]   io_pipe_phv_in_data_67,
  input  [7:0]   io_pipe_phv_in_data_68,
  input  [7:0]   io_pipe_phv_in_data_69,
  input  [7:0]   io_pipe_phv_in_data_70,
  input  [7:0]   io_pipe_phv_in_data_71,
  input  [7:0]   io_pipe_phv_in_data_72,
  input  [7:0]   io_pipe_phv_in_data_73,
  input  [7:0]   io_pipe_phv_in_data_74,
  input  [7:0]   io_pipe_phv_in_data_75,
  input  [7:0]   io_pipe_phv_in_data_76,
  input  [7:0]   io_pipe_phv_in_data_77,
  input  [7:0]   io_pipe_phv_in_data_78,
  input  [7:0]   io_pipe_phv_in_data_79,
  input  [7:0]   io_pipe_phv_in_data_80,
  input  [7:0]   io_pipe_phv_in_data_81,
  input  [7:0]   io_pipe_phv_in_data_82,
  input  [7:0]   io_pipe_phv_in_data_83,
  input  [7:0]   io_pipe_phv_in_data_84,
  input  [7:0]   io_pipe_phv_in_data_85,
  input  [7:0]   io_pipe_phv_in_data_86,
  input  [7:0]   io_pipe_phv_in_data_87,
  input  [7:0]   io_pipe_phv_in_data_88,
  input  [7:0]   io_pipe_phv_in_data_89,
  input  [7:0]   io_pipe_phv_in_data_90,
  input  [7:0]   io_pipe_phv_in_data_91,
  input  [7:0]   io_pipe_phv_in_data_92,
  input  [7:0]   io_pipe_phv_in_data_93,
  input  [7:0]   io_pipe_phv_in_data_94,
  input  [7:0]   io_pipe_phv_in_data_95,
  input  [7:0]   io_pipe_phv_in_data_96,
  input  [7:0]   io_pipe_phv_in_data_97,
  input  [7:0]   io_pipe_phv_in_data_98,
  input  [7:0]   io_pipe_phv_in_data_99,
  input  [7:0]   io_pipe_phv_in_data_100,
  input  [7:0]   io_pipe_phv_in_data_101,
  input  [7:0]   io_pipe_phv_in_data_102,
  input  [7:0]   io_pipe_phv_in_data_103,
  input  [7:0]   io_pipe_phv_in_data_104,
  input  [7:0]   io_pipe_phv_in_data_105,
  input  [7:0]   io_pipe_phv_in_data_106,
  input  [7:0]   io_pipe_phv_in_data_107,
  input  [7:0]   io_pipe_phv_in_data_108,
  input  [7:0]   io_pipe_phv_in_data_109,
  input  [7:0]   io_pipe_phv_in_data_110,
  input  [7:0]   io_pipe_phv_in_data_111,
  input  [7:0]   io_pipe_phv_in_data_112,
  input  [7:0]   io_pipe_phv_in_data_113,
  input  [7:0]   io_pipe_phv_in_data_114,
  input  [7:0]   io_pipe_phv_in_data_115,
  input  [7:0]   io_pipe_phv_in_data_116,
  input  [7:0]   io_pipe_phv_in_data_117,
  input  [7:0]   io_pipe_phv_in_data_118,
  input  [7:0]   io_pipe_phv_in_data_119,
  input  [7:0]   io_pipe_phv_in_data_120,
  input  [7:0]   io_pipe_phv_in_data_121,
  input  [7:0]   io_pipe_phv_in_data_122,
  input  [7:0]   io_pipe_phv_in_data_123,
  input  [7:0]   io_pipe_phv_in_data_124,
  input  [7:0]   io_pipe_phv_in_data_125,
  input  [7:0]   io_pipe_phv_in_data_126,
  input  [7:0]   io_pipe_phv_in_data_127,
  input  [7:0]   io_pipe_phv_in_data_128,
  input  [7:0]   io_pipe_phv_in_data_129,
  input  [7:0]   io_pipe_phv_in_data_130,
  input  [7:0]   io_pipe_phv_in_data_131,
  input  [7:0]   io_pipe_phv_in_data_132,
  input  [7:0]   io_pipe_phv_in_data_133,
  input  [7:0]   io_pipe_phv_in_data_134,
  input  [7:0]   io_pipe_phv_in_data_135,
  input  [7:0]   io_pipe_phv_in_data_136,
  input  [7:0]   io_pipe_phv_in_data_137,
  input  [7:0]   io_pipe_phv_in_data_138,
  input  [7:0]   io_pipe_phv_in_data_139,
  input  [7:0]   io_pipe_phv_in_data_140,
  input  [7:0]   io_pipe_phv_in_data_141,
  input  [7:0]   io_pipe_phv_in_data_142,
  input  [7:0]   io_pipe_phv_in_data_143,
  input  [7:0]   io_pipe_phv_in_data_144,
  input  [7:0]   io_pipe_phv_in_data_145,
  input  [7:0]   io_pipe_phv_in_data_146,
  input  [7:0]   io_pipe_phv_in_data_147,
  input  [7:0]   io_pipe_phv_in_data_148,
  input  [7:0]   io_pipe_phv_in_data_149,
  input  [7:0]   io_pipe_phv_in_data_150,
  input  [7:0]   io_pipe_phv_in_data_151,
  input  [7:0]   io_pipe_phv_in_data_152,
  input  [7:0]   io_pipe_phv_in_data_153,
  input  [7:0]   io_pipe_phv_in_data_154,
  input  [7:0]   io_pipe_phv_in_data_155,
  input  [7:0]   io_pipe_phv_in_data_156,
  input  [7:0]   io_pipe_phv_in_data_157,
  input  [7:0]   io_pipe_phv_in_data_158,
  input  [7:0]   io_pipe_phv_in_data_159,
  input  [7:0]   io_pipe_phv_in_data_160,
  input  [7:0]   io_pipe_phv_in_data_161,
  input  [7:0]   io_pipe_phv_in_data_162,
  input  [7:0]   io_pipe_phv_in_data_163,
  input  [7:0]   io_pipe_phv_in_data_164,
  input  [7:0]   io_pipe_phv_in_data_165,
  input  [7:0]   io_pipe_phv_in_data_166,
  input  [7:0]   io_pipe_phv_in_data_167,
  input  [7:0]   io_pipe_phv_in_data_168,
  input  [7:0]   io_pipe_phv_in_data_169,
  input  [7:0]   io_pipe_phv_in_data_170,
  input  [7:0]   io_pipe_phv_in_data_171,
  input  [7:0]   io_pipe_phv_in_data_172,
  input  [7:0]   io_pipe_phv_in_data_173,
  input  [7:0]   io_pipe_phv_in_data_174,
  input  [7:0]   io_pipe_phv_in_data_175,
  input  [7:0]   io_pipe_phv_in_data_176,
  input  [7:0]   io_pipe_phv_in_data_177,
  input  [7:0]   io_pipe_phv_in_data_178,
  input  [7:0]   io_pipe_phv_in_data_179,
  input  [7:0]   io_pipe_phv_in_data_180,
  input  [7:0]   io_pipe_phv_in_data_181,
  input  [7:0]   io_pipe_phv_in_data_182,
  input  [7:0]   io_pipe_phv_in_data_183,
  input  [7:0]   io_pipe_phv_in_data_184,
  input  [7:0]   io_pipe_phv_in_data_185,
  input  [7:0]   io_pipe_phv_in_data_186,
  input  [7:0]   io_pipe_phv_in_data_187,
  input  [7:0]   io_pipe_phv_in_data_188,
  input  [7:0]   io_pipe_phv_in_data_189,
  input  [7:0]   io_pipe_phv_in_data_190,
  input  [7:0]   io_pipe_phv_in_data_191,
  input  [7:0]   io_pipe_phv_in_data_192,
  input  [7:0]   io_pipe_phv_in_data_193,
  input  [7:0]   io_pipe_phv_in_data_194,
  input  [7:0]   io_pipe_phv_in_data_195,
  input  [7:0]   io_pipe_phv_in_data_196,
  input  [7:0]   io_pipe_phv_in_data_197,
  input  [7:0]   io_pipe_phv_in_data_198,
  input  [7:0]   io_pipe_phv_in_data_199,
  input  [7:0]   io_pipe_phv_in_data_200,
  input  [7:0]   io_pipe_phv_in_data_201,
  input  [7:0]   io_pipe_phv_in_data_202,
  input  [7:0]   io_pipe_phv_in_data_203,
  input  [7:0]   io_pipe_phv_in_data_204,
  input  [7:0]   io_pipe_phv_in_data_205,
  input  [7:0]   io_pipe_phv_in_data_206,
  input  [7:0]   io_pipe_phv_in_data_207,
  input  [7:0]   io_pipe_phv_in_data_208,
  input  [7:0]   io_pipe_phv_in_data_209,
  input  [7:0]   io_pipe_phv_in_data_210,
  input  [7:0]   io_pipe_phv_in_data_211,
  input  [7:0]   io_pipe_phv_in_data_212,
  input  [7:0]   io_pipe_phv_in_data_213,
  input  [7:0]   io_pipe_phv_in_data_214,
  input  [7:0]   io_pipe_phv_in_data_215,
  input  [7:0]   io_pipe_phv_in_data_216,
  input  [7:0]   io_pipe_phv_in_data_217,
  input  [7:0]   io_pipe_phv_in_data_218,
  input  [7:0]   io_pipe_phv_in_data_219,
  input  [7:0]   io_pipe_phv_in_data_220,
  input  [7:0]   io_pipe_phv_in_data_221,
  input  [7:0]   io_pipe_phv_in_data_222,
  input  [7:0]   io_pipe_phv_in_data_223,
  input  [7:0]   io_pipe_phv_in_data_224,
  input  [7:0]   io_pipe_phv_in_data_225,
  input  [7:0]   io_pipe_phv_in_data_226,
  input  [7:0]   io_pipe_phv_in_data_227,
  input  [7:0]   io_pipe_phv_in_data_228,
  input  [7:0]   io_pipe_phv_in_data_229,
  input  [7:0]   io_pipe_phv_in_data_230,
  input  [7:0]   io_pipe_phv_in_data_231,
  input  [7:0]   io_pipe_phv_in_data_232,
  input  [7:0]   io_pipe_phv_in_data_233,
  input  [7:0]   io_pipe_phv_in_data_234,
  input  [7:0]   io_pipe_phv_in_data_235,
  input  [7:0]   io_pipe_phv_in_data_236,
  input  [7:0]   io_pipe_phv_in_data_237,
  input  [7:0]   io_pipe_phv_in_data_238,
  input  [7:0]   io_pipe_phv_in_data_239,
  input  [7:0]   io_pipe_phv_in_data_240,
  input  [7:0]   io_pipe_phv_in_data_241,
  input  [7:0]   io_pipe_phv_in_data_242,
  input  [7:0]   io_pipe_phv_in_data_243,
  input  [7:0]   io_pipe_phv_in_data_244,
  input  [7:0]   io_pipe_phv_in_data_245,
  input  [7:0]   io_pipe_phv_in_data_246,
  input  [7:0]   io_pipe_phv_in_data_247,
  input  [7:0]   io_pipe_phv_in_data_248,
  input  [7:0]   io_pipe_phv_in_data_249,
  input  [7:0]   io_pipe_phv_in_data_250,
  input  [7:0]   io_pipe_phv_in_data_251,
  input  [7:0]   io_pipe_phv_in_data_252,
  input  [7:0]   io_pipe_phv_in_data_253,
  input  [7:0]   io_pipe_phv_in_data_254,
  input  [7:0]   io_pipe_phv_in_data_255,
  input  [3:0]   io_pipe_phv_in_next_processor_id,
  input          io_pipe_phv_in_next_config_id,
  input          io_pipe_phv_in_is_valid_processor,
  output [7:0]   io_pipe_phv_out_data_0,
  output [7:0]   io_pipe_phv_out_data_1,
  output [7:0]   io_pipe_phv_out_data_2,
  output [7:0]   io_pipe_phv_out_data_3,
  output [7:0]   io_pipe_phv_out_data_4,
  output [7:0]   io_pipe_phv_out_data_5,
  output [7:0]   io_pipe_phv_out_data_6,
  output [7:0]   io_pipe_phv_out_data_7,
  output [7:0]   io_pipe_phv_out_data_8,
  output [7:0]   io_pipe_phv_out_data_9,
  output [7:0]   io_pipe_phv_out_data_10,
  output [7:0]   io_pipe_phv_out_data_11,
  output [7:0]   io_pipe_phv_out_data_12,
  output [7:0]   io_pipe_phv_out_data_13,
  output [7:0]   io_pipe_phv_out_data_14,
  output [7:0]   io_pipe_phv_out_data_15,
  output [7:0]   io_pipe_phv_out_data_16,
  output [7:0]   io_pipe_phv_out_data_17,
  output [7:0]   io_pipe_phv_out_data_18,
  output [7:0]   io_pipe_phv_out_data_19,
  output [7:0]   io_pipe_phv_out_data_20,
  output [7:0]   io_pipe_phv_out_data_21,
  output [7:0]   io_pipe_phv_out_data_22,
  output [7:0]   io_pipe_phv_out_data_23,
  output [7:0]   io_pipe_phv_out_data_24,
  output [7:0]   io_pipe_phv_out_data_25,
  output [7:0]   io_pipe_phv_out_data_26,
  output [7:0]   io_pipe_phv_out_data_27,
  output [7:0]   io_pipe_phv_out_data_28,
  output [7:0]   io_pipe_phv_out_data_29,
  output [7:0]   io_pipe_phv_out_data_30,
  output [7:0]   io_pipe_phv_out_data_31,
  output [7:0]   io_pipe_phv_out_data_32,
  output [7:0]   io_pipe_phv_out_data_33,
  output [7:0]   io_pipe_phv_out_data_34,
  output [7:0]   io_pipe_phv_out_data_35,
  output [7:0]   io_pipe_phv_out_data_36,
  output [7:0]   io_pipe_phv_out_data_37,
  output [7:0]   io_pipe_phv_out_data_38,
  output [7:0]   io_pipe_phv_out_data_39,
  output [7:0]   io_pipe_phv_out_data_40,
  output [7:0]   io_pipe_phv_out_data_41,
  output [7:0]   io_pipe_phv_out_data_42,
  output [7:0]   io_pipe_phv_out_data_43,
  output [7:0]   io_pipe_phv_out_data_44,
  output [7:0]   io_pipe_phv_out_data_45,
  output [7:0]   io_pipe_phv_out_data_46,
  output [7:0]   io_pipe_phv_out_data_47,
  output [7:0]   io_pipe_phv_out_data_48,
  output [7:0]   io_pipe_phv_out_data_49,
  output [7:0]   io_pipe_phv_out_data_50,
  output [7:0]   io_pipe_phv_out_data_51,
  output [7:0]   io_pipe_phv_out_data_52,
  output [7:0]   io_pipe_phv_out_data_53,
  output [7:0]   io_pipe_phv_out_data_54,
  output [7:0]   io_pipe_phv_out_data_55,
  output [7:0]   io_pipe_phv_out_data_56,
  output [7:0]   io_pipe_phv_out_data_57,
  output [7:0]   io_pipe_phv_out_data_58,
  output [7:0]   io_pipe_phv_out_data_59,
  output [7:0]   io_pipe_phv_out_data_60,
  output [7:0]   io_pipe_phv_out_data_61,
  output [7:0]   io_pipe_phv_out_data_62,
  output [7:0]   io_pipe_phv_out_data_63,
  output [7:0]   io_pipe_phv_out_data_64,
  output [7:0]   io_pipe_phv_out_data_65,
  output [7:0]   io_pipe_phv_out_data_66,
  output [7:0]   io_pipe_phv_out_data_67,
  output [7:0]   io_pipe_phv_out_data_68,
  output [7:0]   io_pipe_phv_out_data_69,
  output [7:0]   io_pipe_phv_out_data_70,
  output [7:0]   io_pipe_phv_out_data_71,
  output [7:0]   io_pipe_phv_out_data_72,
  output [7:0]   io_pipe_phv_out_data_73,
  output [7:0]   io_pipe_phv_out_data_74,
  output [7:0]   io_pipe_phv_out_data_75,
  output [7:0]   io_pipe_phv_out_data_76,
  output [7:0]   io_pipe_phv_out_data_77,
  output [7:0]   io_pipe_phv_out_data_78,
  output [7:0]   io_pipe_phv_out_data_79,
  output [7:0]   io_pipe_phv_out_data_80,
  output [7:0]   io_pipe_phv_out_data_81,
  output [7:0]   io_pipe_phv_out_data_82,
  output [7:0]   io_pipe_phv_out_data_83,
  output [7:0]   io_pipe_phv_out_data_84,
  output [7:0]   io_pipe_phv_out_data_85,
  output [7:0]   io_pipe_phv_out_data_86,
  output [7:0]   io_pipe_phv_out_data_87,
  output [7:0]   io_pipe_phv_out_data_88,
  output [7:0]   io_pipe_phv_out_data_89,
  output [7:0]   io_pipe_phv_out_data_90,
  output [7:0]   io_pipe_phv_out_data_91,
  output [7:0]   io_pipe_phv_out_data_92,
  output [7:0]   io_pipe_phv_out_data_93,
  output [7:0]   io_pipe_phv_out_data_94,
  output [7:0]   io_pipe_phv_out_data_95,
  output [7:0]   io_pipe_phv_out_data_96,
  output [7:0]   io_pipe_phv_out_data_97,
  output [7:0]   io_pipe_phv_out_data_98,
  output [7:0]   io_pipe_phv_out_data_99,
  output [7:0]   io_pipe_phv_out_data_100,
  output [7:0]   io_pipe_phv_out_data_101,
  output [7:0]   io_pipe_phv_out_data_102,
  output [7:0]   io_pipe_phv_out_data_103,
  output [7:0]   io_pipe_phv_out_data_104,
  output [7:0]   io_pipe_phv_out_data_105,
  output [7:0]   io_pipe_phv_out_data_106,
  output [7:0]   io_pipe_phv_out_data_107,
  output [7:0]   io_pipe_phv_out_data_108,
  output [7:0]   io_pipe_phv_out_data_109,
  output [7:0]   io_pipe_phv_out_data_110,
  output [7:0]   io_pipe_phv_out_data_111,
  output [7:0]   io_pipe_phv_out_data_112,
  output [7:0]   io_pipe_phv_out_data_113,
  output [7:0]   io_pipe_phv_out_data_114,
  output [7:0]   io_pipe_phv_out_data_115,
  output [7:0]   io_pipe_phv_out_data_116,
  output [7:0]   io_pipe_phv_out_data_117,
  output [7:0]   io_pipe_phv_out_data_118,
  output [7:0]   io_pipe_phv_out_data_119,
  output [7:0]   io_pipe_phv_out_data_120,
  output [7:0]   io_pipe_phv_out_data_121,
  output [7:0]   io_pipe_phv_out_data_122,
  output [7:0]   io_pipe_phv_out_data_123,
  output [7:0]   io_pipe_phv_out_data_124,
  output [7:0]   io_pipe_phv_out_data_125,
  output [7:0]   io_pipe_phv_out_data_126,
  output [7:0]   io_pipe_phv_out_data_127,
  output [7:0]   io_pipe_phv_out_data_128,
  output [7:0]   io_pipe_phv_out_data_129,
  output [7:0]   io_pipe_phv_out_data_130,
  output [7:0]   io_pipe_phv_out_data_131,
  output [7:0]   io_pipe_phv_out_data_132,
  output [7:0]   io_pipe_phv_out_data_133,
  output [7:0]   io_pipe_phv_out_data_134,
  output [7:0]   io_pipe_phv_out_data_135,
  output [7:0]   io_pipe_phv_out_data_136,
  output [7:0]   io_pipe_phv_out_data_137,
  output [7:0]   io_pipe_phv_out_data_138,
  output [7:0]   io_pipe_phv_out_data_139,
  output [7:0]   io_pipe_phv_out_data_140,
  output [7:0]   io_pipe_phv_out_data_141,
  output [7:0]   io_pipe_phv_out_data_142,
  output [7:0]   io_pipe_phv_out_data_143,
  output [7:0]   io_pipe_phv_out_data_144,
  output [7:0]   io_pipe_phv_out_data_145,
  output [7:0]   io_pipe_phv_out_data_146,
  output [7:0]   io_pipe_phv_out_data_147,
  output [7:0]   io_pipe_phv_out_data_148,
  output [7:0]   io_pipe_phv_out_data_149,
  output [7:0]   io_pipe_phv_out_data_150,
  output [7:0]   io_pipe_phv_out_data_151,
  output [7:0]   io_pipe_phv_out_data_152,
  output [7:0]   io_pipe_phv_out_data_153,
  output [7:0]   io_pipe_phv_out_data_154,
  output [7:0]   io_pipe_phv_out_data_155,
  output [7:0]   io_pipe_phv_out_data_156,
  output [7:0]   io_pipe_phv_out_data_157,
  output [7:0]   io_pipe_phv_out_data_158,
  output [7:0]   io_pipe_phv_out_data_159,
  output [7:0]   io_pipe_phv_out_data_160,
  output [7:0]   io_pipe_phv_out_data_161,
  output [7:0]   io_pipe_phv_out_data_162,
  output [7:0]   io_pipe_phv_out_data_163,
  output [7:0]   io_pipe_phv_out_data_164,
  output [7:0]   io_pipe_phv_out_data_165,
  output [7:0]   io_pipe_phv_out_data_166,
  output [7:0]   io_pipe_phv_out_data_167,
  output [7:0]   io_pipe_phv_out_data_168,
  output [7:0]   io_pipe_phv_out_data_169,
  output [7:0]   io_pipe_phv_out_data_170,
  output [7:0]   io_pipe_phv_out_data_171,
  output [7:0]   io_pipe_phv_out_data_172,
  output [7:0]   io_pipe_phv_out_data_173,
  output [7:0]   io_pipe_phv_out_data_174,
  output [7:0]   io_pipe_phv_out_data_175,
  output [7:0]   io_pipe_phv_out_data_176,
  output [7:0]   io_pipe_phv_out_data_177,
  output [7:0]   io_pipe_phv_out_data_178,
  output [7:0]   io_pipe_phv_out_data_179,
  output [7:0]   io_pipe_phv_out_data_180,
  output [7:0]   io_pipe_phv_out_data_181,
  output [7:0]   io_pipe_phv_out_data_182,
  output [7:0]   io_pipe_phv_out_data_183,
  output [7:0]   io_pipe_phv_out_data_184,
  output [7:0]   io_pipe_phv_out_data_185,
  output [7:0]   io_pipe_phv_out_data_186,
  output [7:0]   io_pipe_phv_out_data_187,
  output [7:0]   io_pipe_phv_out_data_188,
  output [7:0]   io_pipe_phv_out_data_189,
  output [7:0]   io_pipe_phv_out_data_190,
  output [7:0]   io_pipe_phv_out_data_191,
  output [7:0]   io_pipe_phv_out_data_192,
  output [7:0]   io_pipe_phv_out_data_193,
  output [7:0]   io_pipe_phv_out_data_194,
  output [7:0]   io_pipe_phv_out_data_195,
  output [7:0]   io_pipe_phv_out_data_196,
  output [7:0]   io_pipe_phv_out_data_197,
  output [7:0]   io_pipe_phv_out_data_198,
  output [7:0]   io_pipe_phv_out_data_199,
  output [7:0]   io_pipe_phv_out_data_200,
  output [7:0]   io_pipe_phv_out_data_201,
  output [7:0]   io_pipe_phv_out_data_202,
  output [7:0]   io_pipe_phv_out_data_203,
  output [7:0]   io_pipe_phv_out_data_204,
  output [7:0]   io_pipe_phv_out_data_205,
  output [7:0]   io_pipe_phv_out_data_206,
  output [7:0]   io_pipe_phv_out_data_207,
  output [7:0]   io_pipe_phv_out_data_208,
  output [7:0]   io_pipe_phv_out_data_209,
  output [7:0]   io_pipe_phv_out_data_210,
  output [7:0]   io_pipe_phv_out_data_211,
  output [7:0]   io_pipe_phv_out_data_212,
  output [7:0]   io_pipe_phv_out_data_213,
  output [7:0]   io_pipe_phv_out_data_214,
  output [7:0]   io_pipe_phv_out_data_215,
  output [7:0]   io_pipe_phv_out_data_216,
  output [7:0]   io_pipe_phv_out_data_217,
  output [7:0]   io_pipe_phv_out_data_218,
  output [7:0]   io_pipe_phv_out_data_219,
  output [7:0]   io_pipe_phv_out_data_220,
  output [7:0]   io_pipe_phv_out_data_221,
  output [7:0]   io_pipe_phv_out_data_222,
  output [7:0]   io_pipe_phv_out_data_223,
  output [7:0]   io_pipe_phv_out_data_224,
  output [7:0]   io_pipe_phv_out_data_225,
  output [7:0]   io_pipe_phv_out_data_226,
  output [7:0]   io_pipe_phv_out_data_227,
  output [7:0]   io_pipe_phv_out_data_228,
  output [7:0]   io_pipe_phv_out_data_229,
  output [7:0]   io_pipe_phv_out_data_230,
  output [7:0]   io_pipe_phv_out_data_231,
  output [7:0]   io_pipe_phv_out_data_232,
  output [7:0]   io_pipe_phv_out_data_233,
  output [7:0]   io_pipe_phv_out_data_234,
  output [7:0]   io_pipe_phv_out_data_235,
  output [7:0]   io_pipe_phv_out_data_236,
  output [7:0]   io_pipe_phv_out_data_237,
  output [7:0]   io_pipe_phv_out_data_238,
  output [7:0]   io_pipe_phv_out_data_239,
  output [7:0]   io_pipe_phv_out_data_240,
  output [7:0]   io_pipe_phv_out_data_241,
  output [7:0]   io_pipe_phv_out_data_242,
  output [7:0]   io_pipe_phv_out_data_243,
  output [7:0]   io_pipe_phv_out_data_244,
  output [7:0]   io_pipe_phv_out_data_245,
  output [7:0]   io_pipe_phv_out_data_246,
  output [7:0]   io_pipe_phv_out_data_247,
  output [7:0]   io_pipe_phv_out_data_248,
  output [7:0]   io_pipe_phv_out_data_249,
  output [7:0]   io_pipe_phv_out_data_250,
  output [7:0]   io_pipe_phv_out_data_251,
  output [7:0]   io_pipe_phv_out_data_252,
  output [7:0]   io_pipe_phv_out_data_253,
  output [7:0]   io_pipe_phv_out_data_254,
  output [7:0]   io_pipe_phv_out_data_255,
  output [3:0]   io_pipe_phv_out_next_processor_id,
  output         io_pipe_phv_out_next_config_id,
  output         io_pipe_phv_out_is_valid_processor,
  input  [1:0]   io_key_config_0_field_config_0,
  input  [1:0]   io_key_config_0_field_config_1,
  input  [1:0]   io_key_config_0_field_config_2,
  input  [1:0]   io_key_config_0_field_config_3,
  input  [1:0]   io_key_config_0_field_config_4,
  input  [1:0]   io_key_config_0_field_config_5,
  input          io_key_config_0_field_mask_0_0,
  input          io_key_config_0_field_mask_0_1,
  input          io_key_config_0_field_mask_0_2,
  input          io_key_config_0_field_mask_0_3,
  input          io_key_config_0_field_mask_1_0,
  input          io_key_config_0_field_mask_1_1,
  input          io_key_config_0_field_mask_1_2,
  input          io_key_config_0_field_mask_1_3,
  input          io_key_config_0_field_mask_2_0,
  input          io_key_config_0_field_mask_2_1,
  input          io_key_config_0_field_mask_2_2,
  input          io_key_config_0_field_mask_2_3,
  input          io_key_config_0_field_mask_3_0,
  input          io_key_config_0_field_mask_3_1,
  input          io_key_config_0_field_mask_3_2,
  input          io_key_config_0_field_mask_3_3,
  input          io_key_config_0_field_mask_4_0,
  input          io_key_config_0_field_mask_4_1,
  input          io_key_config_0_field_mask_4_2,
  input          io_key_config_0_field_mask_4_3,
  input          io_key_config_0_field_mask_5_0,
  input          io_key_config_0_field_mask_5_1,
  input          io_key_config_0_field_mask_5_2,
  input          io_key_config_0_field_mask_5_3,
  input  [7:0]   io_key_config_0_field_id_0_0,
  input  [7:0]   io_key_config_0_field_id_0_1,
  input  [7:0]   io_key_config_0_field_id_0_2,
  input  [7:0]   io_key_config_0_field_id_0_3,
  input  [7:0]   io_key_config_0_field_id_1_0,
  input  [7:0]   io_key_config_0_field_id_1_1,
  input  [7:0]   io_key_config_0_field_id_1_2,
  input  [7:0]   io_key_config_0_field_id_1_3,
  input  [7:0]   io_key_config_0_field_id_2_0,
  input  [7:0]   io_key_config_0_field_id_2_1,
  input  [7:0]   io_key_config_0_field_id_2_2,
  input  [7:0]   io_key_config_0_field_id_2_3,
  input  [7:0]   io_key_config_0_field_id_3_0,
  input  [7:0]   io_key_config_0_field_id_3_1,
  input  [7:0]   io_key_config_0_field_id_3_2,
  input  [7:0]   io_key_config_0_field_id_3_3,
  input  [7:0]   io_key_config_0_field_id_4_0,
  input  [7:0]   io_key_config_0_field_id_4_1,
  input  [7:0]   io_key_config_0_field_id_4_2,
  input  [7:0]   io_key_config_0_field_id_4_3,
  input  [7:0]   io_key_config_0_field_id_5_0,
  input  [7:0]   io_key_config_0_field_id_5_1,
  input  [7:0]   io_key_config_0_field_id_5_2,
  input  [7:0]   io_key_config_0_field_id_5_3,
  input  [1:0]   io_key_config_1_field_config_0,
  input  [1:0]   io_key_config_1_field_config_1,
  input  [1:0]   io_key_config_1_field_config_2,
  input  [1:0]   io_key_config_1_field_config_3,
  input  [1:0]   io_key_config_1_field_config_4,
  input  [1:0]   io_key_config_1_field_config_5,
  input          io_key_config_1_field_mask_0_0,
  input          io_key_config_1_field_mask_0_1,
  input          io_key_config_1_field_mask_0_2,
  input          io_key_config_1_field_mask_0_3,
  input          io_key_config_1_field_mask_1_0,
  input          io_key_config_1_field_mask_1_1,
  input          io_key_config_1_field_mask_1_2,
  input          io_key_config_1_field_mask_1_3,
  input          io_key_config_1_field_mask_2_0,
  input          io_key_config_1_field_mask_2_1,
  input          io_key_config_1_field_mask_2_2,
  input          io_key_config_1_field_mask_2_3,
  input          io_key_config_1_field_mask_3_0,
  input          io_key_config_1_field_mask_3_1,
  input          io_key_config_1_field_mask_3_2,
  input          io_key_config_1_field_mask_3_3,
  input          io_key_config_1_field_mask_4_0,
  input          io_key_config_1_field_mask_4_1,
  input          io_key_config_1_field_mask_4_2,
  input          io_key_config_1_field_mask_4_3,
  input          io_key_config_1_field_mask_5_0,
  input          io_key_config_1_field_mask_5_1,
  input          io_key_config_1_field_mask_5_2,
  input          io_key_config_1_field_mask_5_3,
  input  [7:0]   io_key_config_1_field_id_0_0,
  input  [7:0]   io_key_config_1_field_id_0_1,
  input  [7:0]   io_key_config_1_field_id_0_2,
  input  [7:0]   io_key_config_1_field_id_0_3,
  input  [7:0]   io_key_config_1_field_id_1_0,
  input  [7:0]   io_key_config_1_field_id_1_1,
  input  [7:0]   io_key_config_1_field_id_1_2,
  input  [7:0]   io_key_config_1_field_id_1_3,
  input  [7:0]   io_key_config_1_field_id_2_0,
  input  [7:0]   io_key_config_1_field_id_2_1,
  input  [7:0]   io_key_config_1_field_id_2_2,
  input  [7:0]   io_key_config_1_field_id_2_3,
  input  [7:0]   io_key_config_1_field_id_3_0,
  input  [7:0]   io_key_config_1_field_id_3_1,
  input  [7:0]   io_key_config_1_field_id_3_2,
  input  [7:0]   io_key_config_1_field_id_3_3,
  input  [7:0]   io_key_config_1_field_id_4_0,
  input  [7:0]   io_key_config_1_field_id_4_1,
  input  [7:0]   io_key_config_1_field_id_4_2,
  input  [7:0]   io_key_config_1_field_id_4_3,
  input  [7:0]   io_key_config_1_field_id_5_0,
  input  [7:0]   io_key_config_1_field_id_5_1,
  input  [7:0]   io_key_config_1_field_id_5_2,
  input  [7:0]   io_key_config_1_field_id_5_3,
  output [191:0] io_match_key
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_1; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_2; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_3; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_4; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_5; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_6; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_7; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_8; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_9; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_10; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_11; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_12; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_13; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_14; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_15; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_16; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_17; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_18; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_19; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_20; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_21; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_22; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_23; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_24; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_25; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_26; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_27; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_28; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_29; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_30; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_31; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_32; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_33; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_34; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_35; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_36; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_37; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_38; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_39; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_40; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_41; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_42; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_43; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_44; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_45; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_46; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_47; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_48; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_49; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_50; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_51; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_52; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_53; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_54; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_55; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_56; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_57; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_58; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_59; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_60; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_61; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_62; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_63; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_64; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_65; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_66; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_67; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_68; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_69; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_70; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_71; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_72; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_73; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_74; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_75; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_76; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_77; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_78; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_79; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_80; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_81; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_82; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_83; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_84; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_85; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_86; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_87; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_88; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_89; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_90; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_91; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_92; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_93; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_94; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_95; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_96; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_97; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_98; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_99; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_100; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_101; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_102; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_103; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_104; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_105; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_106; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_107; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_108; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_109; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_110; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_111; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_112; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_113; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_114; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_115; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_116; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_117; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_118; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_119; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_120; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_121; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_122; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_123; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_124; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_125; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_126; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_127; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_128; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_129; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_130; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_131; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_132; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_133; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_134; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_135; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_136; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_137; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_138; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_139; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_140; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_141; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_142; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_143; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_144; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_145; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_146; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_147; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_148; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_149; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_150; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_151; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_152; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_153; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_154; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_155; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_156; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_157; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_158; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_159; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_160; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_161; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_162; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_163; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_164; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_165; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_166; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_167; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_168; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_169; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_170; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_171; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_172; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_173; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_174; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_175; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_176; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_177; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_178; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_179; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_180; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_181; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_182; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_183; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_184; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_185; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_186; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_187; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_188; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_189; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_190; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_191; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_192; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_193; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_194; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_195; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_196; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_197; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_198; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_199; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_200; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_201; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_202; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_203; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_204; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_205; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_206; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_207; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_208; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_209; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_210; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_211; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_212; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_213; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_214; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_215; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_216; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_217; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_218; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_219; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_220; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_221; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_222; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_223; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_224; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_225; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_226; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_227; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_228; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_229; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_230; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_231; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_232; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_233; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_234; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_235; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_236; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_237; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_238; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_239; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_240; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_241; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_242; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_243; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_244; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_245; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_246; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_247; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_248; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_249; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_250; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_251; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_252; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_253; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_254; // @[matcher_pisa.scala 110:22]
  reg [7:0] phv_data_255; // @[matcher_pisa.scala 110:22]
  reg [3:0] phv_next_processor_id; // @[matcher_pisa.scala 110:22]
  reg  phv_next_config_id; // @[matcher_pisa.scala 110:22]
  reg  phv_is_valid_processor; // @[matcher_pisa.scala 110:22]
  wire [1:0] _GEN_56 = phv_next_config_id ? io_key_config_1_field_config_0 : io_key_config_0_field_config_0; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [1:0] _GEN_57 = phv_next_config_id ? io_key_config_1_field_config_1 : io_key_config_0_field_config_1; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [1:0] _GEN_58 = phv_next_config_id ? io_key_config_1_field_config_2 : io_key_config_0_field_config_2; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [1:0] _GEN_59 = phv_next_config_id ? io_key_config_1_field_config_3 : io_key_config_0_field_config_3; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [1:0] _GEN_60 = phv_next_config_id ? io_key_config_1_field_config_4 : io_key_config_0_field_config_4; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [1:0] _GEN_61 = phv_next_config_id ? io_key_config_1_field_config_5 : io_key_config_0_field_config_5; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_62 = phv_next_config_id ? io_key_config_1_field_mask_0_0 : io_key_config_0_field_mask_0_0; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_63 = phv_next_config_id ? io_key_config_1_field_mask_0_1 : io_key_config_0_field_mask_0_1; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_64 = phv_next_config_id ? io_key_config_1_field_mask_0_2 : io_key_config_0_field_mask_0_2; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_65 = phv_next_config_id ? io_key_config_1_field_mask_0_3 : io_key_config_0_field_mask_0_3; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_66 = phv_next_config_id ? io_key_config_1_field_mask_1_0 : io_key_config_0_field_mask_1_0; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_67 = phv_next_config_id ? io_key_config_1_field_mask_1_1 : io_key_config_0_field_mask_1_1; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_68 = phv_next_config_id ? io_key_config_1_field_mask_1_2 : io_key_config_0_field_mask_1_2; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_69 = phv_next_config_id ? io_key_config_1_field_mask_1_3 : io_key_config_0_field_mask_1_3; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_70 = phv_next_config_id ? io_key_config_1_field_mask_2_0 : io_key_config_0_field_mask_2_0; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_71 = phv_next_config_id ? io_key_config_1_field_mask_2_1 : io_key_config_0_field_mask_2_1; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_72 = phv_next_config_id ? io_key_config_1_field_mask_2_2 : io_key_config_0_field_mask_2_2; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_73 = phv_next_config_id ? io_key_config_1_field_mask_2_3 : io_key_config_0_field_mask_2_3; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_74 = phv_next_config_id ? io_key_config_1_field_mask_3_0 : io_key_config_0_field_mask_3_0; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_75 = phv_next_config_id ? io_key_config_1_field_mask_3_1 : io_key_config_0_field_mask_3_1; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_76 = phv_next_config_id ? io_key_config_1_field_mask_3_2 : io_key_config_0_field_mask_3_2; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_77 = phv_next_config_id ? io_key_config_1_field_mask_3_3 : io_key_config_0_field_mask_3_3; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_78 = phv_next_config_id ? io_key_config_1_field_mask_4_0 : io_key_config_0_field_mask_4_0; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_79 = phv_next_config_id ? io_key_config_1_field_mask_4_1 : io_key_config_0_field_mask_4_1; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_80 = phv_next_config_id ? io_key_config_1_field_mask_4_2 : io_key_config_0_field_mask_4_2; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_81 = phv_next_config_id ? io_key_config_1_field_mask_4_3 : io_key_config_0_field_mask_4_3; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_82 = phv_next_config_id ? io_key_config_1_field_mask_5_0 : io_key_config_0_field_mask_5_0; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_83 = phv_next_config_id ? io_key_config_1_field_mask_5_1 : io_key_config_0_field_mask_5_1; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_84 = phv_next_config_id ? io_key_config_1_field_mask_5_2 : io_key_config_0_field_mask_5_2; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire  _GEN_85 = phv_next_config_id ? io_key_config_1_field_mask_5_3 : io_key_config_0_field_mask_5_3; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_86 = phv_next_config_id ? io_key_config_1_field_id_0_0 : io_key_config_0_field_id_0_0; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_87 = phv_next_config_id ? io_key_config_1_field_id_0_1 : io_key_config_0_field_id_0_1; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_88 = phv_next_config_id ? io_key_config_1_field_id_0_2 : io_key_config_0_field_id_0_2; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_89 = phv_next_config_id ? io_key_config_1_field_id_0_3 : io_key_config_0_field_id_0_3; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_90 = phv_next_config_id ? io_key_config_1_field_id_1_0 : io_key_config_0_field_id_1_0; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_91 = phv_next_config_id ? io_key_config_1_field_id_1_1 : io_key_config_0_field_id_1_1; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_92 = phv_next_config_id ? io_key_config_1_field_id_1_2 : io_key_config_0_field_id_1_2; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_93 = phv_next_config_id ? io_key_config_1_field_id_1_3 : io_key_config_0_field_id_1_3; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_94 = phv_next_config_id ? io_key_config_1_field_id_2_0 : io_key_config_0_field_id_2_0; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_95 = phv_next_config_id ? io_key_config_1_field_id_2_1 : io_key_config_0_field_id_2_1; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_96 = phv_next_config_id ? io_key_config_1_field_id_2_2 : io_key_config_0_field_id_2_2; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_97 = phv_next_config_id ? io_key_config_1_field_id_2_3 : io_key_config_0_field_id_2_3; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_98 = phv_next_config_id ? io_key_config_1_field_id_3_0 : io_key_config_0_field_id_3_0; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_99 = phv_next_config_id ? io_key_config_1_field_id_3_1 : io_key_config_0_field_id_3_1; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_100 = phv_next_config_id ? io_key_config_1_field_id_3_2 : io_key_config_0_field_id_3_2; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_101 = phv_next_config_id ? io_key_config_1_field_id_3_3 : io_key_config_0_field_id_3_3; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_102 = phv_next_config_id ? io_key_config_1_field_id_4_0 : io_key_config_0_field_id_4_0; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_103 = phv_next_config_id ? io_key_config_1_field_id_4_1 : io_key_config_0_field_id_4_1; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_104 = phv_next_config_id ? io_key_config_1_field_id_4_2 : io_key_config_0_field_id_4_2; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_105 = phv_next_config_id ? io_key_config_1_field_id_4_3 : io_key_config_0_field_id_4_3; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_106 = phv_next_config_id ? io_key_config_1_field_id_5_0 : io_key_config_0_field_id_5_0; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_107 = phv_next_config_id ? io_key_config_1_field_id_5_1 : io_key_config_0_field_id_5_1; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_108 = phv_next_config_id ? io_key_config_1_field_id_5_2 : io_key_config_0_field_id_5_2; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_109 = phv_next_config_id ? io_key_config_1_field_id_5_3 : io_key_config_0_field_id_5_3; // @[matcher_pisa.scala 123:36 matcher_pisa.scala 123:36]
  wire [7:0] _GEN_110 = 8'h0 == _GEN_86 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_111 = 8'h1 == _GEN_86 ? phv_data_1 : _GEN_110; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_112 = 8'h2 == _GEN_86 ? phv_data_2 : _GEN_111; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_113 = 8'h3 == _GEN_86 ? phv_data_3 : _GEN_112; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_114 = 8'h4 == _GEN_86 ? phv_data_4 : _GEN_113; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_115 = 8'h5 == _GEN_86 ? phv_data_5 : _GEN_114; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_116 = 8'h6 == _GEN_86 ? phv_data_6 : _GEN_115; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_117 = 8'h7 == _GEN_86 ? phv_data_7 : _GEN_116; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_118 = 8'h8 == _GEN_86 ? phv_data_8 : _GEN_117; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_119 = 8'h9 == _GEN_86 ? phv_data_9 : _GEN_118; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_120 = 8'ha == _GEN_86 ? phv_data_10 : _GEN_119; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_121 = 8'hb == _GEN_86 ? phv_data_11 : _GEN_120; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_122 = 8'hc == _GEN_86 ? phv_data_12 : _GEN_121; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_123 = 8'hd == _GEN_86 ? phv_data_13 : _GEN_122; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_124 = 8'he == _GEN_86 ? phv_data_14 : _GEN_123; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_125 = 8'hf == _GEN_86 ? phv_data_15 : _GEN_124; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_126 = 8'h10 == _GEN_86 ? phv_data_16 : _GEN_125; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_127 = 8'h11 == _GEN_86 ? phv_data_17 : _GEN_126; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_128 = 8'h12 == _GEN_86 ? phv_data_18 : _GEN_127; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_129 = 8'h13 == _GEN_86 ? phv_data_19 : _GEN_128; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_130 = 8'h14 == _GEN_86 ? phv_data_20 : _GEN_129; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_131 = 8'h15 == _GEN_86 ? phv_data_21 : _GEN_130; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_132 = 8'h16 == _GEN_86 ? phv_data_22 : _GEN_131; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_133 = 8'h17 == _GEN_86 ? phv_data_23 : _GEN_132; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_134 = 8'h18 == _GEN_86 ? phv_data_24 : _GEN_133; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_135 = 8'h19 == _GEN_86 ? phv_data_25 : _GEN_134; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_136 = 8'h1a == _GEN_86 ? phv_data_26 : _GEN_135; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_137 = 8'h1b == _GEN_86 ? phv_data_27 : _GEN_136; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_138 = 8'h1c == _GEN_86 ? phv_data_28 : _GEN_137; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_139 = 8'h1d == _GEN_86 ? phv_data_29 : _GEN_138; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_140 = 8'h1e == _GEN_86 ? phv_data_30 : _GEN_139; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_141 = 8'h1f == _GEN_86 ? phv_data_31 : _GEN_140; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes__0 = _GEN_62 ? _GEN_141 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_143 = 8'h0 == _GEN_87 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_144 = 8'h1 == _GEN_87 ? phv_data_1 : _GEN_143; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_145 = 8'h2 == _GEN_87 ? phv_data_2 : _GEN_144; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_146 = 8'h3 == _GEN_87 ? phv_data_3 : _GEN_145; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_147 = 8'h4 == _GEN_87 ? phv_data_4 : _GEN_146; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_148 = 8'h5 == _GEN_87 ? phv_data_5 : _GEN_147; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_149 = 8'h6 == _GEN_87 ? phv_data_6 : _GEN_148; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_150 = 8'h7 == _GEN_87 ? phv_data_7 : _GEN_149; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_151 = 8'h8 == _GEN_87 ? phv_data_8 : _GEN_150; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_152 = 8'h9 == _GEN_87 ? phv_data_9 : _GEN_151; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_153 = 8'ha == _GEN_87 ? phv_data_10 : _GEN_152; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_154 = 8'hb == _GEN_87 ? phv_data_11 : _GEN_153; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_155 = 8'hc == _GEN_87 ? phv_data_12 : _GEN_154; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_156 = 8'hd == _GEN_87 ? phv_data_13 : _GEN_155; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_157 = 8'he == _GEN_87 ? phv_data_14 : _GEN_156; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_158 = 8'hf == _GEN_87 ? phv_data_15 : _GEN_157; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_159 = 8'h10 == _GEN_87 ? phv_data_16 : _GEN_158; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_160 = 8'h11 == _GEN_87 ? phv_data_17 : _GEN_159; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_161 = 8'h12 == _GEN_87 ? phv_data_18 : _GEN_160; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_162 = 8'h13 == _GEN_87 ? phv_data_19 : _GEN_161; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_163 = 8'h14 == _GEN_87 ? phv_data_20 : _GEN_162; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_164 = 8'h15 == _GEN_87 ? phv_data_21 : _GEN_163; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_165 = 8'h16 == _GEN_87 ? phv_data_22 : _GEN_164; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_166 = 8'h17 == _GEN_87 ? phv_data_23 : _GEN_165; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_167 = 8'h18 == _GEN_87 ? phv_data_24 : _GEN_166; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_168 = 8'h19 == _GEN_87 ? phv_data_25 : _GEN_167; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_169 = 8'h1a == _GEN_87 ? phv_data_26 : _GEN_168; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_170 = 8'h1b == _GEN_87 ? phv_data_27 : _GEN_169; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_171 = 8'h1c == _GEN_87 ? phv_data_28 : _GEN_170; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_172 = 8'h1d == _GEN_87 ? phv_data_29 : _GEN_171; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_173 = 8'h1e == _GEN_87 ? phv_data_30 : _GEN_172; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_174 = 8'h1f == _GEN_87 ? phv_data_31 : _GEN_173; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes__1 = _GEN_63 ? _GEN_174 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_176 = 8'h0 == _GEN_88 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_177 = 8'h1 == _GEN_88 ? phv_data_1 : _GEN_176; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_178 = 8'h2 == _GEN_88 ? phv_data_2 : _GEN_177; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_179 = 8'h3 == _GEN_88 ? phv_data_3 : _GEN_178; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_180 = 8'h4 == _GEN_88 ? phv_data_4 : _GEN_179; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_181 = 8'h5 == _GEN_88 ? phv_data_5 : _GEN_180; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_182 = 8'h6 == _GEN_88 ? phv_data_6 : _GEN_181; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_183 = 8'h7 == _GEN_88 ? phv_data_7 : _GEN_182; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_184 = 8'h8 == _GEN_88 ? phv_data_8 : _GEN_183; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_185 = 8'h9 == _GEN_88 ? phv_data_9 : _GEN_184; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_186 = 8'ha == _GEN_88 ? phv_data_10 : _GEN_185; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_187 = 8'hb == _GEN_88 ? phv_data_11 : _GEN_186; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_188 = 8'hc == _GEN_88 ? phv_data_12 : _GEN_187; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_189 = 8'hd == _GEN_88 ? phv_data_13 : _GEN_188; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_190 = 8'he == _GEN_88 ? phv_data_14 : _GEN_189; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_191 = 8'hf == _GEN_88 ? phv_data_15 : _GEN_190; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_192 = 8'h10 == _GEN_88 ? phv_data_16 : _GEN_191; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_193 = 8'h11 == _GEN_88 ? phv_data_17 : _GEN_192; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_194 = 8'h12 == _GEN_88 ? phv_data_18 : _GEN_193; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_195 = 8'h13 == _GEN_88 ? phv_data_19 : _GEN_194; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_196 = 8'h14 == _GEN_88 ? phv_data_20 : _GEN_195; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_197 = 8'h15 == _GEN_88 ? phv_data_21 : _GEN_196; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_198 = 8'h16 == _GEN_88 ? phv_data_22 : _GEN_197; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_199 = 8'h17 == _GEN_88 ? phv_data_23 : _GEN_198; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_200 = 8'h18 == _GEN_88 ? phv_data_24 : _GEN_199; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_201 = 8'h19 == _GEN_88 ? phv_data_25 : _GEN_200; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_202 = 8'h1a == _GEN_88 ? phv_data_26 : _GEN_201; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_203 = 8'h1b == _GEN_88 ? phv_data_27 : _GEN_202; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_204 = 8'h1c == _GEN_88 ? phv_data_28 : _GEN_203; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_205 = 8'h1d == _GEN_88 ? phv_data_29 : _GEN_204; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_206 = 8'h1e == _GEN_88 ? phv_data_30 : _GEN_205; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_207 = 8'h1f == _GEN_88 ? phv_data_31 : _GEN_206; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes__2 = _GEN_64 ? _GEN_207 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_209 = 8'h0 == _GEN_89 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_210 = 8'h1 == _GEN_89 ? phv_data_1 : _GEN_209; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_211 = 8'h2 == _GEN_89 ? phv_data_2 : _GEN_210; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_212 = 8'h3 == _GEN_89 ? phv_data_3 : _GEN_211; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_213 = 8'h4 == _GEN_89 ? phv_data_4 : _GEN_212; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_214 = 8'h5 == _GEN_89 ? phv_data_5 : _GEN_213; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_215 = 8'h6 == _GEN_89 ? phv_data_6 : _GEN_214; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_216 = 8'h7 == _GEN_89 ? phv_data_7 : _GEN_215; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_217 = 8'h8 == _GEN_89 ? phv_data_8 : _GEN_216; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_218 = 8'h9 == _GEN_89 ? phv_data_9 : _GEN_217; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_219 = 8'ha == _GEN_89 ? phv_data_10 : _GEN_218; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_220 = 8'hb == _GEN_89 ? phv_data_11 : _GEN_219; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_221 = 8'hc == _GEN_89 ? phv_data_12 : _GEN_220; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_222 = 8'hd == _GEN_89 ? phv_data_13 : _GEN_221; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_223 = 8'he == _GEN_89 ? phv_data_14 : _GEN_222; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_224 = 8'hf == _GEN_89 ? phv_data_15 : _GEN_223; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_225 = 8'h10 == _GEN_89 ? phv_data_16 : _GEN_224; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_226 = 8'h11 == _GEN_89 ? phv_data_17 : _GEN_225; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_227 = 8'h12 == _GEN_89 ? phv_data_18 : _GEN_226; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_228 = 8'h13 == _GEN_89 ? phv_data_19 : _GEN_227; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_229 = 8'h14 == _GEN_89 ? phv_data_20 : _GEN_228; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_230 = 8'h15 == _GEN_89 ? phv_data_21 : _GEN_229; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_231 = 8'h16 == _GEN_89 ? phv_data_22 : _GEN_230; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_232 = 8'h17 == _GEN_89 ? phv_data_23 : _GEN_231; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_233 = 8'h18 == _GEN_89 ? phv_data_24 : _GEN_232; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_234 = 8'h19 == _GEN_89 ? phv_data_25 : _GEN_233; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_235 = 8'h1a == _GEN_89 ? phv_data_26 : _GEN_234; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_236 = 8'h1b == _GEN_89 ? phv_data_27 : _GEN_235; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_237 = 8'h1c == _GEN_89 ? phv_data_28 : _GEN_236; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_238 = 8'h1d == _GEN_89 ? phv_data_29 : _GEN_237; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_239 = 8'h1e == _GEN_89 ? phv_data_30 : _GEN_238; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_240 = 8'h1f == _GEN_89 ? phv_data_31 : _GEN_239; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes__3 = _GEN_65 ? _GEN_240 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [31:0] _groups_0_T = {bytes__0,bytes__1,bytes__2,bytes__3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_242 = _GEN_56 == 2'h1 ? _groups_0_T : 32'h0; // @[matcher_pisa.scala 123:50 matcher_pisa.scala 137:31 matcher_pisa.scala 122:27]
  wire [15:0] _double_bytes_0_T = {phv_data_32,phv_data_33}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_243 = 8'h20 == _GEN_86 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53 matcher_pisa.scala 144:41]
  wire [15:0] _double_bytes_0_T_1 = {phv_data_34,phv_data_35}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_244 = 8'h21 == _GEN_86 ? _double_bytes_0_T_1 : _GEN_243; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_2 = {phv_data_36,phv_data_37}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_245 = 8'h22 == _GEN_86 ? _double_bytes_0_T_2 : _GEN_244; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_3 = {phv_data_38,phv_data_39}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_246 = 8'h23 == _GEN_86 ? _double_bytes_0_T_3 : _GEN_245; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_4 = {phv_data_40,phv_data_41}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_247 = 8'h24 == _GEN_86 ? _double_bytes_0_T_4 : _GEN_246; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_5 = {phv_data_42,phv_data_43}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_248 = 8'h25 == _GEN_86 ? _double_bytes_0_T_5 : _GEN_247; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_6 = {phv_data_44,phv_data_45}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_249 = 8'h26 == _GEN_86 ? _double_bytes_0_T_6 : _GEN_248; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_7 = {phv_data_46,phv_data_47}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_250 = 8'h27 == _GEN_86 ? _double_bytes_0_T_7 : _GEN_249; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_8 = {phv_data_48,phv_data_49}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_251 = 8'h28 == _GEN_86 ? _double_bytes_0_T_8 : _GEN_250; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_9 = {phv_data_50,phv_data_51}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_252 = 8'h29 == _GEN_86 ? _double_bytes_0_T_9 : _GEN_251; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_10 = {phv_data_52,phv_data_53}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_253 = 8'h2a == _GEN_86 ? _double_bytes_0_T_10 : _GEN_252; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_11 = {phv_data_54,phv_data_55}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_254 = 8'h2b == _GEN_86 ? _double_bytes_0_T_11 : _GEN_253; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_12 = {phv_data_56,phv_data_57}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_255 = 8'h2c == _GEN_86 ? _double_bytes_0_T_12 : _GEN_254; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_13 = {phv_data_58,phv_data_59}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_256 = 8'h2d == _GEN_86 ? _double_bytes_0_T_13 : _GEN_255; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_14 = {phv_data_60,phv_data_61}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_257 = 8'h2e == _GEN_86 ? _double_bytes_0_T_14 : _GEN_256; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_15 = {phv_data_62,phv_data_63}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_258 = 8'h2f == _GEN_86 ? _double_bytes_0_T_15 : _GEN_257; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_16 = {phv_data_64,phv_data_65}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_259 = 8'h30 == _GEN_86 ? _double_bytes_0_T_16 : _GEN_258; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_17 = {phv_data_66,phv_data_67}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_260 = 8'h31 == _GEN_86 ? _double_bytes_0_T_17 : _GEN_259; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_18 = {phv_data_68,phv_data_69}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_261 = 8'h32 == _GEN_86 ? _double_bytes_0_T_18 : _GEN_260; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_19 = {phv_data_70,phv_data_71}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_262 = 8'h33 == _GEN_86 ? _double_bytes_0_T_19 : _GEN_261; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_20 = {phv_data_72,phv_data_73}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_263 = 8'h34 == _GEN_86 ? _double_bytes_0_T_20 : _GEN_262; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_21 = {phv_data_74,phv_data_75}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_264 = 8'h35 == _GEN_86 ? _double_bytes_0_T_21 : _GEN_263; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_22 = {phv_data_76,phv_data_77}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_265 = 8'h36 == _GEN_86 ? _double_bytes_0_T_22 : _GEN_264; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_23 = {phv_data_78,phv_data_79}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_266 = 8'h37 == _GEN_86 ? _double_bytes_0_T_23 : _GEN_265; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_24 = {phv_data_80,phv_data_81}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_267 = 8'h38 == _GEN_86 ? _double_bytes_0_T_24 : _GEN_266; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_25 = {phv_data_82,phv_data_83}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_268 = 8'h39 == _GEN_86 ? _double_bytes_0_T_25 : _GEN_267; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_26 = {phv_data_84,phv_data_85}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_269 = 8'h3a == _GEN_86 ? _double_bytes_0_T_26 : _GEN_268; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_27 = {phv_data_86,phv_data_87}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_270 = 8'h3b == _GEN_86 ? _double_bytes_0_T_27 : _GEN_269; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_28 = {phv_data_88,phv_data_89}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_271 = 8'h3c == _GEN_86 ? _double_bytes_0_T_28 : _GEN_270; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_29 = {phv_data_90,phv_data_91}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_272 = 8'h3d == _GEN_86 ? _double_bytes_0_T_29 : _GEN_271; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_30 = {phv_data_92,phv_data_93}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_273 = 8'h3e == _GEN_86 ? _double_bytes_0_T_30 : _GEN_272; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_31 = {phv_data_94,phv_data_95}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_274 = 8'h3f == _GEN_86 ? _double_bytes_0_T_31 : _GEN_273; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_32 = {phv_data_96,phv_data_97}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_275 = 8'h40 == _GEN_86 ? _double_bytes_0_T_32 : _GEN_274; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_33 = {phv_data_98,phv_data_99}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_276 = 8'h41 == _GEN_86 ? _double_bytes_0_T_33 : _GEN_275; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_34 = {phv_data_100,phv_data_101}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_277 = 8'h42 == _GEN_86 ? _double_bytes_0_T_34 : _GEN_276; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_35 = {phv_data_102,phv_data_103}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_278 = 8'h43 == _GEN_86 ? _double_bytes_0_T_35 : _GEN_277; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_36 = {phv_data_104,phv_data_105}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_279 = 8'h44 == _GEN_86 ? _double_bytes_0_T_36 : _GEN_278; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_37 = {phv_data_106,phv_data_107}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_280 = 8'h45 == _GEN_86 ? _double_bytes_0_T_37 : _GEN_279; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_38 = {phv_data_108,phv_data_109}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_281 = 8'h46 == _GEN_86 ? _double_bytes_0_T_38 : _GEN_280; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_39 = {phv_data_110,phv_data_111}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_282 = 8'h47 == _GEN_86 ? _double_bytes_0_T_39 : _GEN_281; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_40 = {phv_data_112,phv_data_113}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_283 = 8'h48 == _GEN_86 ? _double_bytes_0_T_40 : _GEN_282; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_41 = {phv_data_114,phv_data_115}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_284 = 8'h49 == _GEN_86 ? _double_bytes_0_T_41 : _GEN_283; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_42 = {phv_data_116,phv_data_117}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_285 = 8'h4a == _GEN_86 ? _double_bytes_0_T_42 : _GEN_284; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_43 = {phv_data_118,phv_data_119}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_286 = 8'h4b == _GEN_86 ? _double_bytes_0_T_43 : _GEN_285; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_44 = {phv_data_120,phv_data_121}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_287 = 8'h4c == _GEN_86 ? _double_bytes_0_T_44 : _GEN_286; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_45 = {phv_data_122,phv_data_123}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_288 = 8'h4d == _GEN_86 ? _double_bytes_0_T_45 : _GEN_287; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_46 = {phv_data_124,phv_data_125}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_289 = 8'h4e == _GEN_86 ? _double_bytes_0_T_46 : _GEN_288; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _double_bytes_0_T_47 = {phv_data_126,phv_data_127}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_290 = 8'h4f == _GEN_86 ? _double_bytes_0_T_47 : _GEN_289; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] double_bytes__0 = _GEN_62 ? _GEN_290 : 16'h0; // @[matcher_pisa.scala 145:46 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_292 = 8'h20 == _GEN_87 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_293 = 8'h21 == _GEN_87 ? _double_bytes_0_T_1 : _GEN_292; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_294 = 8'h22 == _GEN_87 ? _double_bytes_0_T_2 : _GEN_293; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_295 = 8'h23 == _GEN_87 ? _double_bytes_0_T_3 : _GEN_294; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_296 = 8'h24 == _GEN_87 ? _double_bytes_0_T_4 : _GEN_295; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_297 = 8'h25 == _GEN_87 ? _double_bytes_0_T_5 : _GEN_296; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_298 = 8'h26 == _GEN_87 ? _double_bytes_0_T_6 : _GEN_297; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_299 = 8'h27 == _GEN_87 ? _double_bytes_0_T_7 : _GEN_298; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_300 = 8'h28 == _GEN_87 ? _double_bytes_0_T_8 : _GEN_299; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_301 = 8'h29 == _GEN_87 ? _double_bytes_0_T_9 : _GEN_300; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_302 = 8'h2a == _GEN_87 ? _double_bytes_0_T_10 : _GEN_301; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_303 = 8'h2b == _GEN_87 ? _double_bytes_0_T_11 : _GEN_302; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_304 = 8'h2c == _GEN_87 ? _double_bytes_0_T_12 : _GEN_303; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_305 = 8'h2d == _GEN_87 ? _double_bytes_0_T_13 : _GEN_304; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_306 = 8'h2e == _GEN_87 ? _double_bytes_0_T_14 : _GEN_305; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_307 = 8'h2f == _GEN_87 ? _double_bytes_0_T_15 : _GEN_306; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_308 = 8'h30 == _GEN_87 ? _double_bytes_0_T_16 : _GEN_307; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_309 = 8'h31 == _GEN_87 ? _double_bytes_0_T_17 : _GEN_308; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_310 = 8'h32 == _GEN_87 ? _double_bytes_0_T_18 : _GEN_309; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_311 = 8'h33 == _GEN_87 ? _double_bytes_0_T_19 : _GEN_310; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_312 = 8'h34 == _GEN_87 ? _double_bytes_0_T_20 : _GEN_311; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_313 = 8'h35 == _GEN_87 ? _double_bytes_0_T_21 : _GEN_312; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_314 = 8'h36 == _GEN_87 ? _double_bytes_0_T_22 : _GEN_313; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_315 = 8'h37 == _GEN_87 ? _double_bytes_0_T_23 : _GEN_314; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_316 = 8'h38 == _GEN_87 ? _double_bytes_0_T_24 : _GEN_315; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_317 = 8'h39 == _GEN_87 ? _double_bytes_0_T_25 : _GEN_316; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_318 = 8'h3a == _GEN_87 ? _double_bytes_0_T_26 : _GEN_317; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_319 = 8'h3b == _GEN_87 ? _double_bytes_0_T_27 : _GEN_318; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_320 = 8'h3c == _GEN_87 ? _double_bytes_0_T_28 : _GEN_319; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_321 = 8'h3d == _GEN_87 ? _double_bytes_0_T_29 : _GEN_320; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_322 = 8'h3e == _GEN_87 ? _double_bytes_0_T_30 : _GEN_321; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_323 = 8'h3f == _GEN_87 ? _double_bytes_0_T_31 : _GEN_322; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_324 = 8'h40 == _GEN_87 ? _double_bytes_0_T_32 : _GEN_323; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_325 = 8'h41 == _GEN_87 ? _double_bytes_0_T_33 : _GEN_324; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_326 = 8'h42 == _GEN_87 ? _double_bytes_0_T_34 : _GEN_325; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_327 = 8'h43 == _GEN_87 ? _double_bytes_0_T_35 : _GEN_326; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_328 = 8'h44 == _GEN_87 ? _double_bytes_0_T_36 : _GEN_327; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_329 = 8'h45 == _GEN_87 ? _double_bytes_0_T_37 : _GEN_328; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_330 = 8'h46 == _GEN_87 ? _double_bytes_0_T_38 : _GEN_329; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_331 = 8'h47 == _GEN_87 ? _double_bytes_0_T_39 : _GEN_330; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_332 = 8'h48 == _GEN_87 ? _double_bytes_0_T_40 : _GEN_331; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_333 = 8'h49 == _GEN_87 ? _double_bytes_0_T_41 : _GEN_332; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_334 = 8'h4a == _GEN_87 ? _double_bytes_0_T_42 : _GEN_333; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_335 = 8'h4b == _GEN_87 ? _double_bytes_0_T_43 : _GEN_334; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_336 = 8'h4c == _GEN_87 ? _double_bytes_0_T_44 : _GEN_335; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_337 = 8'h4d == _GEN_87 ? _double_bytes_0_T_45 : _GEN_336; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_338 = 8'h4e == _GEN_87 ? _double_bytes_0_T_46 : _GEN_337; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_339 = 8'h4f == _GEN_87 ? _double_bytes_0_T_47 : _GEN_338; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] double_bytes__1 = _GEN_63 ? _GEN_339 : 16'h0; // @[matcher_pisa.scala 145:46 matcher_pisa.scala 144:41]
  wire [31:0] _groups_0_T_1 = {double_bytes__0,double_bytes__1}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_341 = _GEN_56 == 2'h2 ? _groups_0_T_1 : _GEN_242; // @[matcher_pisa.scala 139:50 matcher_pisa.scala 153:31]
  wire [31:0] _groups_0_T_2 = {phv_data_128,phv_data_129,phv_data_130,phv_data_131}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_342 = 8'h50 == _GEN_86 ? _groups_0_T_2 : 32'h0; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39 matcher_pisa.scala 158:31]
  wire [31:0] _groups_0_T_3 = {phv_data_132,phv_data_133,phv_data_134,phv_data_135}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_343 = 8'h51 == _GEN_86 ? _groups_0_T_3 : _GEN_342; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_4 = {phv_data_136,phv_data_137,phv_data_138,phv_data_139}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_344 = 8'h52 == _GEN_86 ? _groups_0_T_4 : _GEN_343; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_5 = {phv_data_140,phv_data_141,phv_data_142,phv_data_143}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_345 = 8'h53 == _GEN_86 ? _groups_0_T_5 : _GEN_344; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_6 = {phv_data_144,phv_data_145,phv_data_146,phv_data_147}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_346 = 8'h54 == _GEN_86 ? _groups_0_T_6 : _GEN_345; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_7 = {phv_data_148,phv_data_149,phv_data_150,phv_data_151}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_347 = 8'h55 == _GEN_86 ? _groups_0_T_7 : _GEN_346; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_8 = {phv_data_152,phv_data_153,phv_data_154,phv_data_155}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_348 = 8'h56 == _GEN_86 ? _groups_0_T_8 : _GEN_347; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_9 = {phv_data_156,phv_data_157,phv_data_158,phv_data_159}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_349 = 8'h57 == _GEN_86 ? _groups_0_T_9 : _GEN_348; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_10 = {phv_data_160,phv_data_161,phv_data_162,phv_data_163}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_350 = 8'h58 == _GEN_86 ? _groups_0_T_10 : _GEN_349; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_11 = {phv_data_164,phv_data_165,phv_data_166,phv_data_167}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_351 = 8'h59 == _GEN_86 ? _groups_0_T_11 : _GEN_350; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_12 = {phv_data_168,phv_data_169,phv_data_170,phv_data_171}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_352 = 8'h5a == _GEN_86 ? _groups_0_T_12 : _GEN_351; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_13 = {phv_data_172,phv_data_173,phv_data_174,phv_data_175}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_353 = 8'h5b == _GEN_86 ? _groups_0_T_13 : _GEN_352; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_14 = {phv_data_176,phv_data_177,phv_data_178,phv_data_179}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_354 = 8'h5c == _GEN_86 ? _groups_0_T_14 : _GEN_353; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_15 = {phv_data_180,phv_data_181,phv_data_182,phv_data_183}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_355 = 8'h5d == _GEN_86 ? _groups_0_T_15 : _GEN_354; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_16 = {phv_data_184,phv_data_185,phv_data_186,phv_data_187}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_356 = 8'h5e == _GEN_86 ? _groups_0_T_16 : _GEN_355; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_17 = {phv_data_188,phv_data_189,phv_data_190,phv_data_191}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_357 = 8'h5f == _GEN_86 ? _groups_0_T_17 : _GEN_356; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_18 = {phv_data_192,phv_data_193,phv_data_194,phv_data_195}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_358 = 8'h60 == _GEN_86 ? _groups_0_T_18 : _GEN_357; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_19 = {phv_data_196,phv_data_197,phv_data_198,phv_data_199}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_359 = 8'h61 == _GEN_86 ? _groups_0_T_19 : _GEN_358; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_20 = {phv_data_200,phv_data_201,phv_data_202,phv_data_203}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_360 = 8'h62 == _GEN_86 ? _groups_0_T_20 : _GEN_359; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_21 = {phv_data_204,phv_data_205,phv_data_206,phv_data_207}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_361 = 8'h63 == _GEN_86 ? _groups_0_T_21 : _GEN_360; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_22 = {phv_data_208,phv_data_209,phv_data_210,phv_data_211}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_362 = 8'h64 == _GEN_86 ? _groups_0_T_22 : _GEN_361; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_23 = {phv_data_212,phv_data_213,phv_data_214,phv_data_215}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_363 = 8'h65 == _GEN_86 ? _groups_0_T_23 : _GEN_362; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_24 = {phv_data_216,phv_data_217,phv_data_218,phv_data_219}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_364 = 8'h66 == _GEN_86 ? _groups_0_T_24 : _GEN_363; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_25 = {phv_data_220,phv_data_221,phv_data_222,phv_data_223}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_365 = 8'h67 == _GEN_86 ? _groups_0_T_25 : _GEN_364; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_26 = {phv_data_224,phv_data_225,phv_data_226,phv_data_227}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_366 = 8'h68 == _GEN_86 ? _groups_0_T_26 : _GEN_365; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_27 = {phv_data_228,phv_data_229,phv_data_230,phv_data_231}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_367 = 8'h69 == _GEN_86 ? _groups_0_T_27 : _GEN_366; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_28 = {phv_data_232,phv_data_233,phv_data_234,phv_data_235}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_368 = 8'h6a == _GEN_86 ? _groups_0_T_28 : _GEN_367; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_29 = {phv_data_236,phv_data_237,phv_data_238,phv_data_239}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_369 = 8'h6b == _GEN_86 ? _groups_0_T_29 : _GEN_368; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_30 = {phv_data_240,phv_data_241,phv_data_242,phv_data_243}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_370 = 8'h6c == _GEN_86 ? _groups_0_T_30 : _GEN_369; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_31 = {phv_data_244,phv_data_245,phv_data_246,phv_data_247}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_371 = 8'h6d == _GEN_86 ? _groups_0_T_31 : _GEN_370; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_32 = {phv_data_248,phv_data_249,phv_data_250,phv_data_251}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_372 = 8'h6e == _GEN_86 ? _groups_0_T_32 : _GEN_371; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _groups_0_T_33 = {phv_data_252,phv_data_253,phv_data_254,phv_data_255}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_373 = 8'h6f == _GEN_86 ? _groups_0_T_33 : _GEN_372; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] groups_0 = _GEN_56 == 2'h3 ? _GEN_373 : _GEN_341; // @[matcher_pisa.scala 155:50]
  wire [7:0] _GEN_375 = 8'h0 == _GEN_90 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_376 = 8'h1 == _GEN_90 ? phv_data_1 : _GEN_375; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_377 = 8'h2 == _GEN_90 ? phv_data_2 : _GEN_376; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_378 = 8'h3 == _GEN_90 ? phv_data_3 : _GEN_377; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_379 = 8'h4 == _GEN_90 ? phv_data_4 : _GEN_378; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_380 = 8'h5 == _GEN_90 ? phv_data_5 : _GEN_379; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_381 = 8'h6 == _GEN_90 ? phv_data_6 : _GEN_380; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_382 = 8'h7 == _GEN_90 ? phv_data_7 : _GEN_381; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_383 = 8'h8 == _GEN_90 ? phv_data_8 : _GEN_382; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_384 = 8'h9 == _GEN_90 ? phv_data_9 : _GEN_383; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_385 = 8'ha == _GEN_90 ? phv_data_10 : _GEN_384; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_386 = 8'hb == _GEN_90 ? phv_data_11 : _GEN_385; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_387 = 8'hc == _GEN_90 ? phv_data_12 : _GEN_386; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_388 = 8'hd == _GEN_90 ? phv_data_13 : _GEN_387; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_389 = 8'he == _GEN_90 ? phv_data_14 : _GEN_388; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_390 = 8'hf == _GEN_90 ? phv_data_15 : _GEN_389; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_391 = 8'h10 == _GEN_90 ? phv_data_16 : _GEN_390; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_392 = 8'h11 == _GEN_90 ? phv_data_17 : _GEN_391; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_393 = 8'h12 == _GEN_90 ? phv_data_18 : _GEN_392; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_394 = 8'h13 == _GEN_90 ? phv_data_19 : _GEN_393; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_395 = 8'h14 == _GEN_90 ? phv_data_20 : _GEN_394; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_396 = 8'h15 == _GEN_90 ? phv_data_21 : _GEN_395; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_397 = 8'h16 == _GEN_90 ? phv_data_22 : _GEN_396; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_398 = 8'h17 == _GEN_90 ? phv_data_23 : _GEN_397; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_399 = 8'h18 == _GEN_90 ? phv_data_24 : _GEN_398; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_400 = 8'h19 == _GEN_90 ? phv_data_25 : _GEN_399; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_401 = 8'h1a == _GEN_90 ? phv_data_26 : _GEN_400; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_402 = 8'h1b == _GEN_90 ? phv_data_27 : _GEN_401; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_403 = 8'h1c == _GEN_90 ? phv_data_28 : _GEN_402; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_404 = 8'h1d == _GEN_90 ? phv_data_29 : _GEN_403; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_405 = 8'h1e == _GEN_90 ? phv_data_30 : _GEN_404; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_406 = 8'h1f == _GEN_90 ? phv_data_31 : _GEN_405; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_1_0 = _GEN_66 ? _GEN_406 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_408 = 8'h0 == _GEN_91 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_409 = 8'h1 == _GEN_91 ? phv_data_1 : _GEN_408; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_410 = 8'h2 == _GEN_91 ? phv_data_2 : _GEN_409; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_411 = 8'h3 == _GEN_91 ? phv_data_3 : _GEN_410; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_412 = 8'h4 == _GEN_91 ? phv_data_4 : _GEN_411; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_413 = 8'h5 == _GEN_91 ? phv_data_5 : _GEN_412; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_414 = 8'h6 == _GEN_91 ? phv_data_6 : _GEN_413; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_415 = 8'h7 == _GEN_91 ? phv_data_7 : _GEN_414; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_416 = 8'h8 == _GEN_91 ? phv_data_8 : _GEN_415; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_417 = 8'h9 == _GEN_91 ? phv_data_9 : _GEN_416; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_418 = 8'ha == _GEN_91 ? phv_data_10 : _GEN_417; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_419 = 8'hb == _GEN_91 ? phv_data_11 : _GEN_418; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_420 = 8'hc == _GEN_91 ? phv_data_12 : _GEN_419; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_421 = 8'hd == _GEN_91 ? phv_data_13 : _GEN_420; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_422 = 8'he == _GEN_91 ? phv_data_14 : _GEN_421; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_423 = 8'hf == _GEN_91 ? phv_data_15 : _GEN_422; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_424 = 8'h10 == _GEN_91 ? phv_data_16 : _GEN_423; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_425 = 8'h11 == _GEN_91 ? phv_data_17 : _GEN_424; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_426 = 8'h12 == _GEN_91 ? phv_data_18 : _GEN_425; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_427 = 8'h13 == _GEN_91 ? phv_data_19 : _GEN_426; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_428 = 8'h14 == _GEN_91 ? phv_data_20 : _GEN_427; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_429 = 8'h15 == _GEN_91 ? phv_data_21 : _GEN_428; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_430 = 8'h16 == _GEN_91 ? phv_data_22 : _GEN_429; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_431 = 8'h17 == _GEN_91 ? phv_data_23 : _GEN_430; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_432 = 8'h18 == _GEN_91 ? phv_data_24 : _GEN_431; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_433 = 8'h19 == _GEN_91 ? phv_data_25 : _GEN_432; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_434 = 8'h1a == _GEN_91 ? phv_data_26 : _GEN_433; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_435 = 8'h1b == _GEN_91 ? phv_data_27 : _GEN_434; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_436 = 8'h1c == _GEN_91 ? phv_data_28 : _GEN_435; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_437 = 8'h1d == _GEN_91 ? phv_data_29 : _GEN_436; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_438 = 8'h1e == _GEN_91 ? phv_data_30 : _GEN_437; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_439 = 8'h1f == _GEN_91 ? phv_data_31 : _GEN_438; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_1_1 = _GEN_67 ? _GEN_439 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_441 = 8'h0 == _GEN_92 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_442 = 8'h1 == _GEN_92 ? phv_data_1 : _GEN_441; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_443 = 8'h2 == _GEN_92 ? phv_data_2 : _GEN_442; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_444 = 8'h3 == _GEN_92 ? phv_data_3 : _GEN_443; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_445 = 8'h4 == _GEN_92 ? phv_data_4 : _GEN_444; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_446 = 8'h5 == _GEN_92 ? phv_data_5 : _GEN_445; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_447 = 8'h6 == _GEN_92 ? phv_data_6 : _GEN_446; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_448 = 8'h7 == _GEN_92 ? phv_data_7 : _GEN_447; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_449 = 8'h8 == _GEN_92 ? phv_data_8 : _GEN_448; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_450 = 8'h9 == _GEN_92 ? phv_data_9 : _GEN_449; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_451 = 8'ha == _GEN_92 ? phv_data_10 : _GEN_450; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_452 = 8'hb == _GEN_92 ? phv_data_11 : _GEN_451; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_453 = 8'hc == _GEN_92 ? phv_data_12 : _GEN_452; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_454 = 8'hd == _GEN_92 ? phv_data_13 : _GEN_453; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_455 = 8'he == _GEN_92 ? phv_data_14 : _GEN_454; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_456 = 8'hf == _GEN_92 ? phv_data_15 : _GEN_455; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_457 = 8'h10 == _GEN_92 ? phv_data_16 : _GEN_456; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_458 = 8'h11 == _GEN_92 ? phv_data_17 : _GEN_457; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_459 = 8'h12 == _GEN_92 ? phv_data_18 : _GEN_458; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_460 = 8'h13 == _GEN_92 ? phv_data_19 : _GEN_459; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_461 = 8'h14 == _GEN_92 ? phv_data_20 : _GEN_460; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_462 = 8'h15 == _GEN_92 ? phv_data_21 : _GEN_461; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_463 = 8'h16 == _GEN_92 ? phv_data_22 : _GEN_462; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_464 = 8'h17 == _GEN_92 ? phv_data_23 : _GEN_463; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_465 = 8'h18 == _GEN_92 ? phv_data_24 : _GEN_464; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_466 = 8'h19 == _GEN_92 ? phv_data_25 : _GEN_465; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_467 = 8'h1a == _GEN_92 ? phv_data_26 : _GEN_466; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_468 = 8'h1b == _GEN_92 ? phv_data_27 : _GEN_467; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_469 = 8'h1c == _GEN_92 ? phv_data_28 : _GEN_468; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_470 = 8'h1d == _GEN_92 ? phv_data_29 : _GEN_469; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_471 = 8'h1e == _GEN_92 ? phv_data_30 : _GEN_470; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_472 = 8'h1f == _GEN_92 ? phv_data_31 : _GEN_471; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_1_2 = _GEN_68 ? _GEN_472 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_474 = 8'h0 == _GEN_93 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_475 = 8'h1 == _GEN_93 ? phv_data_1 : _GEN_474; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_476 = 8'h2 == _GEN_93 ? phv_data_2 : _GEN_475; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_477 = 8'h3 == _GEN_93 ? phv_data_3 : _GEN_476; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_478 = 8'h4 == _GEN_93 ? phv_data_4 : _GEN_477; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_479 = 8'h5 == _GEN_93 ? phv_data_5 : _GEN_478; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_480 = 8'h6 == _GEN_93 ? phv_data_6 : _GEN_479; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_481 = 8'h7 == _GEN_93 ? phv_data_7 : _GEN_480; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_482 = 8'h8 == _GEN_93 ? phv_data_8 : _GEN_481; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_483 = 8'h9 == _GEN_93 ? phv_data_9 : _GEN_482; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_484 = 8'ha == _GEN_93 ? phv_data_10 : _GEN_483; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_485 = 8'hb == _GEN_93 ? phv_data_11 : _GEN_484; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_486 = 8'hc == _GEN_93 ? phv_data_12 : _GEN_485; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_487 = 8'hd == _GEN_93 ? phv_data_13 : _GEN_486; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_488 = 8'he == _GEN_93 ? phv_data_14 : _GEN_487; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_489 = 8'hf == _GEN_93 ? phv_data_15 : _GEN_488; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_490 = 8'h10 == _GEN_93 ? phv_data_16 : _GEN_489; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_491 = 8'h11 == _GEN_93 ? phv_data_17 : _GEN_490; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_492 = 8'h12 == _GEN_93 ? phv_data_18 : _GEN_491; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_493 = 8'h13 == _GEN_93 ? phv_data_19 : _GEN_492; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_494 = 8'h14 == _GEN_93 ? phv_data_20 : _GEN_493; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_495 = 8'h15 == _GEN_93 ? phv_data_21 : _GEN_494; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_496 = 8'h16 == _GEN_93 ? phv_data_22 : _GEN_495; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_497 = 8'h17 == _GEN_93 ? phv_data_23 : _GEN_496; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_498 = 8'h18 == _GEN_93 ? phv_data_24 : _GEN_497; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_499 = 8'h19 == _GEN_93 ? phv_data_25 : _GEN_498; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_500 = 8'h1a == _GEN_93 ? phv_data_26 : _GEN_499; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_501 = 8'h1b == _GEN_93 ? phv_data_27 : _GEN_500; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_502 = 8'h1c == _GEN_93 ? phv_data_28 : _GEN_501; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_503 = 8'h1d == _GEN_93 ? phv_data_29 : _GEN_502; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_504 = 8'h1e == _GEN_93 ? phv_data_30 : _GEN_503; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_505 = 8'h1f == _GEN_93 ? phv_data_31 : _GEN_504; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_1_3 = _GEN_69 ? _GEN_505 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [31:0] _groups_1_T = {bytes_1_0,bytes_1_1,bytes_1_2,bytes_1_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_507 = _GEN_57 == 2'h1 ? _groups_1_T : 32'h0; // @[matcher_pisa.scala 123:50 matcher_pisa.scala 137:31 matcher_pisa.scala 122:27]
  wire [15:0] _GEN_508 = 8'h20 == _GEN_90 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_509 = 8'h21 == _GEN_90 ? _double_bytes_0_T_1 : _GEN_508; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_510 = 8'h22 == _GEN_90 ? _double_bytes_0_T_2 : _GEN_509; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_511 = 8'h23 == _GEN_90 ? _double_bytes_0_T_3 : _GEN_510; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_512 = 8'h24 == _GEN_90 ? _double_bytes_0_T_4 : _GEN_511; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_513 = 8'h25 == _GEN_90 ? _double_bytes_0_T_5 : _GEN_512; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_514 = 8'h26 == _GEN_90 ? _double_bytes_0_T_6 : _GEN_513; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_515 = 8'h27 == _GEN_90 ? _double_bytes_0_T_7 : _GEN_514; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_516 = 8'h28 == _GEN_90 ? _double_bytes_0_T_8 : _GEN_515; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_517 = 8'h29 == _GEN_90 ? _double_bytes_0_T_9 : _GEN_516; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_518 = 8'h2a == _GEN_90 ? _double_bytes_0_T_10 : _GEN_517; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_519 = 8'h2b == _GEN_90 ? _double_bytes_0_T_11 : _GEN_518; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_520 = 8'h2c == _GEN_90 ? _double_bytes_0_T_12 : _GEN_519; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_521 = 8'h2d == _GEN_90 ? _double_bytes_0_T_13 : _GEN_520; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_522 = 8'h2e == _GEN_90 ? _double_bytes_0_T_14 : _GEN_521; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_523 = 8'h2f == _GEN_90 ? _double_bytes_0_T_15 : _GEN_522; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_524 = 8'h30 == _GEN_90 ? _double_bytes_0_T_16 : _GEN_523; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_525 = 8'h31 == _GEN_90 ? _double_bytes_0_T_17 : _GEN_524; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_526 = 8'h32 == _GEN_90 ? _double_bytes_0_T_18 : _GEN_525; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_527 = 8'h33 == _GEN_90 ? _double_bytes_0_T_19 : _GEN_526; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_528 = 8'h34 == _GEN_90 ? _double_bytes_0_T_20 : _GEN_527; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_529 = 8'h35 == _GEN_90 ? _double_bytes_0_T_21 : _GEN_528; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_530 = 8'h36 == _GEN_90 ? _double_bytes_0_T_22 : _GEN_529; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_531 = 8'h37 == _GEN_90 ? _double_bytes_0_T_23 : _GEN_530; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_532 = 8'h38 == _GEN_90 ? _double_bytes_0_T_24 : _GEN_531; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_533 = 8'h39 == _GEN_90 ? _double_bytes_0_T_25 : _GEN_532; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_534 = 8'h3a == _GEN_90 ? _double_bytes_0_T_26 : _GEN_533; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_535 = 8'h3b == _GEN_90 ? _double_bytes_0_T_27 : _GEN_534; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_536 = 8'h3c == _GEN_90 ? _double_bytes_0_T_28 : _GEN_535; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_537 = 8'h3d == _GEN_90 ? _double_bytes_0_T_29 : _GEN_536; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_538 = 8'h3e == _GEN_90 ? _double_bytes_0_T_30 : _GEN_537; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_539 = 8'h3f == _GEN_90 ? _double_bytes_0_T_31 : _GEN_538; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_540 = 8'h40 == _GEN_90 ? _double_bytes_0_T_32 : _GEN_539; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_541 = 8'h41 == _GEN_90 ? _double_bytes_0_T_33 : _GEN_540; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_542 = 8'h42 == _GEN_90 ? _double_bytes_0_T_34 : _GEN_541; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_543 = 8'h43 == _GEN_90 ? _double_bytes_0_T_35 : _GEN_542; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_544 = 8'h44 == _GEN_90 ? _double_bytes_0_T_36 : _GEN_543; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_545 = 8'h45 == _GEN_90 ? _double_bytes_0_T_37 : _GEN_544; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_546 = 8'h46 == _GEN_90 ? _double_bytes_0_T_38 : _GEN_545; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_547 = 8'h47 == _GEN_90 ? _double_bytes_0_T_39 : _GEN_546; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_548 = 8'h48 == _GEN_90 ? _double_bytes_0_T_40 : _GEN_547; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_549 = 8'h49 == _GEN_90 ? _double_bytes_0_T_41 : _GEN_548; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_550 = 8'h4a == _GEN_90 ? _double_bytes_0_T_42 : _GEN_549; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_551 = 8'h4b == _GEN_90 ? _double_bytes_0_T_43 : _GEN_550; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_552 = 8'h4c == _GEN_90 ? _double_bytes_0_T_44 : _GEN_551; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_553 = 8'h4d == _GEN_90 ? _double_bytes_0_T_45 : _GEN_552; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_554 = 8'h4e == _GEN_90 ? _double_bytes_0_T_46 : _GEN_553; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_555 = 8'h4f == _GEN_90 ? _double_bytes_0_T_47 : _GEN_554; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] double_bytes_1_0 = _GEN_66 ? _GEN_555 : 16'h0; // @[matcher_pisa.scala 145:46 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_557 = 8'h20 == _GEN_91 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_558 = 8'h21 == _GEN_91 ? _double_bytes_0_T_1 : _GEN_557; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_559 = 8'h22 == _GEN_91 ? _double_bytes_0_T_2 : _GEN_558; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_560 = 8'h23 == _GEN_91 ? _double_bytes_0_T_3 : _GEN_559; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_561 = 8'h24 == _GEN_91 ? _double_bytes_0_T_4 : _GEN_560; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_562 = 8'h25 == _GEN_91 ? _double_bytes_0_T_5 : _GEN_561; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_563 = 8'h26 == _GEN_91 ? _double_bytes_0_T_6 : _GEN_562; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_564 = 8'h27 == _GEN_91 ? _double_bytes_0_T_7 : _GEN_563; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_565 = 8'h28 == _GEN_91 ? _double_bytes_0_T_8 : _GEN_564; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_566 = 8'h29 == _GEN_91 ? _double_bytes_0_T_9 : _GEN_565; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_567 = 8'h2a == _GEN_91 ? _double_bytes_0_T_10 : _GEN_566; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_568 = 8'h2b == _GEN_91 ? _double_bytes_0_T_11 : _GEN_567; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_569 = 8'h2c == _GEN_91 ? _double_bytes_0_T_12 : _GEN_568; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_570 = 8'h2d == _GEN_91 ? _double_bytes_0_T_13 : _GEN_569; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_571 = 8'h2e == _GEN_91 ? _double_bytes_0_T_14 : _GEN_570; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_572 = 8'h2f == _GEN_91 ? _double_bytes_0_T_15 : _GEN_571; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_573 = 8'h30 == _GEN_91 ? _double_bytes_0_T_16 : _GEN_572; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_574 = 8'h31 == _GEN_91 ? _double_bytes_0_T_17 : _GEN_573; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_575 = 8'h32 == _GEN_91 ? _double_bytes_0_T_18 : _GEN_574; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_576 = 8'h33 == _GEN_91 ? _double_bytes_0_T_19 : _GEN_575; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_577 = 8'h34 == _GEN_91 ? _double_bytes_0_T_20 : _GEN_576; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_578 = 8'h35 == _GEN_91 ? _double_bytes_0_T_21 : _GEN_577; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_579 = 8'h36 == _GEN_91 ? _double_bytes_0_T_22 : _GEN_578; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_580 = 8'h37 == _GEN_91 ? _double_bytes_0_T_23 : _GEN_579; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_581 = 8'h38 == _GEN_91 ? _double_bytes_0_T_24 : _GEN_580; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_582 = 8'h39 == _GEN_91 ? _double_bytes_0_T_25 : _GEN_581; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_583 = 8'h3a == _GEN_91 ? _double_bytes_0_T_26 : _GEN_582; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_584 = 8'h3b == _GEN_91 ? _double_bytes_0_T_27 : _GEN_583; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_585 = 8'h3c == _GEN_91 ? _double_bytes_0_T_28 : _GEN_584; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_586 = 8'h3d == _GEN_91 ? _double_bytes_0_T_29 : _GEN_585; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_587 = 8'h3e == _GEN_91 ? _double_bytes_0_T_30 : _GEN_586; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_588 = 8'h3f == _GEN_91 ? _double_bytes_0_T_31 : _GEN_587; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_589 = 8'h40 == _GEN_91 ? _double_bytes_0_T_32 : _GEN_588; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_590 = 8'h41 == _GEN_91 ? _double_bytes_0_T_33 : _GEN_589; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_591 = 8'h42 == _GEN_91 ? _double_bytes_0_T_34 : _GEN_590; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_592 = 8'h43 == _GEN_91 ? _double_bytes_0_T_35 : _GEN_591; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_593 = 8'h44 == _GEN_91 ? _double_bytes_0_T_36 : _GEN_592; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_594 = 8'h45 == _GEN_91 ? _double_bytes_0_T_37 : _GEN_593; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_595 = 8'h46 == _GEN_91 ? _double_bytes_0_T_38 : _GEN_594; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_596 = 8'h47 == _GEN_91 ? _double_bytes_0_T_39 : _GEN_595; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_597 = 8'h48 == _GEN_91 ? _double_bytes_0_T_40 : _GEN_596; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_598 = 8'h49 == _GEN_91 ? _double_bytes_0_T_41 : _GEN_597; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_599 = 8'h4a == _GEN_91 ? _double_bytes_0_T_42 : _GEN_598; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_600 = 8'h4b == _GEN_91 ? _double_bytes_0_T_43 : _GEN_599; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_601 = 8'h4c == _GEN_91 ? _double_bytes_0_T_44 : _GEN_600; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_602 = 8'h4d == _GEN_91 ? _double_bytes_0_T_45 : _GEN_601; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_603 = 8'h4e == _GEN_91 ? _double_bytes_0_T_46 : _GEN_602; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_604 = 8'h4f == _GEN_91 ? _double_bytes_0_T_47 : _GEN_603; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] double_bytes_1_1 = _GEN_67 ? _GEN_604 : 16'h0; // @[matcher_pisa.scala 145:46 matcher_pisa.scala 144:41]
  wire [31:0] _groups_1_T_1 = {double_bytes_1_0,double_bytes_1_1}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_606 = _GEN_57 == 2'h2 ? _groups_1_T_1 : _GEN_507; // @[matcher_pisa.scala 139:50 matcher_pisa.scala 153:31]
  wire [31:0] _GEN_607 = 8'h50 == _GEN_90 ? _groups_0_T_2 : 32'h0; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39 matcher_pisa.scala 158:31]
  wire [31:0] _GEN_608 = 8'h51 == _GEN_90 ? _groups_0_T_3 : _GEN_607; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_609 = 8'h52 == _GEN_90 ? _groups_0_T_4 : _GEN_608; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_610 = 8'h53 == _GEN_90 ? _groups_0_T_5 : _GEN_609; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_611 = 8'h54 == _GEN_90 ? _groups_0_T_6 : _GEN_610; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_612 = 8'h55 == _GEN_90 ? _groups_0_T_7 : _GEN_611; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_613 = 8'h56 == _GEN_90 ? _groups_0_T_8 : _GEN_612; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_614 = 8'h57 == _GEN_90 ? _groups_0_T_9 : _GEN_613; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_615 = 8'h58 == _GEN_90 ? _groups_0_T_10 : _GEN_614; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_616 = 8'h59 == _GEN_90 ? _groups_0_T_11 : _GEN_615; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_617 = 8'h5a == _GEN_90 ? _groups_0_T_12 : _GEN_616; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_618 = 8'h5b == _GEN_90 ? _groups_0_T_13 : _GEN_617; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_619 = 8'h5c == _GEN_90 ? _groups_0_T_14 : _GEN_618; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_620 = 8'h5d == _GEN_90 ? _groups_0_T_15 : _GEN_619; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_621 = 8'h5e == _GEN_90 ? _groups_0_T_16 : _GEN_620; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_622 = 8'h5f == _GEN_90 ? _groups_0_T_17 : _GEN_621; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_623 = 8'h60 == _GEN_90 ? _groups_0_T_18 : _GEN_622; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_624 = 8'h61 == _GEN_90 ? _groups_0_T_19 : _GEN_623; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_625 = 8'h62 == _GEN_90 ? _groups_0_T_20 : _GEN_624; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_626 = 8'h63 == _GEN_90 ? _groups_0_T_21 : _GEN_625; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_627 = 8'h64 == _GEN_90 ? _groups_0_T_22 : _GEN_626; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_628 = 8'h65 == _GEN_90 ? _groups_0_T_23 : _GEN_627; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_629 = 8'h66 == _GEN_90 ? _groups_0_T_24 : _GEN_628; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_630 = 8'h67 == _GEN_90 ? _groups_0_T_25 : _GEN_629; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_631 = 8'h68 == _GEN_90 ? _groups_0_T_26 : _GEN_630; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_632 = 8'h69 == _GEN_90 ? _groups_0_T_27 : _GEN_631; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_633 = 8'h6a == _GEN_90 ? _groups_0_T_28 : _GEN_632; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_634 = 8'h6b == _GEN_90 ? _groups_0_T_29 : _GEN_633; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_635 = 8'h6c == _GEN_90 ? _groups_0_T_30 : _GEN_634; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_636 = 8'h6d == _GEN_90 ? _groups_0_T_31 : _GEN_635; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_637 = 8'h6e == _GEN_90 ? _groups_0_T_32 : _GEN_636; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_638 = 8'h6f == _GEN_90 ? _groups_0_T_33 : _GEN_637; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] groups_1 = _GEN_57 == 2'h3 ? _GEN_638 : _GEN_606; // @[matcher_pisa.scala 155:50]
  wire [7:0] _GEN_640 = 8'h0 == _GEN_94 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_641 = 8'h1 == _GEN_94 ? phv_data_1 : _GEN_640; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_642 = 8'h2 == _GEN_94 ? phv_data_2 : _GEN_641; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_643 = 8'h3 == _GEN_94 ? phv_data_3 : _GEN_642; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_644 = 8'h4 == _GEN_94 ? phv_data_4 : _GEN_643; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_645 = 8'h5 == _GEN_94 ? phv_data_5 : _GEN_644; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_646 = 8'h6 == _GEN_94 ? phv_data_6 : _GEN_645; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_647 = 8'h7 == _GEN_94 ? phv_data_7 : _GEN_646; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_648 = 8'h8 == _GEN_94 ? phv_data_8 : _GEN_647; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_649 = 8'h9 == _GEN_94 ? phv_data_9 : _GEN_648; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_650 = 8'ha == _GEN_94 ? phv_data_10 : _GEN_649; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_651 = 8'hb == _GEN_94 ? phv_data_11 : _GEN_650; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_652 = 8'hc == _GEN_94 ? phv_data_12 : _GEN_651; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_653 = 8'hd == _GEN_94 ? phv_data_13 : _GEN_652; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_654 = 8'he == _GEN_94 ? phv_data_14 : _GEN_653; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_655 = 8'hf == _GEN_94 ? phv_data_15 : _GEN_654; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_656 = 8'h10 == _GEN_94 ? phv_data_16 : _GEN_655; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_657 = 8'h11 == _GEN_94 ? phv_data_17 : _GEN_656; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_658 = 8'h12 == _GEN_94 ? phv_data_18 : _GEN_657; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_659 = 8'h13 == _GEN_94 ? phv_data_19 : _GEN_658; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_660 = 8'h14 == _GEN_94 ? phv_data_20 : _GEN_659; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_661 = 8'h15 == _GEN_94 ? phv_data_21 : _GEN_660; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_662 = 8'h16 == _GEN_94 ? phv_data_22 : _GEN_661; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_663 = 8'h17 == _GEN_94 ? phv_data_23 : _GEN_662; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_664 = 8'h18 == _GEN_94 ? phv_data_24 : _GEN_663; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_665 = 8'h19 == _GEN_94 ? phv_data_25 : _GEN_664; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_666 = 8'h1a == _GEN_94 ? phv_data_26 : _GEN_665; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_667 = 8'h1b == _GEN_94 ? phv_data_27 : _GEN_666; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_668 = 8'h1c == _GEN_94 ? phv_data_28 : _GEN_667; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_669 = 8'h1d == _GEN_94 ? phv_data_29 : _GEN_668; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_670 = 8'h1e == _GEN_94 ? phv_data_30 : _GEN_669; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_671 = 8'h1f == _GEN_94 ? phv_data_31 : _GEN_670; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_2_0 = _GEN_70 ? _GEN_671 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_673 = 8'h0 == _GEN_95 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_674 = 8'h1 == _GEN_95 ? phv_data_1 : _GEN_673; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_675 = 8'h2 == _GEN_95 ? phv_data_2 : _GEN_674; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_676 = 8'h3 == _GEN_95 ? phv_data_3 : _GEN_675; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_677 = 8'h4 == _GEN_95 ? phv_data_4 : _GEN_676; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_678 = 8'h5 == _GEN_95 ? phv_data_5 : _GEN_677; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_679 = 8'h6 == _GEN_95 ? phv_data_6 : _GEN_678; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_680 = 8'h7 == _GEN_95 ? phv_data_7 : _GEN_679; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_681 = 8'h8 == _GEN_95 ? phv_data_8 : _GEN_680; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_682 = 8'h9 == _GEN_95 ? phv_data_9 : _GEN_681; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_683 = 8'ha == _GEN_95 ? phv_data_10 : _GEN_682; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_684 = 8'hb == _GEN_95 ? phv_data_11 : _GEN_683; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_685 = 8'hc == _GEN_95 ? phv_data_12 : _GEN_684; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_686 = 8'hd == _GEN_95 ? phv_data_13 : _GEN_685; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_687 = 8'he == _GEN_95 ? phv_data_14 : _GEN_686; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_688 = 8'hf == _GEN_95 ? phv_data_15 : _GEN_687; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_689 = 8'h10 == _GEN_95 ? phv_data_16 : _GEN_688; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_690 = 8'h11 == _GEN_95 ? phv_data_17 : _GEN_689; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_691 = 8'h12 == _GEN_95 ? phv_data_18 : _GEN_690; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_692 = 8'h13 == _GEN_95 ? phv_data_19 : _GEN_691; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_693 = 8'h14 == _GEN_95 ? phv_data_20 : _GEN_692; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_694 = 8'h15 == _GEN_95 ? phv_data_21 : _GEN_693; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_695 = 8'h16 == _GEN_95 ? phv_data_22 : _GEN_694; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_696 = 8'h17 == _GEN_95 ? phv_data_23 : _GEN_695; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_697 = 8'h18 == _GEN_95 ? phv_data_24 : _GEN_696; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_698 = 8'h19 == _GEN_95 ? phv_data_25 : _GEN_697; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_699 = 8'h1a == _GEN_95 ? phv_data_26 : _GEN_698; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_700 = 8'h1b == _GEN_95 ? phv_data_27 : _GEN_699; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_701 = 8'h1c == _GEN_95 ? phv_data_28 : _GEN_700; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_702 = 8'h1d == _GEN_95 ? phv_data_29 : _GEN_701; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_703 = 8'h1e == _GEN_95 ? phv_data_30 : _GEN_702; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_704 = 8'h1f == _GEN_95 ? phv_data_31 : _GEN_703; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_2_1 = _GEN_71 ? _GEN_704 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_706 = 8'h0 == _GEN_96 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_707 = 8'h1 == _GEN_96 ? phv_data_1 : _GEN_706; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_708 = 8'h2 == _GEN_96 ? phv_data_2 : _GEN_707; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_709 = 8'h3 == _GEN_96 ? phv_data_3 : _GEN_708; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_710 = 8'h4 == _GEN_96 ? phv_data_4 : _GEN_709; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_711 = 8'h5 == _GEN_96 ? phv_data_5 : _GEN_710; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_712 = 8'h6 == _GEN_96 ? phv_data_6 : _GEN_711; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_713 = 8'h7 == _GEN_96 ? phv_data_7 : _GEN_712; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_714 = 8'h8 == _GEN_96 ? phv_data_8 : _GEN_713; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_715 = 8'h9 == _GEN_96 ? phv_data_9 : _GEN_714; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_716 = 8'ha == _GEN_96 ? phv_data_10 : _GEN_715; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_717 = 8'hb == _GEN_96 ? phv_data_11 : _GEN_716; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_718 = 8'hc == _GEN_96 ? phv_data_12 : _GEN_717; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_719 = 8'hd == _GEN_96 ? phv_data_13 : _GEN_718; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_720 = 8'he == _GEN_96 ? phv_data_14 : _GEN_719; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_721 = 8'hf == _GEN_96 ? phv_data_15 : _GEN_720; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_722 = 8'h10 == _GEN_96 ? phv_data_16 : _GEN_721; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_723 = 8'h11 == _GEN_96 ? phv_data_17 : _GEN_722; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_724 = 8'h12 == _GEN_96 ? phv_data_18 : _GEN_723; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_725 = 8'h13 == _GEN_96 ? phv_data_19 : _GEN_724; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_726 = 8'h14 == _GEN_96 ? phv_data_20 : _GEN_725; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_727 = 8'h15 == _GEN_96 ? phv_data_21 : _GEN_726; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_728 = 8'h16 == _GEN_96 ? phv_data_22 : _GEN_727; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_729 = 8'h17 == _GEN_96 ? phv_data_23 : _GEN_728; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_730 = 8'h18 == _GEN_96 ? phv_data_24 : _GEN_729; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_731 = 8'h19 == _GEN_96 ? phv_data_25 : _GEN_730; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_732 = 8'h1a == _GEN_96 ? phv_data_26 : _GEN_731; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_733 = 8'h1b == _GEN_96 ? phv_data_27 : _GEN_732; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_734 = 8'h1c == _GEN_96 ? phv_data_28 : _GEN_733; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_735 = 8'h1d == _GEN_96 ? phv_data_29 : _GEN_734; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_736 = 8'h1e == _GEN_96 ? phv_data_30 : _GEN_735; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_737 = 8'h1f == _GEN_96 ? phv_data_31 : _GEN_736; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_2_2 = _GEN_72 ? _GEN_737 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_739 = 8'h0 == _GEN_97 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_740 = 8'h1 == _GEN_97 ? phv_data_1 : _GEN_739; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_741 = 8'h2 == _GEN_97 ? phv_data_2 : _GEN_740; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_742 = 8'h3 == _GEN_97 ? phv_data_3 : _GEN_741; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_743 = 8'h4 == _GEN_97 ? phv_data_4 : _GEN_742; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_744 = 8'h5 == _GEN_97 ? phv_data_5 : _GEN_743; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_745 = 8'h6 == _GEN_97 ? phv_data_6 : _GEN_744; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_746 = 8'h7 == _GEN_97 ? phv_data_7 : _GEN_745; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_747 = 8'h8 == _GEN_97 ? phv_data_8 : _GEN_746; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_748 = 8'h9 == _GEN_97 ? phv_data_9 : _GEN_747; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_749 = 8'ha == _GEN_97 ? phv_data_10 : _GEN_748; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_750 = 8'hb == _GEN_97 ? phv_data_11 : _GEN_749; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_751 = 8'hc == _GEN_97 ? phv_data_12 : _GEN_750; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_752 = 8'hd == _GEN_97 ? phv_data_13 : _GEN_751; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_753 = 8'he == _GEN_97 ? phv_data_14 : _GEN_752; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_754 = 8'hf == _GEN_97 ? phv_data_15 : _GEN_753; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_755 = 8'h10 == _GEN_97 ? phv_data_16 : _GEN_754; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_756 = 8'h11 == _GEN_97 ? phv_data_17 : _GEN_755; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_757 = 8'h12 == _GEN_97 ? phv_data_18 : _GEN_756; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_758 = 8'h13 == _GEN_97 ? phv_data_19 : _GEN_757; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_759 = 8'h14 == _GEN_97 ? phv_data_20 : _GEN_758; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_760 = 8'h15 == _GEN_97 ? phv_data_21 : _GEN_759; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_761 = 8'h16 == _GEN_97 ? phv_data_22 : _GEN_760; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_762 = 8'h17 == _GEN_97 ? phv_data_23 : _GEN_761; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_763 = 8'h18 == _GEN_97 ? phv_data_24 : _GEN_762; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_764 = 8'h19 == _GEN_97 ? phv_data_25 : _GEN_763; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_765 = 8'h1a == _GEN_97 ? phv_data_26 : _GEN_764; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_766 = 8'h1b == _GEN_97 ? phv_data_27 : _GEN_765; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_767 = 8'h1c == _GEN_97 ? phv_data_28 : _GEN_766; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_768 = 8'h1d == _GEN_97 ? phv_data_29 : _GEN_767; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_769 = 8'h1e == _GEN_97 ? phv_data_30 : _GEN_768; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_770 = 8'h1f == _GEN_97 ? phv_data_31 : _GEN_769; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_2_3 = _GEN_73 ? _GEN_770 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [31:0] _groups_2_T = {bytes_2_0,bytes_2_1,bytes_2_2,bytes_2_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_772 = _GEN_58 == 2'h1 ? _groups_2_T : 32'h0; // @[matcher_pisa.scala 123:50 matcher_pisa.scala 137:31 matcher_pisa.scala 122:27]
  wire [15:0] _GEN_773 = 8'h20 == _GEN_94 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_774 = 8'h21 == _GEN_94 ? _double_bytes_0_T_1 : _GEN_773; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_775 = 8'h22 == _GEN_94 ? _double_bytes_0_T_2 : _GEN_774; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_776 = 8'h23 == _GEN_94 ? _double_bytes_0_T_3 : _GEN_775; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_777 = 8'h24 == _GEN_94 ? _double_bytes_0_T_4 : _GEN_776; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_778 = 8'h25 == _GEN_94 ? _double_bytes_0_T_5 : _GEN_777; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_779 = 8'h26 == _GEN_94 ? _double_bytes_0_T_6 : _GEN_778; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_780 = 8'h27 == _GEN_94 ? _double_bytes_0_T_7 : _GEN_779; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_781 = 8'h28 == _GEN_94 ? _double_bytes_0_T_8 : _GEN_780; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_782 = 8'h29 == _GEN_94 ? _double_bytes_0_T_9 : _GEN_781; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_783 = 8'h2a == _GEN_94 ? _double_bytes_0_T_10 : _GEN_782; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_784 = 8'h2b == _GEN_94 ? _double_bytes_0_T_11 : _GEN_783; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_785 = 8'h2c == _GEN_94 ? _double_bytes_0_T_12 : _GEN_784; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_786 = 8'h2d == _GEN_94 ? _double_bytes_0_T_13 : _GEN_785; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_787 = 8'h2e == _GEN_94 ? _double_bytes_0_T_14 : _GEN_786; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_788 = 8'h2f == _GEN_94 ? _double_bytes_0_T_15 : _GEN_787; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_789 = 8'h30 == _GEN_94 ? _double_bytes_0_T_16 : _GEN_788; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_790 = 8'h31 == _GEN_94 ? _double_bytes_0_T_17 : _GEN_789; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_791 = 8'h32 == _GEN_94 ? _double_bytes_0_T_18 : _GEN_790; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_792 = 8'h33 == _GEN_94 ? _double_bytes_0_T_19 : _GEN_791; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_793 = 8'h34 == _GEN_94 ? _double_bytes_0_T_20 : _GEN_792; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_794 = 8'h35 == _GEN_94 ? _double_bytes_0_T_21 : _GEN_793; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_795 = 8'h36 == _GEN_94 ? _double_bytes_0_T_22 : _GEN_794; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_796 = 8'h37 == _GEN_94 ? _double_bytes_0_T_23 : _GEN_795; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_797 = 8'h38 == _GEN_94 ? _double_bytes_0_T_24 : _GEN_796; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_798 = 8'h39 == _GEN_94 ? _double_bytes_0_T_25 : _GEN_797; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_799 = 8'h3a == _GEN_94 ? _double_bytes_0_T_26 : _GEN_798; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_800 = 8'h3b == _GEN_94 ? _double_bytes_0_T_27 : _GEN_799; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_801 = 8'h3c == _GEN_94 ? _double_bytes_0_T_28 : _GEN_800; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_802 = 8'h3d == _GEN_94 ? _double_bytes_0_T_29 : _GEN_801; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_803 = 8'h3e == _GEN_94 ? _double_bytes_0_T_30 : _GEN_802; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_804 = 8'h3f == _GEN_94 ? _double_bytes_0_T_31 : _GEN_803; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_805 = 8'h40 == _GEN_94 ? _double_bytes_0_T_32 : _GEN_804; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_806 = 8'h41 == _GEN_94 ? _double_bytes_0_T_33 : _GEN_805; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_807 = 8'h42 == _GEN_94 ? _double_bytes_0_T_34 : _GEN_806; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_808 = 8'h43 == _GEN_94 ? _double_bytes_0_T_35 : _GEN_807; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_809 = 8'h44 == _GEN_94 ? _double_bytes_0_T_36 : _GEN_808; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_810 = 8'h45 == _GEN_94 ? _double_bytes_0_T_37 : _GEN_809; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_811 = 8'h46 == _GEN_94 ? _double_bytes_0_T_38 : _GEN_810; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_812 = 8'h47 == _GEN_94 ? _double_bytes_0_T_39 : _GEN_811; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_813 = 8'h48 == _GEN_94 ? _double_bytes_0_T_40 : _GEN_812; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_814 = 8'h49 == _GEN_94 ? _double_bytes_0_T_41 : _GEN_813; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_815 = 8'h4a == _GEN_94 ? _double_bytes_0_T_42 : _GEN_814; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_816 = 8'h4b == _GEN_94 ? _double_bytes_0_T_43 : _GEN_815; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_817 = 8'h4c == _GEN_94 ? _double_bytes_0_T_44 : _GEN_816; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_818 = 8'h4d == _GEN_94 ? _double_bytes_0_T_45 : _GEN_817; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_819 = 8'h4e == _GEN_94 ? _double_bytes_0_T_46 : _GEN_818; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_820 = 8'h4f == _GEN_94 ? _double_bytes_0_T_47 : _GEN_819; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] double_bytes_2_0 = _GEN_70 ? _GEN_820 : 16'h0; // @[matcher_pisa.scala 145:46 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_822 = 8'h20 == _GEN_95 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_823 = 8'h21 == _GEN_95 ? _double_bytes_0_T_1 : _GEN_822; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_824 = 8'h22 == _GEN_95 ? _double_bytes_0_T_2 : _GEN_823; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_825 = 8'h23 == _GEN_95 ? _double_bytes_0_T_3 : _GEN_824; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_826 = 8'h24 == _GEN_95 ? _double_bytes_0_T_4 : _GEN_825; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_827 = 8'h25 == _GEN_95 ? _double_bytes_0_T_5 : _GEN_826; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_828 = 8'h26 == _GEN_95 ? _double_bytes_0_T_6 : _GEN_827; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_829 = 8'h27 == _GEN_95 ? _double_bytes_0_T_7 : _GEN_828; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_830 = 8'h28 == _GEN_95 ? _double_bytes_0_T_8 : _GEN_829; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_831 = 8'h29 == _GEN_95 ? _double_bytes_0_T_9 : _GEN_830; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_832 = 8'h2a == _GEN_95 ? _double_bytes_0_T_10 : _GEN_831; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_833 = 8'h2b == _GEN_95 ? _double_bytes_0_T_11 : _GEN_832; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_834 = 8'h2c == _GEN_95 ? _double_bytes_0_T_12 : _GEN_833; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_835 = 8'h2d == _GEN_95 ? _double_bytes_0_T_13 : _GEN_834; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_836 = 8'h2e == _GEN_95 ? _double_bytes_0_T_14 : _GEN_835; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_837 = 8'h2f == _GEN_95 ? _double_bytes_0_T_15 : _GEN_836; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_838 = 8'h30 == _GEN_95 ? _double_bytes_0_T_16 : _GEN_837; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_839 = 8'h31 == _GEN_95 ? _double_bytes_0_T_17 : _GEN_838; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_840 = 8'h32 == _GEN_95 ? _double_bytes_0_T_18 : _GEN_839; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_841 = 8'h33 == _GEN_95 ? _double_bytes_0_T_19 : _GEN_840; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_842 = 8'h34 == _GEN_95 ? _double_bytes_0_T_20 : _GEN_841; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_843 = 8'h35 == _GEN_95 ? _double_bytes_0_T_21 : _GEN_842; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_844 = 8'h36 == _GEN_95 ? _double_bytes_0_T_22 : _GEN_843; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_845 = 8'h37 == _GEN_95 ? _double_bytes_0_T_23 : _GEN_844; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_846 = 8'h38 == _GEN_95 ? _double_bytes_0_T_24 : _GEN_845; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_847 = 8'h39 == _GEN_95 ? _double_bytes_0_T_25 : _GEN_846; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_848 = 8'h3a == _GEN_95 ? _double_bytes_0_T_26 : _GEN_847; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_849 = 8'h3b == _GEN_95 ? _double_bytes_0_T_27 : _GEN_848; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_850 = 8'h3c == _GEN_95 ? _double_bytes_0_T_28 : _GEN_849; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_851 = 8'h3d == _GEN_95 ? _double_bytes_0_T_29 : _GEN_850; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_852 = 8'h3e == _GEN_95 ? _double_bytes_0_T_30 : _GEN_851; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_853 = 8'h3f == _GEN_95 ? _double_bytes_0_T_31 : _GEN_852; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_854 = 8'h40 == _GEN_95 ? _double_bytes_0_T_32 : _GEN_853; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_855 = 8'h41 == _GEN_95 ? _double_bytes_0_T_33 : _GEN_854; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_856 = 8'h42 == _GEN_95 ? _double_bytes_0_T_34 : _GEN_855; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_857 = 8'h43 == _GEN_95 ? _double_bytes_0_T_35 : _GEN_856; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_858 = 8'h44 == _GEN_95 ? _double_bytes_0_T_36 : _GEN_857; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_859 = 8'h45 == _GEN_95 ? _double_bytes_0_T_37 : _GEN_858; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_860 = 8'h46 == _GEN_95 ? _double_bytes_0_T_38 : _GEN_859; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_861 = 8'h47 == _GEN_95 ? _double_bytes_0_T_39 : _GEN_860; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_862 = 8'h48 == _GEN_95 ? _double_bytes_0_T_40 : _GEN_861; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_863 = 8'h49 == _GEN_95 ? _double_bytes_0_T_41 : _GEN_862; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_864 = 8'h4a == _GEN_95 ? _double_bytes_0_T_42 : _GEN_863; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_865 = 8'h4b == _GEN_95 ? _double_bytes_0_T_43 : _GEN_864; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_866 = 8'h4c == _GEN_95 ? _double_bytes_0_T_44 : _GEN_865; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_867 = 8'h4d == _GEN_95 ? _double_bytes_0_T_45 : _GEN_866; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_868 = 8'h4e == _GEN_95 ? _double_bytes_0_T_46 : _GEN_867; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_869 = 8'h4f == _GEN_95 ? _double_bytes_0_T_47 : _GEN_868; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] double_bytes_2_1 = _GEN_71 ? _GEN_869 : 16'h0; // @[matcher_pisa.scala 145:46 matcher_pisa.scala 144:41]
  wire [31:0] _groups_2_T_1 = {double_bytes_2_0,double_bytes_2_1}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_871 = _GEN_58 == 2'h2 ? _groups_2_T_1 : _GEN_772; // @[matcher_pisa.scala 139:50 matcher_pisa.scala 153:31]
  wire [31:0] _GEN_872 = 8'h50 == _GEN_94 ? _groups_0_T_2 : 32'h0; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39 matcher_pisa.scala 158:31]
  wire [31:0] _GEN_873 = 8'h51 == _GEN_94 ? _groups_0_T_3 : _GEN_872; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_874 = 8'h52 == _GEN_94 ? _groups_0_T_4 : _GEN_873; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_875 = 8'h53 == _GEN_94 ? _groups_0_T_5 : _GEN_874; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_876 = 8'h54 == _GEN_94 ? _groups_0_T_6 : _GEN_875; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_877 = 8'h55 == _GEN_94 ? _groups_0_T_7 : _GEN_876; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_878 = 8'h56 == _GEN_94 ? _groups_0_T_8 : _GEN_877; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_879 = 8'h57 == _GEN_94 ? _groups_0_T_9 : _GEN_878; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_880 = 8'h58 == _GEN_94 ? _groups_0_T_10 : _GEN_879; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_881 = 8'h59 == _GEN_94 ? _groups_0_T_11 : _GEN_880; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_882 = 8'h5a == _GEN_94 ? _groups_0_T_12 : _GEN_881; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_883 = 8'h5b == _GEN_94 ? _groups_0_T_13 : _GEN_882; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_884 = 8'h5c == _GEN_94 ? _groups_0_T_14 : _GEN_883; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_885 = 8'h5d == _GEN_94 ? _groups_0_T_15 : _GEN_884; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_886 = 8'h5e == _GEN_94 ? _groups_0_T_16 : _GEN_885; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_887 = 8'h5f == _GEN_94 ? _groups_0_T_17 : _GEN_886; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_888 = 8'h60 == _GEN_94 ? _groups_0_T_18 : _GEN_887; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_889 = 8'h61 == _GEN_94 ? _groups_0_T_19 : _GEN_888; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_890 = 8'h62 == _GEN_94 ? _groups_0_T_20 : _GEN_889; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_891 = 8'h63 == _GEN_94 ? _groups_0_T_21 : _GEN_890; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_892 = 8'h64 == _GEN_94 ? _groups_0_T_22 : _GEN_891; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_893 = 8'h65 == _GEN_94 ? _groups_0_T_23 : _GEN_892; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_894 = 8'h66 == _GEN_94 ? _groups_0_T_24 : _GEN_893; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_895 = 8'h67 == _GEN_94 ? _groups_0_T_25 : _GEN_894; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_896 = 8'h68 == _GEN_94 ? _groups_0_T_26 : _GEN_895; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_897 = 8'h69 == _GEN_94 ? _groups_0_T_27 : _GEN_896; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_898 = 8'h6a == _GEN_94 ? _groups_0_T_28 : _GEN_897; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_899 = 8'h6b == _GEN_94 ? _groups_0_T_29 : _GEN_898; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_900 = 8'h6c == _GEN_94 ? _groups_0_T_30 : _GEN_899; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_901 = 8'h6d == _GEN_94 ? _groups_0_T_31 : _GEN_900; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_902 = 8'h6e == _GEN_94 ? _groups_0_T_32 : _GEN_901; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_903 = 8'h6f == _GEN_94 ? _groups_0_T_33 : _GEN_902; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] groups_2 = _GEN_58 == 2'h3 ? _GEN_903 : _GEN_871; // @[matcher_pisa.scala 155:50]
  wire [7:0] _GEN_905 = 8'h0 == _GEN_98 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_906 = 8'h1 == _GEN_98 ? phv_data_1 : _GEN_905; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_907 = 8'h2 == _GEN_98 ? phv_data_2 : _GEN_906; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_908 = 8'h3 == _GEN_98 ? phv_data_3 : _GEN_907; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_909 = 8'h4 == _GEN_98 ? phv_data_4 : _GEN_908; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_910 = 8'h5 == _GEN_98 ? phv_data_5 : _GEN_909; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_911 = 8'h6 == _GEN_98 ? phv_data_6 : _GEN_910; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_912 = 8'h7 == _GEN_98 ? phv_data_7 : _GEN_911; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_913 = 8'h8 == _GEN_98 ? phv_data_8 : _GEN_912; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_914 = 8'h9 == _GEN_98 ? phv_data_9 : _GEN_913; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_915 = 8'ha == _GEN_98 ? phv_data_10 : _GEN_914; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_916 = 8'hb == _GEN_98 ? phv_data_11 : _GEN_915; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_917 = 8'hc == _GEN_98 ? phv_data_12 : _GEN_916; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_918 = 8'hd == _GEN_98 ? phv_data_13 : _GEN_917; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_919 = 8'he == _GEN_98 ? phv_data_14 : _GEN_918; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_920 = 8'hf == _GEN_98 ? phv_data_15 : _GEN_919; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_921 = 8'h10 == _GEN_98 ? phv_data_16 : _GEN_920; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_922 = 8'h11 == _GEN_98 ? phv_data_17 : _GEN_921; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_923 = 8'h12 == _GEN_98 ? phv_data_18 : _GEN_922; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_924 = 8'h13 == _GEN_98 ? phv_data_19 : _GEN_923; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_925 = 8'h14 == _GEN_98 ? phv_data_20 : _GEN_924; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_926 = 8'h15 == _GEN_98 ? phv_data_21 : _GEN_925; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_927 = 8'h16 == _GEN_98 ? phv_data_22 : _GEN_926; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_928 = 8'h17 == _GEN_98 ? phv_data_23 : _GEN_927; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_929 = 8'h18 == _GEN_98 ? phv_data_24 : _GEN_928; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_930 = 8'h19 == _GEN_98 ? phv_data_25 : _GEN_929; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_931 = 8'h1a == _GEN_98 ? phv_data_26 : _GEN_930; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_932 = 8'h1b == _GEN_98 ? phv_data_27 : _GEN_931; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_933 = 8'h1c == _GEN_98 ? phv_data_28 : _GEN_932; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_934 = 8'h1d == _GEN_98 ? phv_data_29 : _GEN_933; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_935 = 8'h1e == _GEN_98 ? phv_data_30 : _GEN_934; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_936 = 8'h1f == _GEN_98 ? phv_data_31 : _GEN_935; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_3_0 = _GEN_74 ? _GEN_936 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_938 = 8'h0 == _GEN_99 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_939 = 8'h1 == _GEN_99 ? phv_data_1 : _GEN_938; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_940 = 8'h2 == _GEN_99 ? phv_data_2 : _GEN_939; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_941 = 8'h3 == _GEN_99 ? phv_data_3 : _GEN_940; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_942 = 8'h4 == _GEN_99 ? phv_data_4 : _GEN_941; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_943 = 8'h5 == _GEN_99 ? phv_data_5 : _GEN_942; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_944 = 8'h6 == _GEN_99 ? phv_data_6 : _GEN_943; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_945 = 8'h7 == _GEN_99 ? phv_data_7 : _GEN_944; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_946 = 8'h8 == _GEN_99 ? phv_data_8 : _GEN_945; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_947 = 8'h9 == _GEN_99 ? phv_data_9 : _GEN_946; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_948 = 8'ha == _GEN_99 ? phv_data_10 : _GEN_947; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_949 = 8'hb == _GEN_99 ? phv_data_11 : _GEN_948; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_950 = 8'hc == _GEN_99 ? phv_data_12 : _GEN_949; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_951 = 8'hd == _GEN_99 ? phv_data_13 : _GEN_950; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_952 = 8'he == _GEN_99 ? phv_data_14 : _GEN_951; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_953 = 8'hf == _GEN_99 ? phv_data_15 : _GEN_952; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_954 = 8'h10 == _GEN_99 ? phv_data_16 : _GEN_953; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_955 = 8'h11 == _GEN_99 ? phv_data_17 : _GEN_954; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_956 = 8'h12 == _GEN_99 ? phv_data_18 : _GEN_955; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_957 = 8'h13 == _GEN_99 ? phv_data_19 : _GEN_956; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_958 = 8'h14 == _GEN_99 ? phv_data_20 : _GEN_957; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_959 = 8'h15 == _GEN_99 ? phv_data_21 : _GEN_958; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_960 = 8'h16 == _GEN_99 ? phv_data_22 : _GEN_959; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_961 = 8'h17 == _GEN_99 ? phv_data_23 : _GEN_960; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_962 = 8'h18 == _GEN_99 ? phv_data_24 : _GEN_961; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_963 = 8'h19 == _GEN_99 ? phv_data_25 : _GEN_962; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_964 = 8'h1a == _GEN_99 ? phv_data_26 : _GEN_963; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_965 = 8'h1b == _GEN_99 ? phv_data_27 : _GEN_964; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_966 = 8'h1c == _GEN_99 ? phv_data_28 : _GEN_965; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_967 = 8'h1d == _GEN_99 ? phv_data_29 : _GEN_966; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_968 = 8'h1e == _GEN_99 ? phv_data_30 : _GEN_967; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_969 = 8'h1f == _GEN_99 ? phv_data_31 : _GEN_968; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_3_1 = _GEN_75 ? _GEN_969 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_971 = 8'h0 == _GEN_100 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_972 = 8'h1 == _GEN_100 ? phv_data_1 : _GEN_971; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_973 = 8'h2 == _GEN_100 ? phv_data_2 : _GEN_972; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_974 = 8'h3 == _GEN_100 ? phv_data_3 : _GEN_973; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_975 = 8'h4 == _GEN_100 ? phv_data_4 : _GEN_974; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_976 = 8'h5 == _GEN_100 ? phv_data_5 : _GEN_975; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_977 = 8'h6 == _GEN_100 ? phv_data_6 : _GEN_976; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_978 = 8'h7 == _GEN_100 ? phv_data_7 : _GEN_977; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_979 = 8'h8 == _GEN_100 ? phv_data_8 : _GEN_978; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_980 = 8'h9 == _GEN_100 ? phv_data_9 : _GEN_979; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_981 = 8'ha == _GEN_100 ? phv_data_10 : _GEN_980; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_982 = 8'hb == _GEN_100 ? phv_data_11 : _GEN_981; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_983 = 8'hc == _GEN_100 ? phv_data_12 : _GEN_982; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_984 = 8'hd == _GEN_100 ? phv_data_13 : _GEN_983; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_985 = 8'he == _GEN_100 ? phv_data_14 : _GEN_984; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_986 = 8'hf == _GEN_100 ? phv_data_15 : _GEN_985; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_987 = 8'h10 == _GEN_100 ? phv_data_16 : _GEN_986; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_988 = 8'h11 == _GEN_100 ? phv_data_17 : _GEN_987; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_989 = 8'h12 == _GEN_100 ? phv_data_18 : _GEN_988; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_990 = 8'h13 == _GEN_100 ? phv_data_19 : _GEN_989; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_991 = 8'h14 == _GEN_100 ? phv_data_20 : _GEN_990; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_992 = 8'h15 == _GEN_100 ? phv_data_21 : _GEN_991; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_993 = 8'h16 == _GEN_100 ? phv_data_22 : _GEN_992; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_994 = 8'h17 == _GEN_100 ? phv_data_23 : _GEN_993; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_995 = 8'h18 == _GEN_100 ? phv_data_24 : _GEN_994; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_996 = 8'h19 == _GEN_100 ? phv_data_25 : _GEN_995; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_997 = 8'h1a == _GEN_100 ? phv_data_26 : _GEN_996; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_998 = 8'h1b == _GEN_100 ? phv_data_27 : _GEN_997; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_999 = 8'h1c == _GEN_100 ? phv_data_28 : _GEN_998; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1000 = 8'h1d == _GEN_100 ? phv_data_29 : _GEN_999; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1001 = 8'h1e == _GEN_100 ? phv_data_30 : _GEN_1000; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1002 = 8'h1f == _GEN_100 ? phv_data_31 : _GEN_1001; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_3_2 = _GEN_76 ? _GEN_1002 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1004 = 8'h0 == _GEN_101 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1005 = 8'h1 == _GEN_101 ? phv_data_1 : _GEN_1004; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1006 = 8'h2 == _GEN_101 ? phv_data_2 : _GEN_1005; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1007 = 8'h3 == _GEN_101 ? phv_data_3 : _GEN_1006; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1008 = 8'h4 == _GEN_101 ? phv_data_4 : _GEN_1007; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1009 = 8'h5 == _GEN_101 ? phv_data_5 : _GEN_1008; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1010 = 8'h6 == _GEN_101 ? phv_data_6 : _GEN_1009; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1011 = 8'h7 == _GEN_101 ? phv_data_7 : _GEN_1010; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1012 = 8'h8 == _GEN_101 ? phv_data_8 : _GEN_1011; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1013 = 8'h9 == _GEN_101 ? phv_data_9 : _GEN_1012; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1014 = 8'ha == _GEN_101 ? phv_data_10 : _GEN_1013; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1015 = 8'hb == _GEN_101 ? phv_data_11 : _GEN_1014; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1016 = 8'hc == _GEN_101 ? phv_data_12 : _GEN_1015; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1017 = 8'hd == _GEN_101 ? phv_data_13 : _GEN_1016; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1018 = 8'he == _GEN_101 ? phv_data_14 : _GEN_1017; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1019 = 8'hf == _GEN_101 ? phv_data_15 : _GEN_1018; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1020 = 8'h10 == _GEN_101 ? phv_data_16 : _GEN_1019; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1021 = 8'h11 == _GEN_101 ? phv_data_17 : _GEN_1020; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1022 = 8'h12 == _GEN_101 ? phv_data_18 : _GEN_1021; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1023 = 8'h13 == _GEN_101 ? phv_data_19 : _GEN_1022; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1024 = 8'h14 == _GEN_101 ? phv_data_20 : _GEN_1023; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1025 = 8'h15 == _GEN_101 ? phv_data_21 : _GEN_1024; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1026 = 8'h16 == _GEN_101 ? phv_data_22 : _GEN_1025; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1027 = 8'h17 == _GEN_101 ? phv_data_23 : _GEN_1026; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1028 = 8'h18 == _GEN_101 ? phv_data_24 : _GEN_1027; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1029 = 8'h19 == _GEN_101 ? phv_data_25 : _GEN_1028; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1030 = 8'h1a == _GEN_101 ? phv_data_26 : _GEN_1029; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1031 = 8'h1b == _GEN_101 ? phv_data_27 : _GEN_1030; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1032 = 8'h1c == _GEN_101 ? phv_data_28 : _GEN_1031; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1033 = 8'h1d == _GEN_101 ? phv_data_29 : _GEN_1032; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1034 = 8'h1e == _GEN_101 ? phv_data_30 : _GEN_1033; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1035 = 8'h1f == _GEN_101 ? phv_data_31 : _GEN_1034; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_3_3 = _GEN_77 ? _GEN_1035 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [31:0] _groups_3_T = {bytes_3_0,bytes_3_1,bytes_3_2,bytes_3_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_1037 = _GEN_59 == 2'h1 ? _groups_3_T : 32'h0; // @[matcher_pisa.scala 123:50 matcher_pisa.scala 137:31 matcher_pisa.scala 122:27]
  wire [15:0] _GEN_1038 = 8'h20 == _GEN_98 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_1039 = 8'h21 == _GEN_98 ? _double_bytes_0_T_1 : _GEN_1038; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1040 = 8'h22 == _GEN_98 ? _double_bytes_0_T_2 : _GEN_1039; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1041 = 8'h23 == _GEN_98 ? _double_bytes_0_T_3 : _GEN_1040; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1042 = 8'h24 == _GEN_98 ? _double_bytes_0_T_4 : _GEN_1041; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1043 = 8'h25 == _GEN_98 ? _double_bytes_0_T_5 : _GEN_1042; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1044 = 8'h26 == _GEN_98 ? _double_bytes_0_T_6 : _GEN_1043; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1045 = 8'h27 == _GEN_98 ? _double_bytes_0_T_7 : _GEN_1044; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1046 = 8'h28 == _GEN_98 ? _double_bytes_0_T_8 : _GEN_1045; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1047 = 8'h29 == _GEN_98 ? _double_bytes_0_T_9 : _GEN_1046; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1048 = 8'h2a == _GEN_98 ? _double_bytes_0_T_10 : _GEN_1047; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1049 = 8'h2b == _GEN_98 ? _double_bytes_0_T_11 : _GEN_1048; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1050 = 8'h2c == _GEN_98 ? _double_bytes_0_T_12 : _GEN_1049; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1051 = 8'h2d == _GEN_98 ? _double_bytes_0_T_13 : _GEN_1050; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1052 = 8'h2e == _GEN_98 ? _double_bytes_0_T_14 : _GEN_1051; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1053 = 8'h2f == _GEN_98 ? _double_bytes_0_T_15 : _GEN_1052; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1054 = 8'h30 == _GEN_98 ? _double_bytes_0_T_16 : _GEN_1053; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1055 = 8'h31 == _GEN_98 ? _double_bytes_0_T_17 : _GEN_1054; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1056 = 8'h32 == _GEN_98 ? _double_bytes_0_T_18 : _GEN_1055; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1057 = 8'h33 == _GEN_98 ? _double_bytes_0_T_19 : _GEN_1056; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1058 = 8'h34 == _GEN_98 ? _double_bytes_0_T_20 : _GEN_1057; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1059 = 8'h35 == _GEN_98 ? _double_bytes_0_T_21 : _GEN_1058; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1060 = 8'h36 == _GEN_98 ? _double_bytes_0_T_22 : _GEN_1059; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1061 = 8'h37 == _GEN_98 ? _double_bytes_0_T_23 : _GEN_1060; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1062 = 8'h38 == _GEN_98 ? _double_bytes_0_T_24 : _GEN_1061; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1063 = 8'h39 == _GEN_98 ? _double_bytes_0_T_25 : _GEN_1062; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1064 = 8'h3a == _GEN_98 ? _double_bytes_0_T_26 : _GEN_1063; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1065 = 8'h3b == _GEN_98 ? _double_bytes_0_T_27 : _GEN_1064; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1066 = 8'h3c == _GEN_98 ? _double_bytes_0_T_28 : _GEN_1065; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1067 = 8'h3d == _GEN_98 ? _double_bytes_0_T_29 : _GEN_1066; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1068 = 8'h3e == _GEN_98 ? _double_bytes_0_T_30 : _GEN_1067; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1069 = 8'h3f == _GEN_98 ? _double_bytes_0_T_31 : _GEN_1068; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1070 = 8'h40 == _GEN_98 ? _double_bytes_0_T_32 : _GEN_1069; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1071 = 8'h41 == _GEN_98 ? _double_bytes_0_T_33 : _GEN_1070; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1072 = 8'h42 == _GEN_98 ? _double_bytes_0_T_34 : _GEN_1071; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1073 = 8'h43 == _GEN_98 ? _double_bytes_0_T_35 : _GEN_1072; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1074 = 8'h44 == _GEN_98 ? _double_bytes_0_T_36 : _GEN_1073; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1075 = 8'h45 == _GEN_98 ? _double_bytes_0_T_37 : _GEN_1074; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1076 = 8'h46 == _GEN_98 ? _double_bytes_0_T_38 : _GEN_1075; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1077 = 8'h47 == _GEN_98 ? _double_bytes_0_T_39 : _GEN_1076; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1078 = 8'h48 == _GEN_98 ? _double_bytes_0_T_40 : _GEN_1077; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1079 = 8'h49 == _GEN_98 ? _double_bytes_0_T_41 : _GEN_1078; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1080 = 8'h4a == _GEN_98 ? _double_bytes_0_T_42 : _GEN_1079; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1081 = 8'h4b == _GEN_98 ? _double_bytes_0_T_43 : _GEN_1080; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1082 = 8'h4c == _GEN_98 ? _double_bytes_0_T_44 : _GEN_1081; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1083 = 8'h4d == _GEN_98 ? _double_bytes_0_T_45 : _GEN_1082; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1084 = 8'h4e == _GEN_98 ? _double_bytes_0_T_46 : _GEN_1083; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1085 = 8'h4f == _GEN_98 ? _double_bytes_0_T_47 : _GEN_1084; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] double_bytes_3_0 = _GEN_74 ? _GEN_1085 : 16'h0; // @[matcher_pisa.scala 145:46 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_1087 = 8'h20 == _GEN_99 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_1088 = 8'h21 == _GEN_99 ? _double_bytes_0_T_1 : _GEN_1087; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1089 = 8'h22 == _GEN_99 ? _double_bytes_0_T_2 : _GEN_1088; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1090 = 8'h23 == _GEN_99 ? _double_bytes_0_T_3 : _GEN_1089; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1091 = 8'h24 == _GEN_99 ? _double_bytes_0_T_4 : _GEN_1090; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1092 = 8'h25 == _GEN_99 ? _double_bytes_0_T_5 : _GEN_1091; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1093 = 8'h26 == _GEN_99 ? _double_bytes_0_T_6 : _GEN_1092; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1094 = 8'h27 == _GEN_99 ? _double_bytes_0_T_7 : _GEN_1093; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1095 = 8'h28 == _GEN_99 ? _double_bytes_0_T_8 : _GEN_1094; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1096 = 8'h29 == _GEN_99 ? _double_bytes_0_T_9 : _GEN_1095; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1097 = 8'h2a == _GEN_99 ? _double_bytes_0_T_10 : _GEN_1096; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1098 = 8'h2b == _GEN_99 ? _double_bytes_0_T_11 : _GEN_1097; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1099 = 8'h2c == _GEN_99 ? _double_bytes_0_T_12 : _GEN_1098; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1100 = 8'h2d == _GEN_99 ? _double_bytes_0_T_13 : _GEN_1099; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1101 = 8'h2e == _GEN_99 ? _double_bytes_0_T_14 : _GEN_1100; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1102 = 8'h2f == _GEN_99 ? _double_bytes_0_T_15 : _GEN_1101; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1103 = 8'h30 == _GEN_99 ? _double_bytes_0_T_16 : _GEN_1102; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1104 = 8'h31 == _GEN_99 ? _double_bytes_0_T_17 : _GEN_1103; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1105 = 8'h32 == _GEN_99 ? _double_bytes_0_T_18 : _GEN_1104; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1106 = 8'h33 == _GEN_99 ? _double_bytes_0_T_19 : _GEN_1105; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1107 = 8'h34 == _GEN_99 ? _double_bytes_0_T_20 : _GEN_1106; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1108 = 8'h35 == _GEN_99 ? _double_bytes_0_T_21 : _GEN_1107; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1109 = 8'h36 == _GEN_99 ? _double_bytes_0_T_22 : _GEN_1108; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1110 = 8'h37 == _GEN_99 ? _double_bytes_0_T_23 : _GEN_1109; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1111 = 8'h38 == _GEN_99 ? _double_bytes_0_T_24 : _GEN_1110; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1112 = 8'h39 == _GEN_99 ? _double_bytes_0_T_25 : _GEN_1111; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1113 = 8'h3a == _GEN_99 ? _double_bytes_0_T_26 : _GEN_1112; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1114 = 8'h3b == _GEN_99 ? _double_bytes_0_T_27 : _GEN_1113; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1115 = 8'h3c == _GEN_99 ? _double_bytes_0_T_28 : _GEN_1114; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1116 = 8'h3d == _GEN_99 ? _double_bytes_0_T_29 : _GEN_1115; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1117 = 8'h3e == _GEN_99 ? _double_bytes_0_T_30 : _GEN_1116; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1118 = 8'h3f == _GEN_99 ? _double_bytes_0_T_31 : _GEN_1117; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1119 = 8'h40 == _GEN_99 ? _double_bytes_0_T_32 : _GEN_1118; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1120 = 8'h41 == _GEN_99 ? _double_bytes_0_T_33 : _GEN_1119; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1121 = 8'h42 == _GEN_99 ? _double_bytes_0_T_34 : _GEN_1120; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1122 = 8'h43 == _GEN_99 ? _double_bytes_0_T_35 : _GEN_1121; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1123 = 8'h44 == _GEN_99 ? _double_bytes_0_T_36 : _GEN_1122; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1124 = 8'h45 == _GEN_99 ? _double_bytes_0_T_37 : _GEN_1123; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1125 = 8'h46 == _GEN_99 ? _double_bytes_0_T_38 : _GEN_1124; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1126 = 8'h47 == _GEN_99 ? _double_bytes_0_T_39 : _GEN_1125; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1127 = 8'h48 == _GEN_99 ? _double_bytes_0_T_40 : _GEN_1126; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1128 = 8'h49 == _GEN_99 ? _double_bytes_0_T_41 : _GEN_1127; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1129 = 8'h4a == _GEN_99 ? _double_bytes_0_T_42 : _GEN_1128; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1130 = 8'h4b == _GEN_99 ? _double_bytes_0_T_43 : _GEN_1129; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1131 = 8'h4c == _GEN_99 ? _double_bytes_0_T_44 : _GEN_1130; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1132 = 8'h4d == _GEN_99 ? _double_bytes_0_T_45 : _GEN_1131; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1133 = 8'h4e == _GEN_99 ? _double_bytes_0_T_46 : _GEN_1132; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1134 = 8'h4f == _GEN_99 ? _double_bytes_0_T_47 : _GEN_1133; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] double_bytes_3_1 = _GEN_75 ? _GEN_1134 : 16'h0; // @[matcher_pisa.scala 145:46 matcher_pisa.scala 144:41]
  wire [31:0] _groups_3_T_1 = {double_bytes_3_0,double_bytes_3_1}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_1136 = _GEN_59 == 2'h2 ? _groups_3_T_1 : _GEN_1037; // @[matcher_pisa.scala 139:50 matcher_pisa.scala 153:31]
  wire [31:0] _GEN_1137 = 8'h50 == _GEN_98 ? _groups_0_T_2 : 32'h0; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39 matcher_pisa.scala 158:31]
  wire [31:0] _GEN_1138 = 8'h51 == _GEN_98 ? _groups_0_T_3 : _GEN_1137; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1139 = 8'h52 == _GEN_98 ? _groups_0_T_4 : _GEN_1138; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1140 = 8'h53 == _GEN_98 ? _groups_0_T_5 : _GEN_1139; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1141 = 8'h54 == _GEN_98 ? _groups_0_T_6 : _GEN_1140; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1142 = 8'h55 == _GEN_98 ? _groups_0_T_7 : _GEN_1141; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1143 = 8'h56 == _GEN_98 ? _groups_0_T_8 : _GEN_1142; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1144 = 8'h57 == _GEN_98 ? _groups_0_T_9 : _GEN_1143; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1145 = 8'h58 == _GEN_98 ? _groups_0_T_10 : _GEN_1144; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1146 = 8'h59 == _GEN_98 ? _groups_0_T_11 : _GEN_1145; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1147 = 8'h5a == _GEN_98 ? _groups_0_T_12 : _GEN_1146; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1148 = 8'h5b == _GEN_98 ? _groups_0_T_13 : _GEN_1147; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1149 = 8'h5c == _GEN_98 ? _groups_0_T_14 : _GEN_1148; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1150 = 8'h5d == _GEN_98 ? _groups_0_T_15 : _GEN_1149; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1151 = 8'h5e == _GEN_98 ? _groups_0_T_16 : _GEN_1150; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1152 = 8'h5f == _GEN_98 ? _groups_0_T_17 : _GEN_1151; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1153 = 8'h60 == _GEN_98 ? _groups_0_T_18 : _GEN_1152; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1154 = 8'h61 == _GEN_98 ? _groups_0_T_19 : _GEN_1153; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1155 = 8'h62 == _GEN_98 ? _groups_0_T_20 : _GEN_1154; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1156 = 8'h63 == _GEN_98 ? _groups_0_T_21 : _GEN_1155; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1157 = 8'h64 == _GEN_98 ? _groups_0_T_22 : _GEN_1156; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1158 = 8'h65 == _GEN_98 ? _groups_0_T_23 : _GEN_1157; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1159 = 8'h66 == _GEN_98 ? _groups_0_T_24 : _GEN_1158; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1160 = 8'h67 == _GEN_98 ? _groups_0_T_25 : _GEN_1159; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1161 = 8'h68 == _GEN_98 ? _groups_0_T_26 : _GEN_1160; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1162 = 8'h69 == _GEN_98 ? _groups_0_T_27 : _GEN_1161; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1163 = 8'h6a == _GEN_98 ? _groups_0_T_28 : _GEN_1162; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1164 = 8'h6b == _GEN_98 ? _groups_0_T_29 : _GEN_1163; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1165 = 8'h6c == _GEN_98 ? _groups_0_T_30 : _GEN_1164; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1166 = 8'h6d == _GEN_98 ? _groups_0_T_31 : _GEN_1165; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1167 = 8'h6e == _GEN_98 ? _groups_0_T_32 : _GEN_1166; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1168 = 8'h6f == _GEN_98 ? _groups_0_T_33 : _GEN_1167; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] groups_3 = _GEN_59 == 2'h3 ? _GEN_1168 : _GEN_1136; // @[matcher_pisa.scala 155:50]
  wire [7:0] _GEN_1170 = 8'h0 == _GEN_102 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1171 = 8'h1 == _GEN_102 ? phv_data_1 : _GEN_1170; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1172 = 8'h2 == _GEN_102 ? phv_data_2 : _GEN_1171; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1173 = 8'h3 == _GEN_102 ? phv_data_3 : _GEN_1172; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1174 = 8'h4 == _GEN_102 ? phv_data_4 : _GEN_1173; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1175 = 8'h5 == _GEN_102 ? phv_data_5 : _GEN_1174; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1176 = 8'h6 == _GEN_102 ? phv_data_6 : _GEN_1175; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1177 = 8'h7 == _GEN_102 ? phv_data_7 : _GEN_1176; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1178 = 8'h8 == _GEN_102 ? phv_data_8 : _GEN_1177; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1179 = 8'h9 == _GEN_102 ? phv_data_9 : _GEN_1178; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1180 = 8'ha == _GEN_102 ? phv_data_10 : _GEN_1179; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1181 = 8'hb == _GEN_102 ? phv_data_11 : _GEN_1180; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1182 = 8'hc == _GEN_102 ? phv_data_12 : _GEN_1181; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1183 = 8'hd == _GEN_102 ? phv_data_13 : _GEN_1182; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1184 = 8'he == _GEN_102 ? phv_data_14 : _GEN_1183; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1185 = 8'hf == _GEN_102 ? phv_data_15 : _GEN_1184; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1186 = 8'h10 == _GEN_102 ? phv_data_16 : _GEN_1185; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1187 = 8'h11 == _GEN_102 ? phv_data_17 : _GEN_1186; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1188 = 8'h12 == _GEN_102 ? phv_data_18 : _GEN_1187; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1189 = 8'h13 == _GEN_102 ? phv_data_19 : _GEN_1188; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1190 = 8'h14 == _GEN_102 ? phv_data_20 : _GEN_1189; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1191 = 8'h15 == _GEN_102 ? phv_data_21 : _GEN_1190; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1192 = 8'h16 == _GEN_102 ? phv_data_22 : _GEN_1191; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1193 = 8'h17 == _GEN_102 ? phv_data_23 : _GEN_1192; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1194 = 8'h18 == _GEN_102 ? phv_data_24 : _GEN_1193; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1195 = 8'h19 == _GEN_102 ? phv_data_25 : _GEN_1194; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1196 = 8'h1a == _GEN_102 ? phv_data_26 : _GEN_1195; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1197 = 8'h1b == _GEN_102 ? phv_data_27 : _GEN_1196; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1198 = 8'h1c == _GEN_102 ? phv_data_28 : _GEN_1197; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1199 = 8'h1d == _GEN_102 ? phv_data_29 : _GEN_1198; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1200 = 8'h1e == _GEN_102 ? phv_data_30 : _GEN_1199; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1201 = 8'h1f == _GEN_102 ? phv_data_31 : _GEN_1200; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_4_0 = _GEN_78 ? _GEN_1201 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1203 = 8'h0 == _GEN_103 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1204 = 8'h1 == _GEN_103 ? phv_data_1 : _GEN_1203; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1205 = 8'h2 == _GEN_103 ? phv_data_2 : _GEN_1204; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1206 = 8'h3 == _GEN_103 ? phv_data_3 : _GEN_1205; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1207 = 8'h4 == _GEN_103 ? phv_data_4 : _GEN_1206; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1208 = 8'h5 == _GEN_103 ? phv_data_5 : _GEN_1207; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1209 = 8'h6 == _GEN_103 ? phv_data_6 : _GEN_1208; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1210 = 8'h7 == _GEN_103 ? phv_data_7 : _GEN_1209; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1211 = 8'h8 == _GEN_103 ? phv_data_8 : _GEN_1210; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1212 = 8'h9 == _GEN_103 ? phv_data_9 : _GEN_1211; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1213 = 8'ha == _GEN_103 ? phv_data_10 : _GEN_1212; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1214 = 8'hb == _GEN_103 ? phv_data_11 : _GEN_1213; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1215 = 8'hc == _GEN_103 ? phv_data_12 : _GEN_1214; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1216 = 8'hd == _GEN_103 ? phv_data_13 : _GEN_1215; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1217 = 8'he == _GEN_103 ? phv_data_14 : _GEN_1216; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1218 = 8'hf == _GEN_103 ? phv_data_15 : _GEN_1217; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1219 = 8'h10 == _GEN_103 ? phv_data_16 : _GEN_1218; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1220 = 8'h11 == _GEN_103 ? phv_data_17 : _GEN_1219; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1221 = 8'h12 == _GEN_103 ? phv_data_18 : _GEN_1220; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1222 = 8'h13 == _GEN_103 ? phv_data_19 : _GEN_1221; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1223 = 8'h14 == _GEN_103 ? phv_data_20 : _GEN_1222; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1224 = 8'h15 == _GEN_103 ? phv_data_21 : _GEN_1223; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1225 = 8'h16 == _GEN_103 ? phv_data_22 : _GEN_1224; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1226 = 8'h17 == _GEN_103 ? phv_data_23 : _GEN_1225; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1227 = 8'h18 == _GEN_103 ? phv_data_24 : _GEN_1226; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1228 = 8'h19 == _GEN_103 ? phv_data_25 : _GEN_1227; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1229 = 8'h1a == _GEN_103 ? phv_data_26 : _GEN_1228; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1230 = 8'h1b == _GEN_103 ? phv_data_27 : _GEN_1229; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1231 = 8'h1c == _GEN_103 ? phv_data_28 : _GEN_1230; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1232 = 8'h1d == _GEN_103 ? phv_data_29 : _GEN_1231; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1233 = 8'h1e == _GEN_103 ? phv_data_30 : _GEN_1232; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1234 = 8'h1f == _GEN_103 ? phv_data_31 : _GEN_1233; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_4_1 = _GEN_79 ? _GEN_1234 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1236 = 8'h0 == _GEN_104 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1237 = 8'h1 == _GEN_104 ? phv_data_1 : _GEN_1236; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1238 = 8'h2 == _GEN_104 ? phv_data_2 : _GEN_1237; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1239 = 8'h3 == _GEN_104 ? phv_data_3 : _GEN_1238; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1240 = 8'h4 == _GEN_104 ? phv_data_4 : _GEN_1239; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1241 = 8'h5 == _GEN_104 ? phv_data_5 : _GEN_1240; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1242 = 8'h6 == _GEN_104 ? phv_data_6 : _GEN_1241; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1243 = 8'h7 == _GEN_104 ? phv_data_7 : _GEN_1242; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1244 = 8'h8 == _GEN_104 ? phv_data_8 : _GEN_1243; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1245 = 8'h9 == _GEN_104 ? phv_data_9 : _GEN_1244; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1246 = 8'ha == _GEN_104 ? phv_data_10 : _GEN_1245; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1247 = 8'hb == _GEN_104 ? phv_data_11 : _GEN_1246; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1248 = 8'hc == _GEN_104 ? phv_data_12 : _GEN_1247; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1249 = 8'hd == _GEN_104 ? phv_data_13 : _GEN_1248; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1250 = 8'he == _GEN_104 ? phv_data_14 : _GEN_1249; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1251 = 8'hf == _GEN_104 ? phv_data_15 : _GEN_1250; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1252 = 8'h10 == _GEN_104 ? phv_data_16 : _GEN_1251; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1253 = 8'h11 == _GEN_104 ? phv_data_17 : _GEN_1252; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1254 = 8'h12 == _GEN_104 ? phv_data_18 : _GEN_1253; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1255 = 8'h13 == _GEN_104 ? phv_data_19 : _GEN_1254; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1256 = 8'h14 == _GEN_104 ? phv_data_20 : _GEN_1255; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1257 = 8'h15 == _GEN_104 ? phv_data_21 : _GEN_1256; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1258 = 8'h16 == _GEN_104 ? phv_data_22 : _GEN_1257; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1259 = 8'h17 == _GEN_104 ? phv_data_23 : _GEN_1258; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1260 = 8'h18 == _GEN_104 ? phv_data_24 : _GEN_1259; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1261 = 8'h19 == _GEN_104 ? phv_data_25 : _GEN_1260; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1262 = 8'h1a == _GEN_104 ? phv_data_26 : _GEN_1261; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1263 = 8'h1b == _GEN_104 ? phv_data_27 : _GEN_1262; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1264 = 8'h1c == _GEN_104 ? phv_data_28 : _GEN_1263; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1265 = 8'h1d == _GEN_104 ? phv_data_29 : _GEN_1264; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1266 = 8'h1e == _GEN_104 ? phv_data_30 : _GEN_1265; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1267 = 8'h1f == _GEN_104 ? phv_data_31 : _GEN_1266; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_4_2 = _GEN_80 ? _GEN_1267 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1269 = 8'h0 == _GEN_105 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1270 = 8'h1 == _GEN_105 ? phv_data_1 : _GEN_1269; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1271 = 8'h2 == _GEN_105 ? phv_data_2 : _GEN_1270; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1272 = 8'h3 == _GEN_105 ? phv_data_3 : _GEN_1271; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1273 = 8'h4 == _GEN_105 ? phv_data_4 : _GEN_1272; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1274 = 8'h5 == _GEN_105 ? phv_data_5 : _GEN_1273; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1275 = 8'h6 == _GEN_105 ? phv_data_6 : _GEN_1274; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1276 = 8'h7 == _GEN_105 ? phv_data_7 : _GEN_1275; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1277 = 8'h8 == _GEN_105 ? phv_data_8 : _GEN_1276; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1278 = 8'h9 == _GEN_105 ? phv_data_9 : _GEN_1277; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1279 = 8'ha == _GEN_105 ? phv_data_10 : _GEN_1278; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1280 = 8'hb == _GEN_105 ? phv_data_11 : _GEN_1279; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1281 = 8'hc == _GEN_105 ? phv_data_12 : _GEN_1280; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1282 = 8'hd == _GEN_105 ? phv_data_13 : _GEN_1281; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1283 = 8'he == _GEN_105 ? phv_data_14 : _GEN_1282; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1284 = 8'hf == _GEN_105 ? phv_data_15 : _GEN_1283; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1285 = 8'h10 == _GEN_105 ? phv_data_16 : _GEN_1284; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1286 = 8'h11 == _GEN_105 ? phv_data_17 : _GEN_1285; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1287 = 8'h12 == _GEN_105 ? phv_data_18 : _GEN_1286; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1288 = 8'h13 == _GEN_105 ? phv_data_19 : _GEN_1287; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1289 = 8'h14 == _GEN_105 ? phv_data_20 : _GEN_1288; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1290 = 8'h15 == _GEN_105 ? phv_data_21 : _GEN_1289; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1291 = 8'h16 == _GEN_105 ? phv_data_22 : _GEN_1290; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1292 = 8'h17 == _GEN_105 ? phv_data_23 : _GEN_1291; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1293 = 8'h18 == _GEN_105 ? phv_data_24 : _GEN_1292; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1294 = 8'h19 == _GEN_105 ? phv_data_25 : _GEN_1293; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1295 = 8'h1a == _GEN_105 ? phv_data_26 : _GEN_1294; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1296 = 8'h1b == _GEN_105 ? phv_data_27 : _GEN_1295; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1297 = 8'h1c == _GEN_105 ? phv_data_28 : _GEN_1296; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1298 = 8'h1d == _GEN_105 ? phv_data_29 : _GEN_1297; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1299 = 8'h1e == _GEN_105 ? phv_data_30 : _GEN_1298; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1300 = 8'h1f == _GEN_105 ? phv_data_31 : _GEN_1299; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_4_3 = _GEN_81 ? _GEN_1300 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [31:0] _groups_4_T = {bytes_4_0,bytes_4_1,bytes_4_2,bytes_4_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_1302 = _GEN_60 == 2'h1 ? _groups_4_T : 32'h0; // @[matcher_pisa.scala 123:50 matcher_pisa.scala 137:31 matcher_pisa.scala 122:27]
  wire [15:0] _GEN_1303 = 8'h20 == _GEN_102 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_1304 = 8'h21 == _GEN_102 ? _double_bytes_0_T_1 : _GEN_1303; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1305 = 8'h22 == _GEN_102 ? _double_bytes_0_T_2 : _GEN_1304; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1306 = 8'h23 == _GEN_102 ? _double_bytes_0_T_3 : _GEN_1305; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1307 = 8'h24 == _GEN_102 ? _double_bytes_0_T_4 : _GEN_1306; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1308 = 8'h25 == _GEN_102 ? _double_bytes_0_T_5 : _GEN_1307; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1309 = 8'h26 == _GEN_102 ? _double_bytes_0_T_6 : _GEN_1308; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1310 = 8'h27 == _GEN_102 ? _double_bytes_0_T_7 : _GEN_1309; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1311 = 8'h28 == _GEN_102 ? _double_bytes_0_T_8 : _GEN_1310; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1312 = 8'h29 == _GEN_102 ? _double_bytes_0_T_9 : _GEN_1311; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1313 = 8'h2a == _GEN_102 ? _double_bytes_0_T_10 : _GEN_1312; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1314 = 8'h2b == _GEN_102 ? _double_bytes_0_T_11 : _GEN_1313; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1315 = 8'h2c == _GEN_102 ? _double_bytes_0_T_12 : _GEN_1314; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1316 = 8'h2d == _GEN_102 ? _double_bytes_0_T_13 : _GEN_1315; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1317 = 8'h2e == _GEN_102 ? _double_bytes_0_T_14 : _GEN_1316; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1318 = 8'h2f == _GEN_102 ? _double_bytes_0_T_15 : _GEN_1317; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1319 = 8'h30 == _GEN_102 ? _double_bytes_0_T_16 : _GEN_1318; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1320 = 8'h31 == _GEN_102 ? _double_bytes_0_T_17 : _GEN_1319; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1321 = 8'h32 == _GEN_102 ? _double_bytes_0_T_18 : _GEN_1320; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1322 = 8'h33 == _GEN_102 ? _double_bytes_0_T_19 : _GEN_1321; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1323 = 8'h34 == _GEN_102 ? _double_bytes_0_T_20 : _GEN_1322; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1324 = 8'h35 == _GEN_102 ? _double_bytes_0_T_21 : _GEN_1323; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1325 = 8'h36 == _GEN_102 ? _double_bytes_0_T_22 : _GEN_1324; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1326 = 8'h37 == _GEN_102 ? _double_bytes_0_T_23 : _GEN_1325; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1327 = 8'h38 == _GEN_102 ? _double_bytes_0_T_24 : _GEN_1326; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1328 = 8'h39 == _GEN_102 ? _double_bytes_0_T_25 : _GEN_1327; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1329 = 8'h3a == _GEN_102 ? _double_bytes_0_T_26 : _GEN_1328; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1330 = 8'h3b == _GEN_102 ? _double_bytes_0_T_27 : _GEN_1329; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1331 = 8'h3c == _GEN_102 ? _double_bytes_0_T_28 : _GEN_1330; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1332 = 8'h3d == _GEN_102 ? _double_bytes_0_T_29 : _GEN_1331; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1333 = 8'h3e == _GEN_102 ? _double_bytes_0_T_30 : _GEN_1332; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1334 = 8'h3f == _GEN_102 ? _double_bytes_0_T_31 : _GEN_1333; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1335 = 8'h40 == _GEN_102 ? _double_bytes_0_T_32 : _GEN_1334; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1336 = 8'h41 == _GEN_102 ? _double_bytes_0_T_33 : _GEN_1335; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1337 = 8'h42 == _GEN_102 ? _double_bytes_0_T_34 : _GEN_1336; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1338 = 8'h43 == _GEN_102 ? _double_bytes_0_T_35 : _GEN_1337; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1339 = 8'h44 == _GEN_102 ? _double_bytes_0_T_36 : _GEN_1338; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1340 = 8'h45 == _GEN_102 ? _double_bytes_0_T_37 : _GEN_1339; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1341 = 8'h46 == _GEN_102 ? _double_bytes_0_T_38 : _GEN_1340; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1342 = 8'h47 == _GEN_102 ? _double_bytes_0_T_39 : _GEN_1341; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1343 = 8'h48 == _GEN_102 ? _double_bytes_0_T_40 : _GEN_1342; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1344 = 8'h49 == _GEN_102 ? _double_bytes_0_T_41 : _GEN_1343; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1345 = 8'h4a == _GEN_102 ? _double_bytes_0_T_42 : _GEN_1344; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1346 = 8'h4b == _GEN_102 ? _double_bytes_0_T_43 : _GEN_1345; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1347 = 8'h4c == _GEN_102 ? _double_bytes_0_T_44 : _GEN_1346; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1348 = 8'h4d == _GEN_102 ? _double_bytes_0_T_45 : _GEN_1347; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1349 = 8'h4e == _GEN_102 ? _double_bytes_0_T_46 : _GEN_1348; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1350 = 8'h4f == _GEN_102 ? _double_bytes_0_T_47 : _GEN_1349; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] double_bytes_4_0 = _GEN_78 ? _GEN_1350 : 16'h0; // @[matcher_pisa.scala 145:46 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_1352 = 8'h20 == _GEN_103 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_1353 = 8'h21 == _GEN_103 ? _double_bytes_0_T_1 : _GEN_1352; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1354 = 8'h22 == _GEN_103 ? _double_bytes_0_T_2 : _GEN_1353; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1355 = 8'h23 == _GEN_103 ? _double_bytes_0_T_3 : _GEN_1354; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1356 = 8'h24 == _GEN_103 ? _double_bytes_0_T_4 : _GEN_1355; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1357 = 8'h25 == _GEN_103 ? _double_bytes_0_T_5 : _GEN_1356; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1358 = 8'h26 == _GEN_103 ? _double_bytes_0_T_6 : _GEN_1357; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1359 = 8'h27 == _GEN_103 ? _double_bytes_0_T_7 : _GEN_1358; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1360 = 8'h28 == _GEN_103 ? _double_bytes_0_T_8 : _GEN_1359; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1361 = 8'h29 == _GEN_103 ? _double_bytes_0_T_9 : _GEN_1360; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1362 = 8'h2a == _GEN_103 ? _double_bytes_0_T_10 : _GEN_1361; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1363 = 8'h2b == _GEN_103 ? _double_bytes_0_T_11 : _GEN_1362; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1364 = 8'h2c == _GEN_103 ? _double_bytes_0_T_12 : _GEN_1363; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1365 = 8'h2d == _GEN_103 ? _double_bytes_0_T_13 : _GEN_1364; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1366 = 8'h2e == _GEN_103 ? _double_bytes_0_T_14 : _GEN_1365; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1367 = 8'h2f == _GEN_103 ? _double_bytes_0_T_15 : _GEN_1366; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1368 = 8'h30 == _GEN_103 ? _double_bytes_0_T_16 : _GEN_1367; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1369 = 8'h31 == _GEN_103 ? _double_bytes_0_T_17 : _GEN_1368; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1370 = 8'h32 == _GEN_103 ? _double_bytes_0_T_18 : _GEN_1369; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1371 = 8'h33 == _GEN_103 ? _double_bytes_0_T_19 : _GEN_1370; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1372 = 8'h34 == _GEN_103 ? _double_bytes_0_T_20 : _GEN_1371; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1373 = 8'h35 == _GEN_103 ? _double_bytes_0_T_21 : _GEN_1372; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1374 = 8'h36 == _GEN_103 ? _double_bytes_0_T_22 : _GEN_1373; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1375 = 8'h37 == _GEN_103 ? _double_bytes_0_T_23 : _GEN_1374; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1376 = 8'h38 == _GEN_103 ? _double_bytes_0_T_24 : _GEN_1375; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1377 = 8'h39 == _GEN_103 ? _double_bytes_0_T_25 : _GEN_1376; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1378 = 8'h3a == _GEN_103 ? _double_bytes_0_T_26 : _GEN_1377; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1379 = 8'h3b == _GEN_103 ? _double_bytes_0_T_27 : _GEN_1378; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1380 = 8'h3c == _GEN_103 ? _double_bytes_0_T_28 : _GEN_1379; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1381 = 8'h3d == _GEN_103 ? _double_bytes_0_T_29 : _GEN_1380; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1382 = 8'h3e == _GEN_103 ? _double_bytes_0_T_30 : _GEN_1381; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1383 = 8'h3f == _GEN_103 ? _double_bytes_0_T_31 : _GEN_1382; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1384 = 8'h40 == _GEN_103 ? _double_bytes_0_T_32 : _GEN_1383; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1385 = 8'h41 == _GEN_103 ? _double_bytes_0_T_33 : _GEN_1384; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1386 = 8'h42 == _GEN_103 ? _double_bytes_0_T_34 : _GEN_1385; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1387 = 8'h43 == _GEN_103 ? _double_bytes_0_T_35 : _GEN_1386; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1388 = 8'h44 == _GEN_103 ? _double_bytes_0_T_36 : _GEN_1387; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1389 = 8'h45 == _GEN_103 ? _double_bytes_0_T_37 : _GEN_1388; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1390 = 8'h46 == _GEN_103 ? _double_bytes_0_T_38 : _GEN_1389; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1391 = 8'h47 == _GEN_103 ? _double_bytes_0_T_39 : _GEN_1390; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1392 = 8'h48 == _GEN_103 ? _double_bytes_0_T_40 : _GEN_1391; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1393 = 8'h49 == _GEN_103 ? _double_bytes_0_T_41 : _GEN_1392; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1394 = 8'h4a == _GEN_103 ? _double_bytes_0_T_42 : _GEN_1393; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1395 = 8'h4b == _GEN_103 ? _double_bytes_0_T_43 : _GEN_1394; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1396 = 8'h4c == _GEN_103 ? _double_bytes_0_T_44 : _GEN_1395; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1397 = 8'h4d == _GEN_103 ? _double_bytes_0_T_45 : _GEN_1396; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1398 = 8'h4e == _GEN_103 ? _double_bytes_0_T_46 : _GEN_1397; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1399 = 8'h4f == _GEN_103 ? _double_bytes_0_T_47 : _GEN_1398; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] double_bytes_4_1 = _GEN_79 ? _GEN_1399 : 16'h0; // @[matcher_pisa.scala 145:46 matcher_pisa.scala 144:41]
  wire [31:0] _groups_4_T_1 = {double_bytes_4_0,double_bytes_4_1}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_1401 = _GEN_60 == 2'h2 ? _groups_4_T_1 : _GEN_1302; // @[matcher_pisa.scala 139:50 matcher_pisa.scala 153:31]
  wire [31:0] _GEN_1402 = 8'h50 == _GEN_102 ? _groups_0_T_2 : 32'h0; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39 matcher_pisa.scala 158:31]
  wire [31:0] _GEN_1403 = 8'h51 == _GEN_102 ? _groups_0_T_3 : _GEN_1402; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1404 = 8'h52 == _GEN_102 ? _groups_0_T_4 : _GEN_1403; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1405 = 8'h53 == _GEN_102 ? _groups_0_T_5 : _GEN_1404; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1406 = 8'h54 == _GEN_102 ? _groups_0_T_6 : _GEN_1405; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1407 = 8'h55 == _GEN_102 ? _groups_0_T_7 : _GEN_1406; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1408 = 8'h56 == _GEN_102 ? _groups_0_T_8 : _GEN_1407; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1409 = 8'h57 == _GEN_102 ? _groups_0_T_9 : _GEN_1408; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1410 = 8'h58 == _GEN_102 ? _groups_0_T_10 : _GEN_1409; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1411 = 8'h59 == _GEN_102 ? _groups_0_T_11 : _GEN_1410; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1412 = 8'h5a == _GEN_102 ? _groups_0_T_12 : _GEN_1411; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1413 = 8'h5b == _GEN_102 ? _groups_0_T_13 : _GEN_1412; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1414 = 8'h5c == _GEN_102 ? _groups_0_T_14 : _GEN_1413; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1415 = 8'h5d == _GEN_102 ? _groups_0_T_15 : _GEN_1414; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1416 = 8'h5e == _GEN_102 ? _groups_0_T_16 : _GEN_1415; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1417 = 8'h5f == _GEN_102 ? _groups_0_T_17 : _GEN_1416; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1418 = 8'h60 == _GEN_102 ? _groups_0_T_18 : _GEN_1417; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1419 = 8'h61 == _GEN_102 ? _groups_0_T_19 : _GEN_1418; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1420 = 8'h62 == _GEN_102 ? _groups_0_T_20 : _GEN_1419; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1421 = 8'h63 == _GEN_102 ? _groups_0_T_21 : _GEN_1420; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1422 = 8'h64 == _GEN_102 ? _groups_0_T_22 : _GEN_1421; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1423 = 8'h65 == _GEN_102 ? _groups_0_T_23 : _GEN_1422; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1424 = 8'h66 == _GEN_102 ? _groups_0_T_24 : _GEN_1423; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1425 = 8'h67 == _GEN_102 ? _groups_0_T_25 : _GEN_1424; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1426 = 8'h68 == _GEN_102 ? _groups_0_T_26 : _GEN_1425; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1427 = 8'h69 == _GEN_102 ? _groups_0_T_27 : _GEN_1426; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1428 = 8'h6a == _GEN_102 ? _groups_0_T_28 : _GEN_1427; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1429 = 8'h6b == _GEN_102 ? _groups_0_T_29 : _GEN_1428; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1430 = 8'h6c == _GEN_102 ? _groups_0_T_30 : _GEN_1429; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1431 = 8'h6d == _GEN_102 ? _groups_0_T_31 : _GEN_1430; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1432 = 8'h6e == _GEN_102 ? _groups_0_T_32 : _GEN_1431; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1433 = 8'h6f == _GEN_102 ? _groups_0_T_33 : _GEN_1432; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] groups_4 = _GEN_60 == 2'h3 ? _GEN_1433 : _GEN_1401; // @[matcher_pisa.scala 155:50]
  wire [7:0] _GEN_1435 = 8'h0 == _GEN_106 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1436 = 8'h1 == _GEN_106 ? phv_data_1 : _GEN_1435; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1437 = 8'h2 == _GEN_106 ? phv_data_2 : _GEN_1436; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1438 = 8'h3 == _GEN_106 ? phv_data_3 : _GEN_1437; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1439 = 8'h4 == _GEN_106 ? phv_data_4 : _GEN_1438; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1440 = 8'h5 == _GEN_106 ? phv_data_5 : _GEN_1439; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1441 = 8'h6 == _GEN_106 ? phv_data_6 : _GEN_1440; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1442 = 8'h7 == _GEN_106 ? phv_data_7 : _GEN_1441; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1443 = 8'h8 == _GEN_106 ? phv_data_8 : _GEN_1442; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1444 = 8'h9 == _GEN_106 ? phv_data_9 : _GEN_1443; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1445 = 8'ha == _GEN_106 ? phv_data_10 : _GEN_1444; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1446 = 8'hb == _GEN_106 ? phv_data_11 : _GEN_1445; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1447 = 8'hc == _GEN_106 ? phv_data_12 : _GEN_1446; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1448 = 8'hd == _GEN_106 ? phv_data_13 : _GEN_1447; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1449 = 8'he == _GEN_106 ? phv_data_14 : _GEN_1448; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1450 = 8'hf == _GEN_106 ? phv_data_15 : _GEN_1449; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1451 = 8'h10 == _GEN_106 ? phv_data_16 : _GEN_1450; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1452 = 8'h11 == _GEN_106 ? phv_data_17 : _GEN_1451; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1453 = 8'h12 == _GEN_106 ? phv_data_18 : _GEN_1452; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1454 = 8'h13 == _GEN_106 ? phv_data_19 : _GEN_1453; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1455 = 8'h14 == _GEN_106 ? phv_data_20 : _GEN_1454; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1456 = 8'h15 == _GEN_106 ? phv_data_21 : _GEN_1455; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1457 = 8'h16 == _GEN_106 ? phv_data_22 : _GEN_1456; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1458 = 8'h17 == _GEN_106 ? phv_data_23 : _GEN_1457; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1459 = 8'h18 == _GEN_106 ? phv_data_24 : _GEN_1458; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1460 = 8'h19 == _GEN_106 ? phv_data_25 : _GEN_1459; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1461 = 8'h1a == _GEN_106 ? phv_data_26 : _GEN_1460; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1462 = 8'h1b == _GEN_106 ? phv_data_27 : _GEN_1461; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1463 = 8'h1c == _GEN_106 ? phv_data_28 : _GEN_1462; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1464 = 8'h1d == _GEN_106 ? phv_data_29 : _GEN_1463; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1465 = 8'h1e == _GEN_106 ? phv_data_30 : _GEN_1464; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1466 = 8'h1f == _GEN_106 ? phv_data_31 : _GEN_1465; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_5_0 = _GEN_82 ? _GEN_1466 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1468 = 8'h0 == _GEN_107 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1469 = 8'h1 == _GEN_107 ? phv_data_1 : _GEN_1468; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1470 = 8'h2 == _GEN_107 ? phv_data_2 : _GEN_1469; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1471 = 8'h3 == _GEN_107 ? phv_data_3 : _GEN_1470; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1472 = 8'h4 == _GEN_107 ? phv_data_4 : _GEN_1471; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1473 = 8'h5 == _GEN_107 ? phv_data_5 : _GEN_1472; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1474 = 8'h6 == _GEN_107 ? phv_data_6 : _GEN_1473; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1475 = 8'h7 == _GEN_107 ? phv_data_7 : _GEN_1474; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1476 = 8'h8 == _GEN_107 ? phv_data_8 : _GEN_1475; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1477 = 8'h9 == _GEN_107 ? phv_data_9 : _GEN_1476; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1478 = 8'ha == _GEN_107 ? phv_data_10 : _GEN_1477; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1479 = 8'hb == _GEN_107 ? phv_data_11 : _GEN_1478; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1480 = 8'hc == _GEN_107 ? phv_data_12 : _GEN_1479; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1481 = 8'hd == _GEN_107 ? phv_data_13 : _GEN_1480; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1482 = 8'he == _GEN_107 ? phv_data_14 : _GEN_1481; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1483 = 8'hf == _GEN_107 ? phv_data_15 : _GEN_1482; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1484 = 8'h10 == _GEN_107 ? phv_data_16 : _GEN_1483; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1485 = 8'h11 == _GEN_107 ? phv_data_17 : _GEN_1484; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1486 = 8'h12 == _GEN_107 ? phv_data_18 : _GEN_1485; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1487 = 8'h13 == _GEN_107 ? phv_data_19 : _GEN_1486; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1488 = 8'h14 == _GEN_107 ? phv_data_20 : _GEN_1487; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1489 = 8'h15 == _GEN_107 ? phv_data_21 : _GEN_1488; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1490 = 8'h16 == _GEN_107 ? phv_data_22 : _GEN_1489; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1491 = 8'h17 == _GEN_107 ? phv_data_23 : _GEN_1490; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1492 = 8'h18 == _GEN_107 ? phv_data_24 : _GEN_1491; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1493 = 8'h19 == _GEN_107 ? phv_data_25 : _GEN_1492; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1494 = 8'h1a == _GEN_107 ? phv_data_26 : _GEN_1493; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1495 = 8'h1b == _GEN_107 ? phv_data_27 : _GEN_1494; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1496 = 8'h1c == _GEN_107 ? phv_data_28 : _GEN_1495; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1497 = 8'h1d == _GEN_107 ? phv_data_29 : _GEN_1496; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1498 = 8'h1e == _GEN_107 ? phv_data_30 : _GEN_1497; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1499 = 8'h1f == _GEN_107 ? phv_data_31 : _GEN_1498; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_5_1 = _GEN_83 ? _GEN_1499 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1501 = 8'h0 == _GEN_108 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1502 = 8'h1 == _GEN_108 ? phv_data_1 : _GEN_1501; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1503 = 8'h2 == _GEN_108 ? phv_data_2 : _GEN_1502; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1504 = 8'h3 == _GEN_108 ? phv_data_3 : _GEN_1503; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1505 = 8'h4 == _GEN_108 ? phv_data_4 : _GEN_1504; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1506 = 8'h5 == _GEN_108 ? phv_data_5 : _GEN_1505; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1507 = 8'h6 == _GEN_108 ? phv_data_6 : _GEN_1506; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1508 = 8'h7 == _GEN_108 ? phv_data_7 : _GEN_1507; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1509 = 8'h8 == _GEN_108 ? phv_data_8 : _GEN_1508; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1510 = 8'h9 == _GEN_108 ? phv_data_9 : _GEN_1509; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1511 = 8'ha == _GEN_108 ? phv_data_10 : _GEN_1510; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1512 = 8'hb == _GEN_108 ? phv_data_11 : _GEN_1511; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1513 = 8'hc == _GEN_108 ? phv_data_12 : _GEN_1512; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1514 = 8'hd == _GEN_108 ? phv_data_13 : _GEN_1513; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1515 = 8'he == _GEN_108 ? phv_data_14 : _GEN_1514; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1516 = 8'hf == _GEN_108 ? phv_data_15 : _GEN_1515; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1517 = 8'h10 == _GEN_108 ? phv_data_16 : _GEN_1516; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1518 = 8'h11 == _GEN_108 ? phv_data_17 : _GEN_1517; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1519 = 8'h12 == _GEN_108 ? phv_data_18 : _GEN_1518; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1520 = 8'h13 == _GEN_108 ? phv_data_19 : _GEN_1519; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1521 = 8'h14 == _GEN_108 ? phv_data_20 : _GEN_1520; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1522 = 8'h15 == _GEN_108 ? phv_data_21 : _GEN_1521; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1523 = 8'h16 == _GEN_108 ? phv_data_22 : _GEN_1522; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1524 = 8'h17 == _GEN_108 ? phv_data_23 : _GEN_1523; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1525 = 8'h18 == _GEN_108 ? phv_data_24 : _GEN_1524; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1526 = 8'h19 == _GEN_108 ? phv_data_25 : _GEN_1525; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1527 = 8'h1a == _GEN_108 ? phv_data_26 : _GEN_1526; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1528 = 8'h1b == _GEN_108 ? phv_data_27 : _GEN_1527; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1529 = 8'h1c == _GEN_108 ? phv_data_28 : _GEN_1528; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1530 = 8'h1d == _GEN_108 ? phv_data_29 : _GEN_1529; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1531 = 8'h1e == _GEN_108 ? phv_data_30 : _GEN_1530; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1532 = 8'h1f == _GEN_108 ? phv_data_31 : _GEN_1531; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_5_2 = _GEN_84 ? _GEN_1532 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1534 = 8'h0 == _GEN_109 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46 matcher_pisa.scala 128:34]
  wire [7:0] _GEN_1535 = 8'h1 == _GEN_109 ? phv_data_1 : _GEN_1534; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1536 = 8'h2 == _GEN_109 ? phv_data_2 : _GEN_1535; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1537 = 8'h3 == _GEN_109 ? phv_data_3 : _GEN_1536; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1538 = 8'h4 == _GEN_109 ? phv_data_4 : _GEN_1537; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1539 = 8'h5 == _GEN_109 ? phv_data_5 : _GEN_1538; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1540 = 8'h6 == _GEN_109 ? phv_data_6 : _GEN_1539; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1541 = 8'h7 == _GEN_109 ? phv_data_7 : _GEN_1540; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1542 = 8'h8 == _GEN_109 ? phv_data_8 : _GEN_1541; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1543 = 8'h9 == _GEN_109 ? phv_data_9 : _GEN_1542; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1544 = 8'ha == _GEN_109 ? phv_data_10 : _GEN_1543; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1545 = 8'hb == _GEN_109 ? phv_data_11 : _GEN_1544; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1546 = 8'hc == _GEN_109 ? phv_data_12 : _GEN_1545; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1547 = 8'hd == _GEN_109 ? phv_data_13 : _GEN_1546; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1548 = 8'he == _GEN_109 ? phv_data_14 : _GEN_1547; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1549 = 8'hf == _GEN_109 ? phv_data_15 : _GEN_1548; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1550 = 8'h10 == _GEN_109 ? phv_data_16 : _GEN_1549; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1551 = 8'h11 == _GEN_109 ? phv_data_17 : _GEN_1550; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1552 = 8'h12 == _GEN_109 ? phv_data_18 : _GEN_1551; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1553 = 8'h13 == _GEN_109 ? phv_data_19 : _GEN_1552; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1554 = 8'h14 == _GEN_109 ? phv_data_20 : _GEN_1553; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1555 = 8'h15 == _GEN_109 ? phv_data_21 : _GEN_1554; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1556 = 8'h16 == _GEN_109 ? phv_data_22 : _GEN_1555; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1557 = 8'h17 == _GEN_109 ? phv_data_23 : _GEN_1556; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1558 = 8'h18 == _GEN_109 ? phv_data_24 : _GEN_1557; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1559 = 8'h19 == _GEN_109 ? phv_data_25 : _GEN_1558; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1560 = 8'h1a == _GEN_109 ? phv_data_26 : _GEN_1559; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1561 = 8'h1b == _GEN_109 ? phv_data_27 : _GEN_1560; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1562 = 8'h1c == _GEN_109 ? phv_data_28 : _GEN_1561; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1563 = 8'h1d == _GEN_109 ? phv_data_29 : _GEN_1562; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1564 = 8'h1e == _GEN_109 ? phv_data_30 : _GEN_1563; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] _GEN_1565 = 8'h1f == _GEN_109 ? phv_data_31 : _GEN_1564; // @[matcher_pisa.scala 131:85 matcher_pisa.scala 132:46]
  wire [7:0] bytes_5_3 = _GEN_85 ? _GEN_1565 : 8'h0; // @[matcher_pisa.scala 129:46 matcher_pisa.scala 128:34]
  wire [31:0] _groups_5_T = {bytes_5_0,bytes_5_1,bytes_5_2,bytes_5_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_1567 = _GEN_61 == 2'h1 ? _groups_5_T : 32'h0; // @[matcher_pisa.scala 123:50 matcher_pisa.scala 137:31 matcher_pisa.scala 122:27]
  wire [15:0] _GEN_1568 = 8'h20 == _GEN_106 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_1569 = 8'h21 == _GEN_106 ? _double_bytes_0_T_1 : _GEN_1568; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1570 = 8'h22 == _GEN_106 ? _double_bytes_0_T_2 : _GEN_1569; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1571 = 8'h23 == _GEN_106 ? _double_bytes_0_T_3 : _GEN_1570; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1572 = 8'h24 == _GEN_106 ? _double_bytes_0_T_4 : _GEN_1571; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1573 = 8'h25 == _GEN_106 ? _double_bytes_0_T_5 : _GEN_1572; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1574 = 8'h26 == _GEN_106 ? _double_bytes_0_T_6 : _GEN_1573; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1575 = 8'h27 == _GEN_106 ? _double_bytes_0_T_7 : _GEN_1574; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1576 = 8'h28 == _GEN_106 ? _double_bytes_0_T_8 : _GEN_1575; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1577 = 8'h29 == _GEN_106 ? _double_bytes_0_T_9 : _GEN_1576; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1578 = 8'h2a == _GEN_106 ? _double_bytes_0_T_10 : _GEN_1577; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1579 = 8'h2b == _GEN_106 ? _double_bytes_0_T_11 : _GEN_1578; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1580 = 8'h2c == _GEN_106 ? _double_bytes_0_T_12 : _GEN_1579; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1581 = 8'h2d == _GEN_106 ? _double_bytes_0_T_13 : _GEN_1580; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1582 = 8'h2e == _GEN_106 ? _double_bytes_0_T_14 : _GEN_1581; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1583 = 8'h2f == _GEN_106 ? _double_bytes_0_T_15 : _GEN_1582; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1584 = 8'h30 == _GEN_106 ? _double_bytes_0_T_16 : _GEN_1583; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1585 = 8'h31 == _GEN_106 ? _double_bytes_0_T_17 : _GEN_1584; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1586 = 8'h32 == _GEN_106 ? _double_bytes_0_T_18 : _GEN_1585; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1587 = 8'h33 == _GEN_106 ? _double_bytes_0_T_19 : _GEN_1586; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1588 = 8'h34 == _GEN_106 ? _double_bytes_0_T_20 : _GEN_1587; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1589 = 8'h35 == _GEN_106 ? _double_bytes_0_T_21 : _GEN_1588; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1590 = 8'h36 == _GEN_106 ? _double_bytes_0_T_22 : _GEN_1589; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1591 = 8'h37 == _GEN_106 ? _double_bytes_0_T_23 : _GEN_1590; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1592 = 8'h38 == _GEN_106 ? _double_bytes_0_T_24 : _GEN_1591; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1593 = 8'h39 == _GEN_106 ? _double_bytes_0_T_25 : _GEN_1592; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1594 = 8'h3a == _GEN_106 ? _double_bytes_0_T_26 : _GEN_1593; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1595 = 8'h3b == _GEN_106 ? _double_bytes_0_T_27 : _GEN_1594; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1596 = 8'h3c == _GEN_106 ? _double_bytes_0_T_28 : _GEN_1595; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1597 = 8'h3d == _GEN_106 ? _double_bytes_0_T_29 : _GEN_1596; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1598 = 8'h3e == _GEN_106 ? _double_bytes_0_T_30 : _GEN_1597; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1599 = 8'h3f == _GEN_106 ? _double_bytes_0_T_31 : _GEN_1598; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1600 = 8'h40 == _GEN_106 ? _double_bytes_0_T_32 : _GEN_1599; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1601 = 8'h41 == _GEN_106 ? _double_bytes_0_T_33 : _GEN_1600; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1602 = 8'h42 == _GEN_106 ? _double_bytes_0_T_34 : _GEN_1601; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1603 = 8'h43 == _GEN_106 ? _double_bytes_0_T_35 : _GEN_1602; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1604 = 8'h44 == _GEN_106 ? _double_bytes_0_T_36 : _GEN_1603; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1605 = 8'h45 == _GEN_106 ? _double_bytes_0_T_37 : _GEN_1604; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1606 = 8'h46 == _GEN_106 ? _double_bytes_0_T_38 : _GEN_1605; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1607 = 8'h47 == _GEN_106 ? _double_bytes_0_T_39 : _GEN_1606; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1608 = 8'h48 == _GEN_106 ? _double_bytes_0_T_40 : _GEN_1607; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1609 = 8'h49 == _GEN_106 ? _double_bytes_0_T_41 : _GEN_1608; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1610 = 8'h4a == _GEN_106 ? _double_bytes_0_T_42 : _GEN_1609; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1611 = 8'h4b == _GEN_106 ? _double_bytes_0_T_43 : _GEN_1610; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1612 = 8'h4c == _GEN_106 ? _double_bytes_0_T_44 : _GEN_1611; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1613 = 8'h4d == _GEN_106 ? _double_bytes_0_T_45 : _GEN_1612; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1614 = 8'h4e == _GEN_106 ? _double_bytes_0_T_46 : _GEN_1613; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1615 = 8'h4f == _GEN_106 ? _double_bytes_0_T_47 : _GEN_1614; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] double_bytes_5_0 = _GEN_82 ? _GEN_1615 : 16'h0; // @[matcher_pisa.scala 145:46 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_1617 = 8'h20 == _GEN_107 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53 matcher_pisa.scala 144:41]
  wire [15:0] _GEN_1618 = 8'h21 == _GEN_107 ? _double_bytes_0_T_1 : _GEN_1617; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1619 = 8'h22 == _GEN_107 ? _double_bytes_0_T_2 : _GEN_1618; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1620 = 8'h23 == _GEN_107 ? _double_bytes_0_T_3 : _GEN_1619; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1621 = 8'h24 == _GEN_107 ? _double_bytes_0_T_4 : _GEN_1620; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1622 = 8'h25 == _GEN_107 ? _double_bytes_0_T_5 : _GEN_1621; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1623 = 8'h26 == _GEN_107 ? _double_bytes_0_T_6 : _GEN_1622; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1624 = 8'h27 == _GEN_107 ? _double_bytes_0_T_7 : _GEN_1623; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1625 = 8'h28 == _GEN_107 ? _double_bytes_0_T_8 : _GEN_1624; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1626 = 8'h29 == _GEN_107 ? _double_bytes_0_T_9 : _GEN_1625; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1627 = 8'h2a == _GEN_107 ? _double_bytes_0_T_10 : _GEN_1626; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1628 = 8'h2b == _GEN_107 ? _double_bytes_0_T_11 : _GEN_1627; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1629 = 8'h2c == _GEN_107 ? _double_bytes_0_T_12 : _GEN_1628; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1630 = 8'h2d == _GEN_107 ? _double_bytes_0_T_13 : _GEN_1629; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1631 = 8'h2e == _GEN_107 ? _double_bytes_0_T_14 : _GEN_1630; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1632 = 8'h2f == _GEN_107 ? _double_bytes_0_T_15 : _GEN_1631; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1633 = 8'h30 == _GEN_107 ? _double_bytes_0_T_16 : _GEN_1632; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1634 = 8'h31 == _GEN_107 ? _double_bytes_0_T_17 : _GEN_1633; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1635 = 8'h32 == _GEN_107 ? _double_bytes_0_T_18 : _GEN_1634; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1636 = 8'h33 == _GEN_107 ? _double_bytes_0_T_19 : _GEN_1635; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1637 = 8'h34 == _GEN_107 ? _double_bytes_0_T_20 : _GEN_1636; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1638 = 8'h35 == _GEN_107 ? _double_bytes_0_T_21 : _GEN_1637; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1639 = 8'h36 == _GEN_107 ? _double_bytes_0_T_22 : _GEN_1638; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1640 = 8'h37 == _GEN_107 ? _double_bytes_0_T_23 : _GEN_1639; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1641 = 8'h38 == _GEN_107 ? _double_bytes_0_T_24 : _GEN_1640; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1642 = 8'h39 == _GEN_107 ? _double_bytes_0_T_25 : _GEN_1641; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1643 = 8'h3a == _GEN_107 ? _double_bytes_0_T_26 : _GEN_1642; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1644 = 8'h3b == _GEN_107 ? _double_bytes_0_T_27 : _GEN_1643; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1645 = 8'h3c == _GEN_107 ? _double_bytes_0_T_28 : _GEN_1644; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1646 = 8'h3d == _GEN_107 ? _double_bytes_0_T_29 : _GEN_1645; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1647 = 8'h3e == _GEN_107 ? _double_bytes_0_T_30 : _GEN_1646; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1648 = 8'h3f == _GEN_107 ? _double_bytes_0_T_31 : _GEN_1647; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1649 = 8'h40 == _GEN_107 ? _double_bytes_0_T_32 : _GEN_1648; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1650 = 8'h41 == _GEN_107 ? _double_bytes_0_T_33 : _GEN_1649; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1651 = 8'h42 == _GEN_107 ? _double_bytes_0_T_34 : _GEN_1650; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1652 = 8'h43 == _GEN_107 ? _double_bytes_0_T_35 : _GEN_1651; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1653 = 8'h44 == _GEN_107 ? _double_bytes_0_T_36 : _GEN_1652; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1654 = 8'h45 == _GEN_107 ? _double_bytes_0_T_37 : _GEN_1653; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1655 = 8'h46 == _GEN_107 ? _double_bytes_0_T_38 : _GEN_1654; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1656 = 8'h47 == _GEN_107 ? _double_bytes_0_T_39 : _GEN_1655; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1657 = 8'h48 == _GEN_107 ? _double_bytes_0_T_40 : _GEN_1656; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1658 = 8'h49 == _GEN_107 ? _double_bytes_0_T_41 : _GEN_1657; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1659 = 8'h4a == _GEN_107 ? _double_bytes_0_T_42 : _GEN_1658; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1660 = 8'h4b == _GEN_107 ? _double_bytes_0_T_43 : _GEN_1659; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1661 = 8'h4c == _GEN_107 ? _double_bytes_0_T_44 : _GEN_1660; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1662 = 8'h4d == _GEN_107 ? _double_bytes_0_T_45 : _GEN_1661; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1663 = 8'h4e == _GEN_107 ? _double_bytes_0_T_46 : _GEN_1662; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] _GEN_1664 = 8'h4f == _GEN_107 ? _double_bytes_0_T_47 : _GEN_1663; // @[matcher_pisa.scala 147:85 matcher_pisa.scala 148:53]
  wire [15:0] double_bytes_5_1 = _GEN_83 ? _GEN_1664 : 16'h0; // @[matcher_pisa.scala 145:46 matcher_pisa.scala 144:41]
  wire [31:0] _groups_5_T_1 = {double_bytes_5_0,double_bytes_5_1}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_1666 = _GEN_61 == 2'h2 ? _groups_5_T_1 : _GEN_1567; // @[matcher_pisa.scala 139:50 matcher_pisa.scala 153:31]
  wire [31:0] _GEN_1667 = 8'h50 == _GEN_106 ? _groups_0_T_2 : 32'h0; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39 matcher_pisa.scala 158:31]
  wire [31:0] _GEN_1668 = 8'h51 == _GEN_106 ? _groups_0_T_3 : _GEN_1667; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1669 = 8'h52 == _GEN_106 ? _groups_0_T_4 : _GEN_1668; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1670 = 8'h53 == _GEN_106 ? _groups_0_T_5 : _GEN_1669; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1671 = 8'h54 == _GEN_106 ? _groups_0_T_6 : _GEN_1670; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1672 = 8'h55 == _GEN_106 ? _groups_0_T_7 : _GEN_1671; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1673 = 8'h56 == _GEN_106 ? _groups_0_T_8 : _GEN_1672; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1674 = 8'h57 == _GEN_106 ? _groups_0_T_9 : _GEN_1673; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1675 = 8'h58 == _GEN_106 ? _groups_0_T_10 : _GEN_1674; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1676 = 8'h59 == _GEN_106 ? _groups_0_T_11 : _GEN_1675; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1677 = 8'h5a == _GEN_106 ? _groups_0_T_12 : _GEN_1676; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1678 = 8'h5b == _GEN_106 ? _groups_0_T_13 : _GEN_1677; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1679 = 8'h5c == _GEN_106 ? _groups_0_T_14 : _GEN_1678; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1680 = 8'h5d == _GEN_106 ? _groups_0_T_15 : _GEN_1679; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1681 = 8'h5e == _GEN_106 ? _groups_0_T_16 : _GEN_1680; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1682 = 8'h5f == _GEN_106 ? _groups_0_T_17 : _GEN_1681; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1683 = 8'h60 == _GEN_106 ? _groups_0_T_18 : _GEN_1682; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1684 = 8'h61 == _GEN_106 ? _groups_0_T_19 : _GEN_1683; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1685 = 8'h62 == _GEN_106 ? _groups_0_T_20 : _GEN_1684; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1686 = 8'h63 == _GEN_106 ? _groups_0_T_21 : _GEN_1685; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1687 = 8'h64 == _GEN_106 ? _groups_0_T_22 : _GEN_1686; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1688 = 8'h65 == _GEN_106 ? _groups_0_T_23 : _GEN_1687; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1689 = 8'h66 == _GEN_106 ? _groups_0_T_24 : _GEN_1688; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1690 = 8'h67 == _GEN_106 ? _groups_0_T_25 : _GEN_1689; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1691 = 8'h68 == _GEN_106 ? _groups_0_T_26 : _GEN_1690; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1692 = 8'h69 == _GEN_106 ? _groups_0_T_27 : _GEN_1691; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1693 = 8'h6a == _GEN_106 ? _groups_0_T_28 : _GEN_1692; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1694 = 8'h6b == _GEN_106 ? _groups_0_T_29 : _GEN_1693; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1695 = 8'h6c == _GEN_106 ? _groups_0_T_30 : _GEN_1694; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1696 = 8'h6d == _GEN_106 ? _groups_0_T_31 : _GEN_1695; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1697 = 8'h6e == _GEN_106 ? _groups_0_T_32 : _GEN_1696; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] _GEN_1698 = 8'h6f == _GEN_106 ? _groups_0_T_33 : _GEN_1697; // @[matcher_pisa.scala 160:77 matcher_pisa.scala 161:39]
  wire [31:0] groups_5 = _GEN_61 == 2'h3 ? _GEN_1698 : _GEN_1666; // @[matcher_pisa.scala 155:50]
  wire [191:0] _io_match_key_T = {groups_0,groups_1,groups_2,groups_3,groups_4,groups_5}; // @[Cat.scala 30:58]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_96 = phv_data_96; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_97 = phv_data_97; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_98 = phv_data_98; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_99 = phv_data_99; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_100 = phv_data_100; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_101 = phv_data_101; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_102 = phv_data_102; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_103 = phv_data_103; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_104 = phv_data_104; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_105 = phv_data_105; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_106 = phv_data_106; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_107 = phv_data_107; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_108 = phv_data_108; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_109 = phv_data_109; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_110 = phv_data_110; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_111 = phv_data_111; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_112 = phv_data_112; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_113 = phv_data_113; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_114 = phv_data_114; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_115 = phv_data_115; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_116 = phv_data_116; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_117 = phv_data_117; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_118 = phv_data_118; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_119 = phv_data_119; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_120 = phv_data_120; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_121 = phv_data_121; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_122 = phv_data_122; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_123 = phv_data_123; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_124 = phv_data_124; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_125 = phv_data_125; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_126 = phv_data_126; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_127 = phv_data_127; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_128 = phv_data_128; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_129 = phv_data_129; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_130 = phv_data_130; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_131 = phv_data_131; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_132 = phv_data_132; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_133 = phv_data_133; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_134 = phv_data_134; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_135 = phv_data_135; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_136 = phv_data_136; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_137 = phv_data_137; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_138 = phv_data_138; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_139 = phv_data_139; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_140 = phv_data_140; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_141 = phv_data_141; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_142 = phv_data_142; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_143 = phv_data_143; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_144 = phv_data_144; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_145 = phv_data_145; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_146 = phv_data_146; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_147 = phv_data_147; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_148 = phv_data_148; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_149 = phv_data_149; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_150 = phv_data_150; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_151 = phv_data_151; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_152 = phv_data_152; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_153 = phv_data_153; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_154 = phv_data_154; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_155 = phv_data_155; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_156 = phv_data_156; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_157 = phv_data_157; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_158 = phv_data_158; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_159 = phv_data_159; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_160 = phv_data_160; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_161 = phv_data_161; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_162 = phv_data_162; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_163 = phv_data_163; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_164 = phv_data_164; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_165 = phv_data_165; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_166 = phv_data_166; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_167 = phv_data_167; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_168 = phv_data_168; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_169 = phv_data_169; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_170 = phv_data_170; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_171 = phv_data_171; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_172 = phv_data_172; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_173 = phv_data_173; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_174 = phv_data_174; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_175 = phv_data_175; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_176 = phv_data_176; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_177 = phv_data_177; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_178 = phv_data_178; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_179 = phv_data_179; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_180 = phv_data_180; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_181 = phv_data_181; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_182 = phv_data_182; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_183 = phv_data_183; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_184 = phv_data_184; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_185 = phv_data_185; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_186 = phv_data_186; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_187 = phv_data_187; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_188 = phv_data_188; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_189 = phv_data_189; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_190 = phv_data_190; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_191 = phv_data_191; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_192 = phv_data_192; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_193 = phv_data_193; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_194 = phv_data_194; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_195 = phv_data_195; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_196 = phv_data_196; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_197 = phv_data_197; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_198 = phv_data_198; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_199 = phv_data_199; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_200 = phv_data_200; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_201 = phv_data_201; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_202 = phv_data_202; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_203 = phv_data_203; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_204 = phv_data_204; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_205 = phv_data_205; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_206 = phv_data_206; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_207 = phv_data_207; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_208 = phv_data_208; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_209 = phv_data_209; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_210 = phv_data_210; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_211 = phv_data_211; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_212 = phv_data_212; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_213 = phv_data_213; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_214 = phv_data_214; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_215 = phv_data_215; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_216 = phv_data_216; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_217 = phv_data_217; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_218 = phv_data_218; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_219 = phv_data_219; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_220 = phv_data_220; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_221 = phv_data_221; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_222 = phv_data_222; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_223 = phv_data_223; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_224 = phv_data_224; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_225 = phv_data_225; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_226 = phv_data_226; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_227 = phv_data_227; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_228 = phv_data_228; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_229 = phv_data_229; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_230 = phv_data_230; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_231 = phv_data_231; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_232 = phv_data_232; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_233 = phv_data_233; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_234 = phv_data_234; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_235 = phv_data_235; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_236 = phv_data_236; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_237 = phv_data_237; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_238 = phv_data_238; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_239 = phv_data_239; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_240 = phv_data_240; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_241 = phv_data_241; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_242 = phv_data_242; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_243 = phv_data_243; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_244 = phv_data_244; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_245 = phv_data_245; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_246 = phv_data_246; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_247 = phv_data_247; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_248 = phv_data_248; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_249 = phv_data_249; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_250 = phv_data_250; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_251 = phv_data_251; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_252 = phv_data_252; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_253 = phv_data_253; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_254 = phv_data_254; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_data_255 = phv_data_255; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[matcher_pisa.scala 112:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[matcher_pisa.scala 112:25]
  assign io_match_key = phv_is_valid_processor ? _io_match_key_T : 192'h0; // @[matcher_pisa.scala 116:39 matcher_pisa.scala 166:26 matcher_pisa.scala 168:26]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[matcher_pisa.scala 111:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[matcher_pisa.scala 111:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[matcher_pisa.scala 111:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[matcher_pisa.scala 111:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[matcher_pisa.scala 111:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[matcher_pisa.scala 111:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[matcher_pisa.scala 111:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[matcher_pisa.scala 111:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[matcher_pisa.scala 111:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[matcher_pisa.scala 111:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[matcher_pisa.scala 111:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[matcher_pisa.scala 111:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[matcher_pisa.scala 111:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[matcher_pisa.scala 111:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[matcher_pisa.scala 111:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[matcher_pisa.scala 111:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[matcher_pisa.scala 111:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[matcher_pisa.scala 111:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[matcher_pisa.scala 111:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[matcher_pisa.scala 111:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[matcher_pisa.scala 111:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[matcher_pisa.scala 111:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[matcher_pisa.scala 111:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[matcher_pisa.scala 111:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[matcher_pisa.scala 111:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[matcher_pisa.scala 111:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[matcher_pisa.scala 111:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[matcher_pisa.scala 111:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[matcher_pisa.scala 111:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[matcher_pisa.scala 111:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[matcher_pisa.scala 111:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[matcher_pisa.scala 111:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[matcher_pisa.scala 111:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[matcher_pisa.scala 111:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[matcher_pisa.scala 111:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[matcher_pisa.scala 111:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[matcher_pisa.scala 111:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[matcher_pisa.scala 111:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[matcher_pisa.scala 111:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[matcher_pisa.scala 111:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[matcher_pisa.scala 111:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[matcher_pisa.scala 111:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[matcher_pisa.scala 111:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[matcher_pisa.scala 111:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[matcher_pisa.scala 111:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[matcher_pisa.scala 111:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[matcher_pisa.scala 111:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[matcher_pisa.scala 111:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[matcher_pisa.scala 111:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[matcher_pisa.scala 111:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[matcher_pisa.scala 111:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[matcher_pisa.scala 111:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[matcher_pisa.scala 111:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[matcher_pisa.scala 111:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[matcher_pisa.scala 111:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[matcher_pisa.scala 111:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[matcher_pisa.scala 111:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[matcher_pisa.scala 111:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[matcher_pisa.scala 111:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[matcher_pisa.scala 111:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[matcher_pisa.scala 111:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[matcher_pisa.scala 111:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[matcher_pisa.scala 111:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[matcher_pisa.scala 111:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[matcher_pisa.scala 111:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[matcher_pisa.scala 111:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[matcher_pisa.scala 111:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[matcher_pisa.scala 111:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[matcher_pisa.scala 111:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[matcher_pisa.scala 111:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[matcher_pisa.scala 111:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[matcher_pisa.scala 111:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[matcher_pisa.scala 111:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[matcher_pisa.scala 111:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[matcher_pisa.scala 111:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[matcher_pisa.scala 111:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[matcher_pisa.scala 111:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[matcher_pisa.scala 111:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[matcher_pisa.scala 111:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[matcher_pisa.scala 111:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[matcher_pisa.scala 111:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[matcher_pisa.scala 111:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[matcher_pisa.scala 111:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[matcher_pisa.scala 111:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[matcher_pisa.scala 111:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[matcher_pisa.scala 111:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[matcher_pisa.scala 111:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[matcher_pisa.scala 111:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[matcher_pisa.scala 111:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[matcher_pisa.scala 111:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[matcher_pisa.scala 111:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[matcher_pisa.scala 111:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[matcher_pisa.scala 111:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[matcher_pisa.scala 111:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[matcher_pisa.scala 111:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[matcher_pisa.scala 111:13]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[matcher_pisa.scala 111:13]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[matcher_pisa.scala 111:13]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[matcher_pisa.scala 111:13]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[matcher_pisa.scala 111:13]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[matcher_pisa.scala 111:13]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[matcher_pisa.scala 111:13]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[matcher_pisa.scala 111:13]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[matcher_pisa.scala 111:13]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[matcher_pisa.scala 111:13]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[matcher_pisa.scala 111:13]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[matcher_pisa.scala 111:13]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[matcher_pisa.scala 111:13]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[matcher_pisa.scala 111:13]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[matcher_pisa.scala 111:13]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[matcher_pisa.scala 111:13]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[matcher_pisa.scala 111:13]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[matcher_pisa.scala 111:13]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[matcher_pisa.scala 111:13]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[matcher_pisa.scala 111:13]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[matcher_pisa.scala 111:13]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[matcher_pisa.scala 111:13]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[matcher_pisa.scala 111:13]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[matcher_pisa.scala 111:13]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[matcher_pisa.scala 111:13]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[matcher_pisa.scala 111:13]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[matcher_pisa.scala 111:13]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[matcher_pisa.scala 111:13]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[matcher_pisa.scala 111:13]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[matcher_pisa.scala 111:13]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[matcher_pisa.scala 111:13]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[matcher_pisa.scala 111:13]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[matcher_pisa.scala 111:13]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[matcher_pisa.scala 111:13]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[matcher_pisa.scala 111:13]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[matcher_pisa.scala 111:13]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[matcher_pisa.scala 111:13]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[matcher_pisa.scala 111:13]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[matcher_pisa.scala 111:13]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[matcher_pisa.scala 111:13]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[matcher_pisa.scala 111:13]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[matcher_pisa.scala 111:13]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[matcher_pisa.scala 111:13]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[matcher_pisa.scala 111:13]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[matcher_pisa.scala 111:13]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[matcher_pisa.scala 111:13]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[matcher_pisa.scala 111:13]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[matcher_pisa.scala 111:13]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[matcher_pisa.scala 111:13]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[matcher_pisa.scala 111:13]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[matcher_pisa.scala 111:13]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[matcher_pisa.scala 111:13]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[matcher_pisa.scala 111:13]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[matcher_pisa.scala 111:13]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[matcher_pisa.scala 111:13]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[matcher_pisa.scala 111:13]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[matcher_pisa.scala 111:13]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[matcher_pisa.scala 111:13]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[matcher_pisa.scala 111:13]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[matcher_pisa.scala 111:13]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[matcher_pisa.scala 111:13]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[matcher_pisa.scala 111:13]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[matcher_pisa.scala 111:13]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[matcher_pisa.scala 111:13]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[matcher_pisa.scala 111:13]
    phv_data_160 <= io_pipe_phv_in_data_160; // @[matcher_pisa.scala 111:13]
    phv_data_161 <= io_pipe_phv_in_data_161; // @[matcher_pisa.scala 111:13]
    phv_data_162 <= io_pipe_phv_in_data_162; // @[matcher_pisa.scala 111:13]
    phv_data_163 <= io_pipe_phv_in_data_163; // @[matcher_pisa.scala 111:13]
    phv_data_164 <= io_pipe_phv_in_data_164; // @[matcher_pisa.scala 111:13]
    phv_data_165 <= io_pipe_phv_in_data_165; // @[matcher_pisa.scala 111:13]
    phv_data_166 <= io_pipe_phv_in_data_166; // @[matcher_pisa.scala 111:13]
    phv_data_167 <= io_pipe_phv_in_data_167; // @[matcher_pisa.scala 111:13]
    phv_data_168 <= io_pipe_phv_in_data_168; // @[matcher_pisa.scala 111:13]
    phv_data_169 <= io_pipe_phv_in_data_169; // @[matcher_pisa.scala 111:13]
    phv_data_170 <= io_pipe_phv_in_data_170; // @[matcher_pisa.scala 111:13]
    phv_data_171 <= io_pipe_phv_in_data_171; // @[matcher_pisa.scala 111:13]
    phv_data_172 <= io_pipe_phv_in_data_172; // @[matcher_pisa.scala 111:13]
    phv_data_173 <= io_pipe_phv_in_data_173; // @[matcher_pisa.scala 111:13]
    phv_data_174 <= io_pipe_phv_in_data_174; // @[matcher_pisa.scala 111:13]
    phv_data_175 <= io_pipe_phv_in_data_175; // @[matcher_pisa.scala 111:13]
    phv_data_176 <= io_pipe_phv_in_data_176; // @[matcher_pisa.scala 111:13]
    phv_data_177 <= io_pipe_phv_in_data_177; // @[matcher_pisa.scala 111:13]
    phv_data_178 <= io_pipe_phv_in_data_178; // @[matcher_pisa.scala 111:13]
    phv_data_179 <= io_pipe_phv_in_data_179; // @[matcher_pisa.scala 111:13]
    phv_data_180 <= io_pipe_phv_in_data_180; // @[matcher_pisa.scala 111:13]
    phv_data_181 <= io_pipe_phv_in_data_181; // @[matcher_pisa.scala 111:13]
    phv_data_182 <= io_pipe_phv_in_data_182; // @[matcher_pisa.scala 111:13]
    phv_data_183 <= io_pipe_phv_in_data_183; // @[matcher_pisa.scala 111:13]
    phv_data_184 <= io_pipe_phv_in_data_184; // @[matcher_pisa.scala 111:13]
    phv_data_185 <= io_pipe_phv_in_data_185; // @[matcher_pisa.scala 111:13]
    phv_data_186 <= io_pipe_phv_in_data_186; // @[matcher_pisa.scala 111:13]
    phv_data_187 <= io_pipe_phv_in_data_187; // @[matcher_pisa.scala 111:13]
    phv_data_188 <= io_pipe_phv_in_data_188; // @[matcher_pisa.scala 111:13]
    phv_data_189 <= io_pipe_phv_in_data_189; // @[matcher_pisa.scala 111:13]
    phv_data_190 <= io_pipe_phv_in_data_190; // @[matcher_pisa.scala 111:13]
    phv_data_191 <= io_pipe_phv_in_data_191; // @[matcher_pisa.scala 111:13]
    phv_data_192 <= io_pipe_phv_in_data_192; // @[matcher_pisa.scala 111:13]
    phv_data_193 <= io_pipe_phv_in_data_193; // @[matcher_pisa.scala 111:13]
    phv_data_194 <= io_pipe_phv_in_data_194; // @[matcher_pisa.scala 111:13]
    phv_data_195 <= io_pipe_phv_in_data_195; // @[matcher_pisa.scala 111:13]
    phv_data_196 <= io_pipe_phv_in_data_196; // @[matcher_pisa.scala 111:13]
    phv_data_197 <= io_pipe_phv_in_data_197; // @[matcher_pisa.scala 111:13]
    phv_data_198 <= io_pipe_phv_in_data_198; // @[matcher_pisa.scala 111:13]
    phv_data_199 <= io_pipe_phv_in_data_199; // @[matcher_pisa.scala 111:13]
    phv_data_200 <= io_pipe_phv_in_data_200; // @[matcher_pisa.scala 111:13]
    phv_data_201 <= io_pipe_phv_in_data_201; // @[matcher_pisa.scala 111:13]
    phv_data_202 <= io_pipe_phv_in_data_202; // @[matcher_pisa.scala 111:13]
    phv_data_203 <= io_pipe_phv_in_data_203; // @[matcher_pisa.scala 111:13]
    phv_data_204 <= io_pipe_phv_in_data_204; // @[matcher_pisa.scala 111:13]
    phv_data_205 <= io_pipe_phv_in_data_205; // @[matcher_pisa.scala 111:13]
    phv_data_206 <= io_pipe_phv_in_data_206; // @[matcher_pisa.scala 111:13]
    phv_data_207 <= io_pipe_phv_in_data_207; // @[matcher_pisa.scala 111:13]
    phv_data_208 <= io_pipe_phv_in_data_208; // @[matcher_pisa.scala 111:13]
    phv_data_209 <= io_pipe_phv_in_data_209; // @[matcher_pisa.scala 111:13]
    phv_data_210 <= io_pipe_phv_in_data_210; // @[matcher_pisa.scala 111:13]
    phv_data_211 <= io_pipe_phv_in_data_211; // @[matcher_pisa.scala 111:13]
    phv_data_212 <= io_pipe_phv_in_data_212; // @[matcher_pisa.scala 111:13]
    phv_data_213 <= io_pipe_phv_in_data_213; // @[matcher_pisa.scala 111:13]
    phv_data_214 <= io_pipe_phv_in_data_214; // @[matcher_pisa.scala 111:13]
    phv_data_215 <= io_pipe_phv_in_data_215; // @[matcher_pisa.scala 111:13]
    phv_data_216 <= io_pipe_phv_in_data_216; // @[matcher_pisa.scala 111:13]
    phv_data_217 <= io_pipe_phv_in_data_217; // @[matcher_pisa.scala 111:13]
    phv_data_218 <= io_pipe_phv_in_data_218; // @[matcher_pisa.scala 111:13]
    phv_data_219 <= io_pipe_phv_in_data_219; // @[matcher_pisa.scala 111:13]
    phv_data_220 <= io_pipe_phv_in_data_220; // @[matcher_pisa.scala 111:13]
    phv_data_221 <= io_pipe_phv_in_data_221; // @[matcher_pisa.scala 111:13]
    phv_data_222 <= io_pipe_phv_in_data_222; // @[matcher_pisa.scala 111:13]
    phv_data_223 <= io_pipe_phv_in_data_223; // @[matcher_pisa.scala 111:13]
    phv_data_224 <= io_pipe_phv_in_data_224; // @[matcher_pisa.scala 111:13]
    phv_data_225 <= io_pipe_phv_in_data_225; // @[matcher_pisa.scala 111:13]
    phv_data_226 <= io_pipe_phv_in_data_226; // @[matcher_pisa.scala 111:13]
    phv_data_227 <= io_pipe_phv_in_data_227; // @[matcher_pisa.scala 111:13]
    phv_data_228 <= io_pipe_phv_in_data_228; // @[matcher_pisa.scala 111:13]
    phv_data_229 <= io_pipe_phv_in_data_229; // @[matcher_pisa.scala 111:13]
    phv_data_230 <= io_pipe_phv_in_data_230; // @[matcher_pisa.scala 111:13]
    phv_data_231 <= io_pipe_phv_in_data_231; // @[matcher_pisa.scala 111:13]
    phv_data_232 <= io_pipe_phv_in_data_232; // @[matcher_pisa.scala 111:13]
    phv_data_233 <= io_pipe_phv_in_data_233; // @[matcher_pisa.scala 111:13]
    phv_data_234 <= io_pipe_phv_in_data_234; // @[matcher_pisa.scala 111:13]
    phv_data_235 <= io_pipe_phv_in_data_235; // @[matcher_pisa.scala 111:13]
    phv_data_236 <= io_pipe_phv_in_data_236; // @[matcher_pisa.scala 111:13]
    phv_data_237 <= io_pipe_phv_in_data_237; // @[matcher_pisa.scala 111:13]
    phv_data_238 <= io_pipe_phv_in_data_238; // @[matcher_pisa.scala 111:13]
    phv_data_239 <= io_pipe_phv_in_data_239; // @[matcher_pisa.scala 111:13]
    phv_data_240 <= io_pipe_phv_in_data_240; // @[matcher_pisa.scala 111:13]
    phv_data_241 <= io_pipe_phv_in_data_241; // @[matcher_pisa.scala 111:13]
    phv_data_242 <= io_pipe_phv_in_data_242; // @[matcher_pisa.scala 111:13]
    phv_data_243 <= io_pipe_phv_in_data_243; // @[matcher_pisa.scala 111:13]
    phv_data_244 <= io_pipe_phv_in_data_244; // @[matcher_pisa.scala 111:13]
    phv_data_245 <= io_pipe_phv_in_data_245; // @[matcher_pisa.scala 111:13]
    phv_data_246 <= io_pipe_phv_in_data_246; // @[matcher_pisa.scala 111:13]
    phv_data_247 <= io_pipe_phv_in_data_247; // @[matcher_pisa.scala 111:13]
    phv_data_248 <= io_pipe_phv_in_data_248; // @[matcher_pisa.scala 111:13]
    phv_data_249 <= io_pipe_phv_in_data_249; // @[matcher_pisa.scala 111:13]
    phv_data_250 <= io_pipe_phv_in_data_250; // @[matcher_pisa.scala 111:13]
    phv_data_251 <= io_pipe_phv_in_data_251; // @[matcher_pisa.scala 111:13]
    phv_data_252 <= io_pipe_phv_in_data_252; // @[matcher_pisa.scala 111:13]
    phv_data_253 <= io_pipe_phv_in_data_253; // @[matcher_pisa.scala 111:13]
    phv_data_254 <= io_pipe_phv_in_data_254; // @[matcher_pisa.scala 111:13]
    phv_data_255 <= io_pipe_phv_in_data_255; // @[matcher_pisa.scala 111:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[matcher_pisa.scala 111:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[matcher_pisa.scala 111:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[matcher_pisa.scala 111:13]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_data_160 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  phv_data_161 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  phv_data_162 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  phv_data_163 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  phv_data_164 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  phv_data_165 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  phv_data_166 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  phv_data_167 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  phv_data_168 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  phv_data_169 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  phv_data_170 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  phv_data_171 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  phv_data_172 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  phv_data_173 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  phv_data_174 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  phv_data_175 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  phv_data_176 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_data_177 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_data_178 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  phv_data_179 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  phv_data_180 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  phv_data_181 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  phv_data_182 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  phv_data_183 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  phv_data_184 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  phv_data_185 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  phv_data_186 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  phv_data_187 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  phv_data_188 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  phv_data_189 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  phv_data_190 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  phv_data_191 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  phv_data_192 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  phv_data_193 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  phv_data_194 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  phv_data_195 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  phv_data_196 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  phv_data_197 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  phv_data_198 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  phv_data_199 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  phv_data_200 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  phv_data_201 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  phv_data_202 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  phv_data_203 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  phv_data_204 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  phv_data_205 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  phv_data_206 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  phv_data_207 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  phv_data_208 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  phv_data_209 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  phv_data_210 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  phv_data_211 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  phv_data_212 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  phv_data_213 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  phv_data_214 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  phv_data_215 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  phv_data_216 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  phv_data_217 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  phv_data_218 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  phv_data_219 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  phv_data_220 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  phv_data_221 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  phv_data_222 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  phv_data_223 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  phv_data_224 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  phv_data_225 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  phv_data_226 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  phv_data_227 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  phv_data_228 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  phv_data_229 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  phv_data_230 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  phv_data_231 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  phv_data_232 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  phv_data_233 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  phv_data_234 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  phv_data_235 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  phv_data_236 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  phv_data_237 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  phv_data_238 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  phv_data_239 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  phv_data_240 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  phv_data_241 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  phv_data_242 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  phv_data_243 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  phv_data_244 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  phv_data_245 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  phv_data_246 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  phv_data_247 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  phv_data_248 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  phv_data_249 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  phv_data_250 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  phv_data_251 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  phv_data_252 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  phv_data_253 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  phv_data_254 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  phv_data_255 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_256[3:0];
  _RAND_257 = {1{`RANDOM}};
  phv_next_config_id = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_258[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
