module PrimitiveGetSource(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [3:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  input         io_pipe_phv_in_valid,
  input         io_pipe_phv_in_last,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [3:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  output        io_pipe_phv_out_valid,
  output        io_pipe_phv_out_last,
  input  [31:0] io_vliw_in_0,
  input  [31:0] io_vliw_in_1,
  input  [31:0] io_vliw_in_2,
  input  [31:0] io_vliw_in_3,
  input  [7:0]  io_offset_in_0,
  input  [7:0]  io_offset_in_1,
  input  [7:0]  io_offset_in_2,
  input  [7:0]  io_offset_in_3,
  input  [7:0]  io_length_in_0,
  input  [7:0]  io_length_in_1,
  input  [7:0]  io_length_in_2,
  input  [7:0]  io_length_in_3,
  output [31:0] io_vliw_out_0,
  output [31:0] io_vliw_out_1,
  output [31:0] io_vliw_out_2,
  output [31:0] io_vliw_out_3,
  output [31:0] io_field_out_0,
  output [31:0] io_field_out_1,
  output [31:0] io_field_out_2,
  output [31:0] io_field_out_3,
  output [3:0]  io_mask_out_0,
  output [3:0]  io_mask_out_1,
  output [3:0]  io_mask_out_2,
  output [3:0]  io_mask_out_3,
  output [1:0]  io_bias_out_0,
  output [1:0]  io_bias_out_1,
  output [1:0]  io_bias_out_2,
  output [1:0]  io_bias_out_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[executor.scala 151:22]
  reg [7:0] phv_data_1; // @[executor.scala 151:22]
  reg [7:0] phv_data_2; // @[executor.scala 151:22]
  reg [7:0] phv_data_3; // @[executor.scala 151:22]
  reg [7:0] phv_data_4; // @[executor.scala 151:22]
  reg [7:0] phv_data_5; // @[executor.scala 151:22]
  reg [7:0] phv_data_6; // @[executor.scala 151:22]
  reg [7:0] phv_data_7; // @[executor.scala 151:22]
  reg [7:0] phv_data_8; // @[executor.scala 151:22]
  reg [7:0] phv_data_9; // @[executor.scala 151:22]
  reg [7:0] phv_data_10; // @[executor.scala 151:22]
  reg [7:0] phv_data_11; // @[executor.scala 151:22]
  reg [7:0] phv_data_12; // @[executor.scala 151:22]
  reg [7:0] phv_data_13; // @[executor.scala 151:22]
  reg [7:0] phv_data_14; // @[executor.scala 151:22]
  reg [7:0] phv_data_15; // @[executor.scala 151:22]
  reg [7:0] phv_data_16; // @[executor.scala 151:22]
  reg [7:0] phv_data_17; // @[executor.scala 151:22]
  reg [7:0] phv_data_18; // @[executor.scala 151:22]
  reg [7:0] phv_data_19; // @[executor.scala 151:22]
  reg [7:0] phv_data_20; // @[executor.scala 151:22]
  reg [7:0] phv_data_21; // @[executor.scala 151:22]
  reg [7:0] phv_data_22; // @[executor.scala 151:22]
  reg [7:0] phv_data_23; // @[executor.scala 151:22]
  reg [7:0] phv_data_24; // @[executor.scala 151:22]
  reg [7:0] phv_data_25; // @[executor.scala 151:22]
  reg [7:0] phv_data_26; // @[executor.scala 151:22]
  reg [7:0] phv_data_27; // @[executor.scala 151:22]
  reg [7:0] phv_data_28; // @[executor.scala 151:22]
  reg [7:0] phv_data_29; // @[executor.scala 151:22]
  reg [7:0] phv_data_30; // @[executor.scala 151:22]
  reg [7:0] phv_data_31; // @[executor.scala 151:22]
  reg [7:0] phv_data_32; // @[executor.scala 151:22]
  reg [7:0] phv_data_33; // @[executor.scala 151:22]
  reg [7:0] phv_data_34; // @[executor.scala 151:22]
  reg [7:0] phv_data_35; // @[executor.scala 151:22]
  reg [7:0] phv_data_36; // @[executor.scala 151:22]
  reg [7:0] phv_data_37; // @[executor.scala 151:22]
  reg [7:0] phv_data_38; // @[executor.scala 151:22]
  reg [7:0] phv_data_39; // @[executor.scala 151:22]
  reg [7:0] phv_data_40; // @[executor.scala 151:22]
  reg [7:0] phv_data_41; // @[executor.scala 151:22]
  reg [7:0] phv_data_42; // @[executor.scala 151:22]
  reg [7:0] phv_data_43; // @[executor.scala 151:22]
  reg [7:0] phv_data_44; // @[executor.scala 151:22]
  reg [7:0] phv_data_45; // @[executor.scala 151:22]
  reg [7:0] phv_data_46; // @[executor.scala 151:22]
  reg [7:0] phv_data_47; // @[executor.scala 151:22]
  reg [7:0] phv_data_48; // @[executor.scala 151:22]
  reg [7:0] phv_data_49; // @[executor.scala 151:22]
  reg [7:0] phv_data_50; // @[executor.scala 151:22]
  reg [7:0] phv_data_51; // @[executor.scala 151:22]
  reg [7:0] phv_data_52; // @[executor.scala 151:22]
  reg [7:0] phv_data_53; // @[executor.scala 151:22]
  reg [7:0] phv_data_54; // @[executor.scala 151:22]
  reg [7:0] phv_data_55; // @[executor.scala 151:22]
  reg [7:0] phv_data_56; // @[executor.scala 151:22]
  reg [7:0] phv_data_57; // @[executor.scala 151:22]
  reg [7:0] phv_data_58; // @[executor.scala 151:22]
  reg [7:0] phv_data_59; // @[executor.scala 151:22]
  reg [7:0] phv_data_60; // @[executor.scala 151:22]
  reg [7:0] phv_data_61; // @[executor.scala 151:22]
  reg [7:0] phv_data_62; // @[executor.scala 151:22]
  reg [7:0] phv_data_63; // @[executor.scala 151:22]
  reg [7:0] phv_data_64; // @[executor.scala 151:22]
  reg [7:0] phv_data_65; // @[executor.scala 151:22]
  reg [7:0] phv_data_66; // @[executor.scala 151:22]
  reg [7:0] phv_data_67; // @[executor.scala 151:22]
  reg [7:0] phv_data_68; // @[executor.scala 151:22]
  reg [7:0] phv_data_69; // @[executor.scala 151:22]
  reg [7:0] phv_data_70; // @[executor.scala 151:22]
  reg [7:0] phv_data_71; // @[executor.scala 151:22]
  reg [7:0] phv_data_72; // @[executor.scala 151:22]
  reg [7:0] phv_data_73; // @[executor.scala 151:22]
  reg [7:0] phv_data_74; // @[executor.scala 151:22]
  reg [7:0] phv_data_75; // @[executor.scala 151:22]
  reg [7:0] phv_data_76; // @[executor.scala 151:22]
  reg [7:0] phv_data_77; // @[executor.scala 151:22]
  reg [7:0] phv_data_78; // @[executor.scala 151:22]
  reg [7:0] phv_data_79; // @[executor.scala 151:22]
  reg [7:0] phv_data_80; // @[executor.scala 151:22]
  reg [7:0] phv_data_81; // @[executor.scala 151:22]
  reg [7:0] phv_data_82; // @[executor.scala 151:22]
  reg [7:0] phv_data_83; // @[executor.scala 151:22]
  reg [7:0] phv_data_84; // @[executor.scala 151:22]
  reg [7:0] phv_data_85; // @[executor.scala 151:22]
  reg [7:0] phv_data_86; // @[executor.scala 151:22]
  reg [7:0] phv_data_87; // @[executor.scala 151:22]
  reg [7:0] phv_data_88; // @[executor.scala 151:22]
  reg [7:0] phv_data_89; // @[executor.scala 151:22]
  reg [7:0] phv_data_90; // @[executor.scala 151:22]
  reg [7:0] phv_data_91; // @[executor.scala 151:22]
  reg [7:0] phv_data_92; // @[executor.scala 151:22]
  reg [7:0] phv_data_93; // @[executor.scala 151:22]
  reg [7:0] phv_data_94; // @[executor.scala 151:22]
  reg [7:0] phv_data_95; // @[executor.scala 151:22]
  reg [7:0] phv_data_96; // @[executor.scala 151:22]
  reg [7:0] phv_data_97; // @[executor.scala 151:22]
  reg [7:0] phv_data_98; // @[executor.scala 151:22]
  reg [7:0] phv_data_99; // @[executor.scala 151:22]
  reg [7:0] phv_data_100; // @[executor.scala 151:22]
  reg [7:0] phv_data_101; // @[executor.scala 151:22]
  reg [7:0] phv_data_102; // @[executor.scala 151:22]
  reg [7:0] phv_data_103; // @[executor.scala 151:22]
  reg [7:0] phv_data_104; // @[executor.scala 151:22]
  reg [7:0] phv_data_105; // @[executor.scala 151:22]
  reg [7:0] phv_data_106; // @[executor.scala 151:22]
  reg [7:0] phv_data_107; // @[executor.scala 151:22]
  reg [7:0] phv_data_108; // @[executor.scala 151:22]
  reg [7:0] phv_data_109; // @[executor.scala 151:22]
  reg [7:0] phv_data_110; // @[executor.scala 151:22]
  reg [7:0] phv_data_111; // @[executor.scala 151:22]
  reg [7:0] phv_data_112; // @[executor.scala 151:22]
  reg [7:0] phv_data_113; // @[executor.scala 151:22]
  reg [7:0] phv_data_114; // @[executor.scala 151:22]
  reg [7:0] phv_data_115; // @[executor.scala 151:22]
  reg [7:0] phv_data_116; // @[executor.scala 151:22]
  reg [7:0] phv_data_117; // @[executor.scala 151:22]
  reg [7:0] phv_data_118; // @[executor.scala 151:22]
  reg [7:0] phv_data_119; // @[executor.scala 151:22]
  reg [7:0] phv_data_120; // @[executor.scala 151:22]
  reg [7:0] phv_data_121; // @[executor.scala 151:22]
  reg [7:0] phv_data_122; // @[executor.scala 151:22]
  reg [7:0] phv_data_123; // @[executor.scala 151:22]
  reg [7:0] phv_data_124; // @[executor.scala 151:22]
  reg [7:0] phv_data_125; // @[executor.scala 151:22]
  reg [7:0] phv_data_126; // @[executor.scala 151:22]
  reg [7:0] phv_data_127; // @[executor.scala 151:22]
  reg [7:0] phv_data_128; // @[executor.scala 151:22]
  reg [7:0] phv_data_129; // @[executor.scala 151:22]
  reg [7:0] phv_data_130; // @[executor.scala 151:22]
  reg [7:0] phv_data_131; // @[executor.scala 151:22]
  reg [7:0] phv_data_132; // @[executor.scala 151:22]
  reg [7:0] phv_data_133; // @[executor.scala 151:22]
  reg [7:0] phv_data_134; // @[executor.scala 151:22]
  reg [7:0] phv_data_135; // @[executor.scala 151:22]
  reg [7:0] phv_data_136; // @[executor.scala 151:22]
  reg [7:0] phv_data_137; // @[executor.scala 151:22]
  reg [7:0] phv_data_138; // @[executor.scala 151:22]
  reg [7:0] phv_data_139; // @[executor.scala 151:22]
  reg [7:0] phv_data_140; // @[executor.scala 151:22]
  reg [7:0] phv_data_141; // @[executor.scala 151:22]
  reg [7:0] phv_data_142; // @[executor.scala 151:22]
  reg [7:0] phv_data_143; // @[executor.scala 151:22]
  reg [7:0] phv_data_144; // @[executor.scala 151:22]
  reg [7:0] phv_data_145; // @[executor.scala 151:22]
  reg [7:0] phv_data_146; // @[executor.scala 151:22]
  reg [7:0] phv_data_147; // @[executor.scala 151:22]
  reg [7:0] phv_data_148; // @[executor.scala 151:22]
  reg [7:0] phv_data_149; // @[executor.scala 151:22]
  reg [7:0] phv_data_150; // @[executor.scala 151:22]
  reg [7:0] phv_data_151; // @[executor.scala 151:22]
  reg [7:0] phv_data_152; // @[executor.scala 151:22]
  reg [7:0] phv_data_153; // @[executor.scala 151:22]
  reg [7:0] phv_data_154; // @[executor.scala 151:22]
  reg [7:0] phv_data_155; // @[executor.scala 151:22]
  reg [7:0] phv_data_156; // @[executor.scala 151:22]
  reg [7:0] phv_data_157; // @[executor.scala 151:22]
  reg [7:0] phv_data_158; // @[executor.scala 151:22]
  reg [7:0] phv_data_159; // @[executor.scala 151:22]
  reg [15:0] phv_header_0; // @[executor.scala 151:22]
  reg [15:0] phv_header_1; // @[executor.scala 151:22]
  reg [15:0] phv_header_2; // @[executor.scala 151:22]
  reg [15:0] phv_header_3; // @[executor.scala 151:22]
  reg [15:0] phv_header_4; // @[executor.scala 151:22]
  reg [15:0] phv_header_5; // @[executor.scala 151:22]
  reg [15:0] phv_header_6; // @[executor.scala 151:22]
  reg [15:0] phv_header_7; // @[executor.scala 151:22]
  reg [15:0] phv_header_8; // @[executor.scala 151:22]
  reg [15:0] phv_header_9; // @[executor.scala 151:22]
  reg [15:0] phv_header_10; // @[executor.scala 151:22]
  reg [15:0] phv_header_11; // @[executor.scala 151:22]
  reg [15:0] phv_header_12; // @[executor.scala 151:22]
  reg [15:0] phv_header_13; // @[executor.scala 151:22]
  reg [15:0] phv_header_14; // @[executor.scala 151:22]
  reg [15:0] phv_header_15; // @[executor.scala 151:22]
  reg [7:0] phv_parse_current_state; // @[executor.scala 151:22]
  reg [7:0] phv_parse_current_offset; // @[executor.scala 151:22]
  reg [15:0] phv_parse_transition_field; // @[executor.scala 151:22]
  reg [3:0] phv_next_processor_id; // @[executor.scala 151:22]
  reg  phv_next_config_id; // @[executor.scala 151:22]
  reg  phv_is_valid_processor; // @[executor.scala 151:22]
  reg  phv_valid; // @[executor.scala 151:22]
  reg  phv_last; // @[executor.scala 151:22]
  reg [31:0] vliw_0; // @[executor.scala 158:23]
  reg [31:0] vliw_1; // @[executor.scala 158:23]
  reg [31:0] vliw_2; // @[executor.scala 158:23]
  reg [31:0] vliw_3; // @[executor.scala 158:23]
  reg [7:0] offset_0; // @[executor.scala 162:25]
  reg [7:0] offset_1; // @[executor.scala 162:25]
  reg [7:0] offset_2; // @[executor.scala 162:25]
  reg [7:0] offset_3; // @[executor.scala 162:25]
  reg [7:0] length_0; // @[executor.scala 163:25]
  reg [7:0] length_1; // @[executor.scala 163:25]
  reg [7:0] length_2; // @[executor.scala 163:25]
  reg [7:0] length_3; // @[executor.scala 163:25]
  wire [3:0] opcode = vliw_0[31:28]; // @[primitive.scala 9:44]
  wire [13:0] io_field_out_0_lo = vliw_0[13:0]; // @[primitive.scala 11:44]
  wire  from_header = length_0 != 8'h0; // @[executor.scala 177:45]
  wire [5:0] total_offset_hi = offset_0[7:2]; // @[executor.scala 191:57]
  wire [7:0] _ending_T_1 = offset_0 + length_0; // @[executor.scala 193:46]
  wire [1:0] ending = _ending_T_1[1:0]; // @[executor.scala 193:58]
  wire [3:0] _GEN_3488 = {{2'd0}, ending}; // @[executor.scala 194:45]
  wire [3:0] _bias_T_1 = 4'h4 - _GEN_3488; // @[executor.scala 194:45]
  wire [1:0] bias = _bias_T_1[1:0]; // @[executor.scala 194:54]
  wire [7:0] total_offset = {total_offset_hi,2'h0}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_1 = 8'h1 == total_offset ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2 = 8'h2 == total_offset ? phv_data_2 : _GEN_1; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3 = 8'h3 == total_offset ? phv_data_3 : _GEN_2; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4 = 8'h4 == total_offset ? phv_data_4 : _GEN_3; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5 = 8'h5 == total_offset ? phv_data_5 : _GEN_4; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6 = 8'h6 == total_offset ? phv_data_6 : _GEN_5; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7 = 8'h7 == total_offset ? phv_data_7 : _GEN_6; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8 = 8'h8 == total_offset ? phv_data_8 : _GEN_7; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_9 = 8'h9 == total_offset ? phv_data_9 : _GEN_8; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_10 = 8'ha == total_offset ? phv_data_10 : _GEN_9; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_11 = 8'hb == total_offset ? phv_data_11 : _GEN_10; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_12 = 8'hc == total_offset ? phv_data_12 : _GEN_11; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_13 = 8'hd == total_offset ? phv_data_13 : _GEN_12; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_14 = 8'he == total_offset ? phv_data_14 : _GEN_13; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_15 = 8'hf == total_offset ? phv_data_15 : _GEN_14; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_16 = 8'h10 == total_offset ? phv_data_16 : _GEN_15; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_17 = 8'h11 == total_offset ? phv_data_17 : _GEN_16; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_18 = 8'h12 == total_offset ? phv_data_18 : _GEN_17; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_19 = 8'h13 == total_offset ? phv_data_19 : _GEN_18; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_20 = 8'h14 == total_offset ? phv_data_20 : _GEN_19; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_21 = 8'h15 == total_offset ? phv_data_21 : _GEN_20; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_22 = 8'h16 == total_offset ? phv_data_22 : _GEN_21; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_23 = 8'h17 == total_offset ? phv_data_23 : _GEN_22; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_24 = 8'h18 == total_offset ? phv_data_24 : _GEN_23; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_25 = 8'h19 == total_offset ? phv_data_25 : _GEN_24; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_26 = 8'h1a == total_offset ? phv_data_26 : _GEN_25; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_27 = 8'h1b == total_offset ? phv_data_27 : _GEN_26; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_28 = 8'h1c == total_offset ? phv_data_28 : _GEN_27; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_29 = 8'h1d == total_offset ? phv_data_29 : _GEN_28; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_30 = 8'h1e == total_offset ? phv_data_30 : _GEN_29; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_31 = 8'h1f == total_offset ? phv_data_31 : _GEN_30; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_32 = 8'h20 == total_offset ? phv_data_32 : _GEN_31; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_33 = 8'h21 == total_offset ? phv_data_33 : _GEN_32; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_34 = 8'h22 == total_offset ? phv_data_34 : _GEN_33; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_35 = 8'h23 == total_offset ? phv_data_35 : _GEN_34; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_36 = 8'h24 == total_offset ? phv_data_36 : _GEN_35; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_37 = 8'h25 == total_offset ? phv_data_37 : _GEN_36; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_38 = 8'h26 == total_offset ? phv_data_38 : _GEN_37; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_39 = 8'h27 == total_offset ? phv_data_39 : _GEN_38; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_40 = 8'h28 == total_offset ? phv_data_40 : _GEN_39; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_41 = 8'h29 == total_offset ? phv_data_41 : _GEN_40; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_42 = 8'h2a == total_offset ? phv_data_42 : _GEN_41; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_43 = 8'h2b == total_offset ? phv_data_43 : _GEN_42; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_44 = 8'h2c == total_offset ? phv_data_44 : _GEN_43; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_45 = 8'h2d == total_offset ? phv_data_45 : _GEN_44; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_46 = 8'h2e == total_offset ? phv_data_46 : _GEN_45; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_47 = 8'h2f == total_offset ? phv_data_47 : _GEN_46; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_48 = 8'h30 == total_offset ? phv_data_48 : _GEN_47; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_49 = 8'h31 == total_offset ? phv_data_49 : _GEN_48; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_50 = 8'h32 == total_offset ? phv_data_50 : _GEN_49; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_51 = 8'h33 == total_offset ? phv_data_51 : _GEN_50; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_52 = 8'h34 == total_offset ? phv_data_52 : _GEN_51; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_53 = 8'h35 == total_offset ? phv_data_53 : _GEN_52; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_54 = 8'h36 == total_offset ? phv_data_54 : _GEN_53; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_55 = 8'h37 == total_offset ? phv_data_55 : _GEN_54; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_56 = 8'h38 == total_offset ? phv_data_56 : _GEN_55; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_57 = 8'h39 == total_offset ? phv_data_57 : _GEN_56; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_58 = 8'h3a == total_offset ? phv_data_58 : _GEN_57; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_59 = 8'h3b == total_offset ? phv_data_59 : _GEN_58; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_60 = 8'h3c == total_offset ? phv_data_60 : _GEN_59; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_61 = 8'h3d == total_offset ? phv_data_61 : _GEN_60; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_62 = 8'h3e == total_offset ? phv_data_62 : _GEN_61; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_63 = 8'h3f == total_offset ? phv_data_63 : _GEN_62; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_64 = 8'h40 == total_offset ? phv_data_64 : _GEN_63; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_65 = 8'h41 == total_offset ? phv_data_65 : _GEN_64; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_66 = 8'h42 == total_offset ? phv_data_66 : _GEN_65; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_67 = 8'h43 == total_offset ? phv_data_67 : _GEN_66; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_68 = 8'h44 == total_offset ? phv_data_68 : _GEN_67; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_69 = 8'h45 == total_offset ? phv_data_69 : _GEN_68; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_70 = 8'h46 == total_offset ? phv_data_70 : _GEN_69; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_71 = 8'h47 == total_offset ? phv_data_71 : _GEN_70; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_72 = 8'h48 == total_offset ? phv_data_72 : _GEN_71; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_73 = 8'h49 == total_offset ? phv_data_73 : _GEN_72; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_74 = 8'h4a == total_offset ? phv_data_74 : _GEN_73; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_75 = 8'h4b == total_offset ? phv_data_75 : _GEN_74; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_76 = 8'h4c == total_offset ? phv_data_76 : _GEN_75; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_77 = 8'h4d == total_offset ? phv_data_77 : _GEN_76; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_78 = 8'h4e == total_offset ? phv_data_78 : _GEN_77; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_79 = 8'h4f == total_offset ? phv_data_79 : _GEN_78; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_80 = 8'h50 == total_offset ? phv_data_80 : _GEN_79; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_81 = 8'h51 == total_offset ? phv_data_81 : _GEN_80; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_82 = 8'h52 == total_offset ? phv_data_82 : _GEN_81; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_83 = 8'h53 == total_offset ? phv_data_83 : _GEN_82; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_84 = 8'h54 == total_offset ? phv_data_84 : _GEN_83; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_85 = 8'h55 == total_offset ? phv_data_85 : _GEN_84; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_86 = 8'h56 == total_offset ? phv_data_86 : _GEN_85; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_87 = 8'h57 == total_offset ? phv_data_87 : _GEN_86; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_88 = 8'h58 == total_offset ? phv_data_88 : _GEN_87; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_89 = 8'h59 == total_offset ? phv_data_89 : _GEN_88; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_90 = 8'h5a == total_offset ? phv_data_90 : _GEN_89; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_91 = 8'h5b == total_offset ? phv_data_91 : _GEN_90; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_92 = 8'h5c == total_offset ? phv_data_92 : _GEN_91; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_93 = 8'h5d == total_offset ? phv_data_93 : _GEN_92; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_94 = 8'h5e == total_offset ? phv_data_94 : _GEN_93; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_95 = 8'h5f == total_offset ? phv_data_95 : _GEN_94; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_96 = 8'h60 == total_offset ? phv_data_96 : _GEN_95; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_97 = 8'h61 == total_offset ? phv_data_97 : _GEN_96; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_98 = 8'h62 == total_offset ? phv_data_98 : _GEN_97; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_99 = 8'h63 == total_offset ? phv_data_99 : _GEN_98; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_100 = 8'h64 == total_offset ? phv_data_100 : _GEN_99; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_101 = 8'h65 == total_offset ? phv_data_101 : _GEN_100; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_102 = 8'h66 == total_offset ? phv_data_102 : _GEN_101; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_103 = 8'h67 == total_offset ? phv_data_103 : _GEN_102; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_104 = 8'h68 == total_offset ? phv_data_104 : _GEN_103; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_105 = 8'h69 == total_offset ? phv_data_105 : _GEN_104; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_106 = 8'h6a == total_offset ? phv_data_106 : _GEN_105; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_107 = 8'h6b == total_offset ? phv_data_107 : _GEN_106; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_108 = 8'h6c == total_offset ? phv_data_108 : _GEN_107; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_109 = 8'h6d == total_offset ? phv_data_109 : _GEN_108; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_110 = 8'h6e == total_offset ? phv_data_110 : _GEN_109; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_111 = 8'h6f == total_offset ? phv_data_111 : _GEN_110; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_112 = 8'h70 == total_offset ? phv_data_112 : _GEN_111; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_113 = 8'h71 == total_offset ? phv_data_113 : _GEN_112; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_114 = 8'h72 == total_offset ? phv_data_114 : _GEN_113; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_115 = 8'h73 == total_offset ? phv_data_115 : _GEN_114; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_116 = 8'h74 == total_offset ? phv_data_116 : _GEN_115; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_117 = 8'h75 == total_offset ? phv_data_117 : _GEN_116; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_118 = 8'h76 == total_offset ? phv_data_118 : _GEN_117; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_119 = 8'h77 == total_offset ? phv_data_119 : _GEN_118; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_120 = 8'h78 == total_offset ? phv_data_120 : _GEN_119; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_121 = 8'h79 == total_offset ? phv_data_121 : _GEN_120; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_122 = 8'h7a == total_offset ? phv_data_122 : _GEN_121; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_123 = 8'h7b == total_offset ? phv_data_123 : _GEN_122; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_124 = 8'h7c == total_offset ? phv_data_124 : _GEN_123; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_125 = 8'h7d == total_offset ? phv_data_125 : _GEN_124; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_126 = 8'h7e == total_offset ? phv_data_126 : _GEN_125; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_127 = 8'h7f == total_offset ? phv_data_127 : _GEN_126; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_128 = 8'h80 == total_offset ? phv_data_128 : _GEN_127; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_129 = 8'h81 == total_offset ? phv_data_129 : _GEN_128; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_130 = 8'h82 == total_offset ? phv_data_130 : _GEN_129; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_131 = 8'h83 == total_offset ? phv_data_131 : _GEN_130; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_132 = 8'h84 == total_offset ? phv_data_132 : _GEN_131; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_133 = 8'h85 == total_offset ? phv_data_133 : _GEN_132; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_134 = 8'h86 == total_offset ? phv_data_134 : _GEN_133; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_135 = 8'h87 == total_offset ? phv_data_135 : _GEN_134; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_136 = 8'h88 == total_offset ? phv_data_136 : _GEN_135; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_137 = 8'h89 == total_offset ? phv_data_137 : _GEN_136; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_138 = 8'h8a == total_offset ? phv_data_138 : _GEN_137; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_139 = 8'h8b == total_offset ? phv_data_139 : _GEN_138; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_140 = 8'h8c == total_offset ? phv_data_140 : _GEN_139; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_141 = 8'h8d == total_offset ? phv_data_141 : _GEN_140; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_142 = 8'h8e == total_offset ? phv_data_142 : _GEN_141; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_143 = 8'h8f == total_offset ? phv_data_143 : _GEN_142; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_144 = 8'h90 == total_offset ? phv_data_144 : _GEN_143; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_145 = 8'h91 == total_offset ? phv_data_145 : _GEN_144; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_146 = 8'h92 == total_offset ? phv_data_146 : _GEN_145; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_147 = 8'h93 == total_offset ? phv_data_147 : _GEN_146; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_148 = 8'h94 == total_offset ? phv_data_148 : _GEN_147; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_149 = 8'h95 == total_offset ? phv_data_149 : _GEN_148; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_150 = 8'h96 == total_offset ? phv_data_150 : _GEN_149; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_151 = 8'h97 == total_offset ? phv_data_151 : _GEN_150; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_152 = 8'h98 == total_offset ? phv_data_152 : _GEN_151; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_153 = 8'h99 == total_offset ? phv_data_153 : _GEN_152; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_154 = 8'h9a == total_offset ? phv_data_154 : _GEN_153; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_155 = 8'h9b == total_offset ? phv_data_155 : _GEN_154; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_156 = 8'h9c == total_offset ? phv_data_156 : _GEN_155; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_157 = 8'h9d == total_offset ? phv_data_157 : _GEN_156; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_158 = 8'h9e == total_offset ? phv_data_158 : _GEN_157; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes__3 = 8'h9f == total_offset ? phv_data_159 : _GEN_158; // @[executor.scala 197:66 executor.scala 197:66]
  wire  _mask_3_T_3 = ending == 2'h0; // @[executor.scala 199:88]
  wire  mask__3 = 2'h0 >= offset_0[1:0] & (2'h0 < ending | ending == 2'h0); // @[executor.scala 199:56]
  wire [7:0] total_offset_1 = {total_offset_hi,2'h1}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_161 = 8'h1 == total_offset_1 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_162 = 8'h2 == total_offset_1 ? phv_data_2 : _GEN_161; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_163 = 8'h3 == total_offset_1 ? phv_data_3 : _GEN_162; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_164 = 8'h4 == total_offset_1 ? phv_data_4 : _GEN_163; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_165 = 8'h5 == total_offset_1 ? phv_data_5 : _GEN_164; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_166 = 8'h6 == total_offset_1 ? phv_data_6 : _GEN_165; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_167 = 8'h7 == total_offset_1 ? phv_data_7 : _GEN_166; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_168 = 8'h8 == total_offset_1 ? phv_data_8 : _GEN_167; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_169 = 8'h9 == total_offset_1 ? phv_data_9 : _GEN_168; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_170 = 8'ha == total_offset_1 ? phv_data_10 : _GEN_169; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_171 = 8'hb == total_offset_1 ? phv_data_11 : _GEN_170; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_172 = 8'hc == total_offset_1 ? phv_data_12 : _GEN_171; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_173 = 8'hd == total_offset_1 ? phv_data_13 : _GEN_172; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_174 = 8'he == total_offset_1 ? phv_data_14 : _GEN_173; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_175 = 8'hf == total_offset_1 ? phv_data_15 : _GEN_174; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_176 = 8'h10 == total_offset_1 ? phv_data_16 : _GEN_175; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_177 = 8'h11 == total_offset_1 ? phv_data_17 : _GEN_176; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_178 = 8'h12 == total_offset_1 ? phv_data_18 : _GEN_177; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_179 = 8'h13 == total_offset_1 ? phv_data_19 : _GEN_178; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_180 = 8'h14 == total_offset_1 ? phv_data_20 : _GEN_179; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_181 = 8'h15 == total_offset_1 ? phv_data_21 : _GEN_180; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_182 = 8'h16 == total_offset_1 ? phv_data_22 : _GEN_181; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_183 = 8'h17 == total_offset_1 ? phv_data_23 : _GEN_182; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_184 = 8'h18 == total_offset_1 ? phv_data_24 : _GEN_183; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_185 = 8'h19 == total_offset_1 ? phv_data_25 : _GEN_184; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_186 = 8'h1a == total_offset_1 ? phv_data_26 : _GEN_185; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_187 = 8'h1b == total_offset_1 ? phv_data_27 : _GEN_186; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_188 = 8'h1c == total_offset_1 ? phv_data_28 : _GEN_187; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_189 = 8'h1d == total_offset_1 ? phv_data_29 : _GEN_188; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_190 = 8'h1e == total_offset_1 ? phv_data_30 : _GEN_189; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_191 = 8'h1f == total_offset_1 ? phv_data_31 : _GEN_190; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_192 = 8'h20 == total_offset_1 ? phv_data_32 : _GEN_191; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_193 = 8'h21 == total_offset_1 ? phv_data_33 : _GEN_192; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_194 = 8'h22 == total_offset_1 ? phv_data_34 : _GEN_193; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_195 = 8'h23 == total_offset_1 ? phv_data_35 : _GEN_194; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_196 = 8'h24 == total_offset_1 ? phv_data_36 : _GEN_195; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_197 = 8'h25 == total_offset_1 ? phv_data_37 : _GEN_196; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_198 = 8'h26 == total_offset_1 ? phv_data_38 : _GEN_197; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_199 = 8'h27 == total_offset_1 ? phv_data_39 : _GEN_198; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_200 = 8'h28 == total_offset_1 ? phv_data_40 : _GEN_199; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_201 = 8'h29 == total_offset_1 ? phv_data_41 : _GEN_200; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_202 = 8'h2a == total_offset_1 ? phv_data_42 : _GEN_201; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_203 = 8'h2b == total_offset_1 ? phv_data_43 : _GEN_202; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_204 = 8'h2c == total_offset_1 ? phv_data_44 : _GEN_203; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_205 = 8'h2d == total_offset_1 ? phv_data_45 : _GEN_204; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_206 = 8'h2e == total_offset_1 ? phv_data_46 : _GEN_205; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_207 = 8'h2f == total_offset_1 ? phv_data_47 : _GEN_206; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_208 = 8'h30 == total_offset_1 ? phv_data_48 : _GEN_207; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_209 = 8'h31 == total_offset_1 ? phv_data_49 : _GEN_208; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_210 = 8'h32 == total_offset_1 ? phv_data_50 : _GEN_209; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_211 = 8'h33 == total_offset_1 ? phv_data_51 : _GEN_210; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_212 = 8'h34 == total_offset_1 ? phv_data_52 : _GEN_211; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_213 = 8'h35 == total_offset_1 ? phv_data_53 : _GEN_212; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_214 = 8'h36 == total_offset_1 ? phv_data_54 : _GEN_213; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_215 = 8'h37 == total_offset_1 ? phv_data_55 : _GEN_214; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_216 = 8'h38 == total_offset_1 ? phv_data_56 : _GEN_215; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_217 = 8'h39 == total_offset_1 ? phv_data_57 : _GEN_216; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_218 = 8'h3a == total_offset_1 ? phv_data_58 : _GEN_217; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_219 = 8'h3b == total_offset_1 ? phv_data_59 : _GEN_218; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_220 = 8'h3c == total_offset_1 ? phv_data_60 : _GEN_219; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_221 = 8'h3d == total_offset_1 ? phv_data_61 : _GEN_220; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_222 = 8'h3e == total_offset_1 ? phv_data_62 : _GEN_221; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_223 = 8'h3f == total_offset_1 ? phv_data_63 : _GEN_222; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_224 = 8'h40 == total_offset_1 ? phv_data_64 : _GEN_223; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_225 = 8'h41 == total_offset_1 ? phv_data_65 : _GEN_224; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_226 = 8'h42 == total_offset_1 ? phv_data_66 : _GEN_225; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_227 = 8'h43 == total_offset_1 ? phv_data_67 : _GEN_226; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_228 = 8'h44 == total_offset_1 ? phv_data_68 : _GEN_227; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_229 = 8'h45 == total_offset_1 ? phv_data_69 : _GEN_228; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_230 = 8'h46 == total_offset_1 ? phv_data_70 : _GEN_229; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_231 = 8'h47 == total_offset_1 ? phv_data_71 : _GEN_230; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_232 = 8'h48 == total_offset_1 ? phv_data_72 : _GEN_231; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_233 = 8'h49 == total_offset_1 ? phv_data_73 : _GEN_232; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_234 = 8'h4a == total_offset_1 ? phv_data_74 : _GEN_233; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_235 = 8'h4b == total_offset_1 ? phv_data_75 : _GEN_234; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_236 = 8'h4c == total_offset_1 ? phv_data_76 : _GEN_235; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_237 = 8'h4d == total_offset_1 ? phv_data_77 : _GEN_236; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_238 = 8'h4e == total_offset_1 ? phv_data_78 : _GEN_237; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_239 = 8'h4f == total_offset_1 ? phv_data_79 : _GEN_238; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_240 = 8'h50 == total_offset_1 ? phv_data_80 : _GEN_239; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_241 = 8'h51 == total_offset_1 ? phv_data_81 : _GEN_240; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_242 = 8'h52 == total_offset_1 ? phv_data_82 : _GEN_241; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_243 = 8'h53 == total_offset_1 ? phv_data_83 : _GEN_242; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_244 = 8'h54 == total_offset_1 ? phv_data_84 : _GEN_243; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_245 = 8'h55 == total_offset_1 ? phv_data_85 : _GEN_244; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_246 = 8'h56 == total_offset_1 ? phv_data_86 : _GEN_245; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_247 = 8'h57 == total_offset_1 ? phv_data_87 : _GEN_246; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_248 = 8'h58 == total_offset_1 ? phv_data_88 : _GEN_247; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_249 = 8'h59 == total_offset_1 ? phv_data_89 : _GEN_248; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_250 = 8'h5a == total_offset_1 ? phv_data_90 : _GEN_249; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_251 = 8'h5b == total_offset_1 ? phv_data_91 : _GEN_250; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_252 = 8'h5c == total_offset_1 ? phv_data_92 : _GEN_251; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_253 = 8'h5d == total_offset_1 ? phv_data_93 : _GEN_252; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_254 = 8'h5e == total_offset_1 ? phv_data_94 : _GEN_253; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_255 = 8'h5f == total_offset_1 ? phv_data_95 : _GEN_254; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_256 = 8'h60 == total_offset_1 ? phv_data_96 : _GEN_255; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_257 = 8'h61 == total_offset_1 ? phv_data_97 : _GEN_256; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_258 = 8'h62 == total_offset_1 ? phv_data_98 : _GEN_257; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_259 = 8'h63 == total_offset_1 ? phv_data_99 : _GEN_258; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_260 = 8'h64 == total_offset_1 ? phv_data_100 : _GEN_259; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_261 = 8'h65 == total_offset_1 ? phv_data_101 : _GEN_260; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_262 = 8'h66 == total_offset_1 ? phv_data_102 : _GEN_261; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_263 = 8'h67 == total_offset_1 ? phv_data_103 : _GEN_262; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_264 = 8'h68 == total_offset_1 ? phv_data_104 : _GEN_263; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_265 = 8'h69 == total_offset_1 ? phv_data_105 : _GEN_264; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_266 = 8'h6a == total_offset_1 ? phv_data_106 : _GEN_265; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_267 = 8'h6b == total_offset_1 ? phv_data_107 : _GEN_266; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_268 = 8'h6c == total_offset_1 ? phv_data_108 : _GEN_267; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_269 = 8'h6d == total_offset_1 ? phv_data_109 : _GEN_268; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_270 = 8'h6e == total_offset_1 ? phv_data_110 : _GEN_269; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_271 = 8'h6f == total_offset_1 ? phv_data_111 : _GEN_270; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_272 = 8'h70 == total_offset_1 ? phv_data_112 : _GEN_271; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_273 = 8'h71 == total_offset_1 ? phv_data_113 : _GEN_272; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_274 = 8'h72 == total_offset_1 ? phv_data_114 : _GEN_273; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_275 = 8'h73 == total_offset_1 ? phv_data_115 : _GEN_274; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_276 = 8'h74 == total_offset_1 ? phv_data_116 : _GEN_275; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_277 = 8'h75 == total_offset_1 ? phv_data_117 : _GEN_276; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_278 = 8'h76 == total_offset_1 ? phv_data_118 : _GEN_277; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_279 = 8'h77 == total_offset_1 ? phv_data_119 : _GEN_278; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_280 = 8'h78 == total_offset_1 ? phv_data_120 : _GEN_279; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_281 = 8'h79 == total_offset_1 ? phv_data_121 : _GEN_280; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_282 = 8'h7a == total_offset_1 ? phv_data_122 : _GEN_281; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_283 = 8'h7b == total_offset_1 ? phv_data_123 : _GEN_282; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_284 = 8'h7c == total_offset_1 ? phv_data_124 : _GEN_283; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_285 = 8'h7d == total_offset_1 ? phv_data_125 : _GEN_284; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_286 = 8'h7e == total_offset_1 ? phv_data_126 : _GEN_285; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_287 = 8'h7f == total_offset_1 ? phv_data_127 : _GEN_286; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_288 = 8'h80 == total_offset_1 ? phv_data_128 : _GEN_287; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_289 = 8'h81 == total_offset_1 ? phv_data_129 : _GEN_288; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_290 = 8'h82 == total_offset_1 ? phv_data_130 : _GEN_289; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_291 = 8'h83 == total_offset_1 ? phv_data_131 : _GEN_290; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_292 = 8'h84 == total_offset_1 ? phv_data_132 : _GEN_291; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_293 = 8'h85 == total_offset_1 ? phv_data_133 : _GEN_292; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_294 = 8'h86 == total_offset_1 ? phv_data_134 : _GEN_293; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_295 = 8'h87 == total_offset_1 ? phv_data_135 : _GEN_294; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_296 = 8'h88 == total_offset_1 ? phv_data_136 : _GEN_295; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_297 = 8'h89 == total_offset_1 ? phv_data_137 : _GEN_296; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_298 = 8'h8a == total_offset_1 ? phv_data_138 : _GEN_297; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_299 = 8'h8b == total_offset_1 ? phv_data_139 : _GEN_298; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_300 = 8'h8c == total_offset_1 ? phv_data_140 : _GEN_299; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_301 = 8'h8d == total_offset_1 ? phv_data_141 : _GEN_300; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_302 = 8'h8e == total_offset_1 ? phv_data_142 : _GEN_301; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_303 = 8'h8f == total_offset_1 ? phv_data_143 : _GEN_302; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_304 = 8'h90 == total_offset_1 ? phv_data_144 : _GEN_303; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_305 = 8'h91 == total_offset_1 ? phv_data_145 : _GEN_304; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_306 = 8'h92 == total_offset_1 ? phv_data_146 : _GEN_305; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_307 = 8'h93 == total_offset_1 ? phv_data_147 : _GEN_306; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_308 = 8'h94 == total_offset_1 ? phv_data_148 : _GEN_307; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_309 = 8'h95 == total_offset_1 ? phv_data_149 : _GEN_308; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_310 = 8'h96 == total_offset_1 ? phv_data_150 : _GEN_309; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_311 = 8'h97 == total_offset_1 ? phv_data_151 : _GEN_310; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_312 = 8'h98 == total_offset_1 ? phv_data_152 : _GEN_311; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_313 = 8'h99 == total_offset_1 ? phv_data_153 : _GEN_312; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_314 = 8'h9a == total_offset_1 ? phv_data_154 : _GEN_313; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_315 = 8'h9b == total_offset_1 ? phv_data_155 : _GEN_314; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_316 = 8'h9c == total_offset_1 ? phv_data_156 : _GEN_315; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_317 = 8'h9d == total_offset_1 ? phv_data_157 : _GEN_316; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_318 = 8'h9e == total_offset_1 ? phv_data_158 : _GEN_317; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes__2 = 8'h9f == total_offset_1 ? phv_data_159 : _GEN_318; // @[executor.scala 197:66 executor.scala 197:66]
  wire  mask__2 = 2'h1 >= offset_0[1:0] & (2'h1 < ending | ending == 2'h0); // @[executor.scala 199:56]
  wire [7:0] total_offset_2 = {total_offset_hi,2'h2}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_321 = 8'h1 == total_offset_2 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_322 = 8'h2 == total_offset_2 ? phv_data_2 : _GEN_321; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_323 = 8'h3 == total_offset_2 ? phv_data_3 : _GEN_322; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_324 = 8'h4 == total_offset_2 ? phv_data_4 : _GEN_323; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_325 = 8'h5 == total_offset_2 ? phv_data_5 : _GEN_324; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_326 = 8'h6 == total_offset_2 ? phv_data_6 : _GEN_325; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_327 = 8'h7 == total_offset_2 ? phv_data_7 : _GEN_326; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_328 = 8'h8 == total_offset_2 ? phv_data_8 : _GEN_327; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_329 = 8'h9 == total_offset_2 ? phv_data_9 : _GEN_328; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_330 = 8'ha == total_offset_2 ? phv_data_10 : _GEN_329; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_331 = 8'hb == total_offset_2 ? phv_data_11 : _GEN_330; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_332 = 8'hc == total_offset_2 ? phv_data_12 : _GEN_331; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_333 = 8'hd == total_offset_2 ? phv_data_13 : _GEN_332; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_334 = 8'he == total_offset_2 ? phv_data_14 : _GEN_333; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_335 = 8'hf == total_offset_2 ? phv_data_15 : _GEN_334; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_336 = 8'h10 == total_offset_2 ? phv_data_16 : _GEN_335; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_337 = 8'h11 == total_offset_2 ? phv_data_17 : _GEN_336; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_338 = 8'h12 == total_offset_2 ? phv_data_18 : _GEN_337; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_339 = 8'h13 == total_offset_2 ? phv_data_19 : _GEN_338; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_340 = 8'h14 == total_offset_2 ? phv_data_20 : _GEN_339; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_341 = 8'h15 == total_offset_2 ? phv_data_21 : _GEN_340; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_342 = 8'h16 == total_offset_2 ? phv_data_22 : _GEN_341; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_343 = 8'h17 == total_offset_2 ? phv_data_23 : _GEN_342; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_344 = 8'h18 == total_offset_2 ? phv_data_24 : _GEN_343; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_345 = 8'h19 == total_offset_2 ? phv_data_25 : _GEN_344; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_346 = 8'h1a == total_offset_2 ? phv_data_26 : _GEN_345; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_347 = 8'h1b == total_offset_2 ? phv_data_27 : _GEN_346; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_348 = 8'h1c == total_offset_2 ? phv_data_28 : _GEN_347; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_349 = 8'h1d == total_offset_2 ? phv_data_29 : _GEN_348; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_350 = 8'h1e == total_offset_2 ? phv_data_30 : _GEN_349; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_351 = 8'h1f == total_offset_2 ? phv_data_31 : _GEN_350; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_352 = 8'h20 == total_offset_2 ? phv_data_32 : _GEN_351; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_353 = 8'h21 == total_offset_2 ? phv_data_33 : _GEN_352; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_354 = 8'h22 == total_offset_2 ? phv_data_34 : _GEN_353; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_355 = 8'h23 == total_offset_2 ? phv_data_35 : _GEN_354; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_356 = 8'h24 == total_offset_2 ? phv_data_36 : _GEN_355; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_357 = 8'h25 == total_offset_2 ? phv_data_37 : _GEN_356; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_358 = 8'h26 == total_offset_2 ? phv_data_38 : _GEN_357; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_359 = 8'h27 == total_offset_2 ? phv_data_39 : _GEN_358; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_360 = 8'h28 == total_offset_2 ? phv_data_40 : _GEN_359; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_361 = 8'h29 == total_offset_2 ? phv_data_41 : _GEN_360; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_362 = 8'h2a == total_offset_2 ? phv_data_42 : _GEN_361; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_363 = 8'h2b == total_offset_2 ? phv_data_43 : _GEN_362; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_364 = 8'h2c == total_offset_2 ? phv_data_44 : _GEN_363; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_365 = 8'h2d == total_offset_2 ? phv_data_45 : _GEN_364; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_366 = 8'h2e == total_offset_2 ? phv_data_46 : _GEN_365; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_367 = 8'h2f == total_offset_2 ? phv_data_47 : _GEN_366; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_368 = 8'h30 == total_offset_2 ? phv_data_48 : _GEN_367; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_369 = 8'h31 == total_offset_2 ? phv_data_49 : _GEN_368; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_370 = 8'h32 == total_offset_2 ? phv_data_50 : _GEN_369; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_371 = 8'h33 == total_offset_2 ? phv_data_51 : _GEN_370; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_372 = 8'h34 == total_offset_2 ? phv_data_52 : _GEN_371; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_373 = 8'h35 == total_offset_2 ? phv_data_53 : _GEN_372; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_374 = 8'h36 == total_offset_2 ? phv_data_54 : _GEN_373; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_375 = 8'h37 == total_offset_2 ? phv_data_55 : _GEN_374; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_376 = 8'h38 == total_offset_2 ? phv_data_56 : _GEN_375; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_377 = 8'h39 == total_offset_2 ? phv_data_57 : _GEN_376; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_378 = 8'h3a == total_offset_2 ? phv_data_58 : _GEN_377; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_379 = 8'h3b == total_offset_2 ? phv_data_59 : _GEN_378; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_380 = 8'h3c == total_offset_2 ? phv_data_60 : _GEN_379; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_381 = 8'h3d == total_offset_2 ? phv_data_61 : _GEN_380; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_382 = 8'h3e == total_offset_2 ? phv_data_62 : _GEN_381; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_383 = 8'h3f == total_offset_2 ? phv_data_63 : _GEN_382; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_384 = 8'h40 == total_offset_2 ? phv_data_64 : _GEN_383; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_385 = 8'h41 == total_offset_2 ? phv_data_65 : _GEN_384; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_386 = 8'h42 == total_offset_2 ? phv_data_66 : _GEN_385; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_387 = 8'h43 == total_offset_2 ? phv_data_67 : _GEN_386; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_388 = 8'h44 == total_offset_2 ? phv_data_68 : _GEN_387; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_389 = 8'h45 == total_offset_2 ? phv_data_69 : _GEN_388; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_390 = 8'h46 == total_offset_2 ? phv_data_70 : _GEN_389; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_391 = 8'h47 == total_offset_2 ? phv_data_71 : _GEN_390; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_392 = 8'h48 == total_offset_2 ? phv_data_72 : _GEN_391; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_393 = 8'h49 == total_offset_2 ? phv_data_73 : _GEN_392; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_394 = 8'h4a == total_offset_2 ? phv_data_74 : _GEN_393; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_395 = 8'h4b == total_offset_2 ? phv_data_75 : _GEN_394; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_396 = 8'h4c == total_offset_2 ? phv_data_76 : _GEN_395; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_397 = 8'h4d == total_offset_2 ? phv_data_77 : _GEN_396; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_398 = 8'h4e == total_offset_2 ? phv_data_78 : _GEN_397; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_399 = 8'h4f == total_offset_2 ? phv_data_79 : _GEN_398; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_400 = 8'h50 == total_offset_2 ? phv_data_80 : _GEN_399; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_401 = 8'h51 == total_offset_2 ? phv_data_81 : _GEN_400; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_402 = 8'h52 == total_offset_2 ? phv_data_82 : _GEN_401; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_403 = 8'h53 == total_offset_2 ? phv_data_83 : _GEN_402; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_404 = 8'h54 == total_offset_2 ? phv_data_84 : _GEN_403; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_405 = 8'h55 == total_offset_2 ? phv_data_85 : _GEN_404; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_406 = 8'h56 == total_offset_2 ? phv_data_86 : _GEN_405; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_407 = 8'h57 == total_offset_2 ? phv_data_87 : _GEN_406; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_408 = 8'h58 == total_offset_2 ? phv_data_88 : _GEN_407; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_409 = 8'h59 == total_offset_2 ? phv_data_89 : _GEN_408; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_410 = 8'h5a == total_offset_2 ? phv_data_90 : _GEN_409; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_411 = 8'h5b == total_offset_2 ? phv_data_91 : _GEN_410; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_412 = 8'h5c == total_offset_2 ? phv_data_92 : _GEN_411; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_413 = 8'h5d == total_offset_2 ? phv_data_93 : _GEN_412; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_414 = 8'h5e == total_offset_2 ? phv_data_94 : _GEN_413; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_415 = 8'h5f == total_offset_2 ? phv_data_95 : _GEN_414; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_416 = 8'h60 == total_offset_2 ? phv_data_96 : _GEN_415; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_417 = 8'h61 == total_offset_2 ? phv_data_97 : _GEN_416; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_418 = 8'h62 == total_offset_2 ? phv_data_98 : _GEN_417; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_419 = 8'h63 == total_offset_2 ? phv_data_99 : _GEN_418; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_420 = 8'h64 == total_offset_2 ? phv_data_100 : _GEN_419; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_421 = 8'h65 == total_offset_2 ? phv_data_101 : _GEN_420; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_422 = 8'h66 == total_offset_2 ? phv_data_102 : _GEN_421; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_423 = 8'h67 == total_offset_2 ? phv_data_103 : _GEN_422; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_424 = 8'h68 == total_offset_2 ? phv_data_104 : _GEN_423; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_425 = 8'h69 == total_offset_2 ? phv_data_105 : _GEN_424; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_426 = 8'h6a == total_offset_2 ? phv_data_106 : _GEN_425; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_427 = 8'h6b == total_offset_2 ? phv_data_107 : _GEN_426; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_428 = 8'h6c == total_offset_2 ? phv_data_108 : _GEN_427; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_429 = 8'h6d == total_offset_2 ? phv_data_109 : _GEN_428; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_430 = 8'h6e == total_offset_2 ? phv_data_110 : _GEN_429; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_431 = 8'h6f == total_offset_2 ? phv_data_111 : _GEN_430; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_432 = 8'h70 == total_offset_2 ? phv_data_112 : _GEN_431; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_433 = 8'h71 == total_offset_2 ? phv_data_113 : _GEN_432; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_434 = 8'h72 == total_offset_2 ? phv_data_114 : _GEN_433; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_435 = 8'h73 == total_offset_2 ? phv_data_115 : _GEN_434; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_436 = 8'h74 == total_offset_2 ? phv_data_116 : _GEN_435; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_437 = 8'h75 == total_offset_2 ? phv_data_117 : _GEN_436; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_438 = 8'h76 == total_offset_2 ? phv_data_118 : _GEN_437; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_439 = 8'h77 == total_offset_2 ? phv_data_119 : _GEN_438; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_440 = 8'h78 == total_offset_2 ? phv_data_120 : _GEN_439; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_441 = 8'h79 == total_offset_2 ? phv_data_121 : _GEN_440; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_442 = 8'h7a == total_offset_2 ? phv_data_122 : _GEN_441; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_443 = 8'h7b == total_offset_2 ? phv_data_123 : _GEN_442; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_444 = 8'h7c == total_offset_2 ? phv_data_124 : _GEN_443; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_445 = 8'h7d == total_offset_2 ? phv_data_125 : _GEN_444; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_446 = 8'h7e == total_offset_2 ? phv_data_126 : _GEN_445; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_447 = 8'h7f == total_offset_2 ? phv_data_127 : _GEN_446; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_448 = 8'h80 == total_offset_2 ? phv_data_128 : _GEN_447; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_449 = 8'h81 == total_offset_2 ? phv_data_129 : _GEN_448; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_450 = 8'h82 == total_offset_2 ? phv_data_130 : _GEN_449; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_451 = 8'h83 == total_offset_2 ? phv_data_131 : _GEN_450; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_452 = 8'h84 == total_offset_2 ? phv_data_132 : _GEN_451; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_453 = 8'h85 == total_offset_2 ? phv_data_133 : _GEN_452; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_454 = 8'h86 == total_offset_2 ? phv_data_134 : _GEN_453; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_455 = 8'h87 == total_offset_2 ? phv_data_135 : _GEN_454; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_456 = 8'h88 == total_offset_2 ? phv_data_136 : _GEN_455; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_457 = 8'h89 == total_offset_2 ? phv_data_137 : _GEN_456; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_458 = 8'h8a == total_offset_2 ? phv_data_138 : _GEN_457; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_459 = 8'h8b == total_offset_2 ? phv_data_139 : _GEN_458; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_460 = 8'h8c == total_offset_2 ? phv_data_140 : _GEN_459; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_461 = 8'h8d == total_offset_2 ? phv_data_141 : _GEN_460; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_462 = 8'h8e == total_offset_2 ? phv_data_142 : _GEN_461; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_463 = 8'h8f == total_offset_2 ? phv_data_143 : _GEN_462; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_464 = 8'h90 == total_offset_2 ? phv_data_144 : _GEN_463; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_465 = 8'h91 == total_offset_2 ? phv_data_145 : _GEN_464; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_466 = 8'h92 == total_offset_2 ? phv_data_146 : _GEN_465; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_467 = 8'h93 == total_offset_2 ? phv_data_147 : _GEN_466; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_468 = 8'h94 == total_offset_2 ? phv_data_148 : _GEN_467; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_469 = 8'h95 == total_offset_2 ? phv_data_149 : _GEN_468; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_470 = 8'h96 == total_offset_2 ? phv_data_150 : _GEN_469; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_471 = 8'h97 == total_offset_2 ? phv_data_151 : _GEN_470; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_472 = 8'h98 == total_offset_2 ? phv_data_152 : _GEN_471; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_473 = 8'h99 == total_offset_2 ? phv_data_153 : _GEN_472; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_474 = 8'h9a == total_offset_2 ? phv_data_154 : _GEN_473; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_475 = 8'h9b == total_offset_2 ? phv_data_155 : _GEN_474; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_476 = 8'h9c == total_offset_2 ? phv_data_156 : _GEN_475; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_477 = 8'h9d == total_offset_2 ? phv_data_157 : _GEN_476; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_478 = 8'h9e == total_offset_2 ? phv_data_158 : _GEN_477; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes__1 = 8'h9f == total_offset_2 ? phv_data_159 : _GEN_478; // @[executor.scala 197:66 executor.scala 197:66]
  wire  mask__1 = 2'h2 >= offset_0[1:0] & (2'h2 < ending | ending == 2'h0); // @[executor.scala 199:56]
  wire [7:0] total_offset_3 = {total_offset_hi,2'h3}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_481 = 8'h1 == total_offset_3 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_482 = 8'h2 == total_offset_3 ? phv_data_2 : _GEN_481; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_483 = 8'h3 == total_offset_3 ? phv_data_3 : _GEN_482; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_484 = 8'h4 == total_offset_3 ? phv_data_4 : _GEN_483; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_485 = 8'h5 == total_offset_3 ? phv_data_5 : _GEN_484; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_486 = 8'h6 == total_offset_3 ? phv_data_6 : _GEN_485; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_487 = 8'h7 == total_offset_3 ? phv_data_7 : _GEN_486; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_488 = 8'h8 == total_offset_3 ? phv_data_8 : _GEN_487; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_489 = 8'h9 == total_offset_3 ? phv_data_9 : _GEN_488; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_490 = 8'ha == total_offset_3 ? phv_data_10 : _GEN_489; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_491 = 8'hb == total_offset_3 ? phv_data_11 : _GEN_490; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_492 = 8'hc == total_offset_3 ? phv_data_12 : _GEN_491; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_493 = 8'hd == total_offset_3 ? phv_data_13 : _GEN_492; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_494 = 8'he == total_offset_3 ? phv_data_14 : _GEN_493; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_495 = 8'hf == total_offset_3 ? phv_data_15 : _GEN_494; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_496 = 8'h10 == total_offset_3 ? phv_data_16 : _GEN_495; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_497 = 8'h11 == total_offset_3 ? phv_data_17 : _GEN_496; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_498 = 8'h12 == total_offset_3 ? phv_data_18 : _GEN_497; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_499 = 8'h13 == total_offset_3 ? phv_data_19 : _GEN_498; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_500 = 8'h14 == total_offset_3 ? phv_data_20 : _GEN_499; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_501 = 8'h15 == total_offset_3 ? phv_data_21 : _GEN_500; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_502 = 8'h16 == total_offset_3 ? phv_data_22 : _GEN_501; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_503 = 8'h17 == total_offset_3 ? phv_data_23 : _GEN_502; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_504 = 8'h18 == total_offset_3 ? phv_data_24 : _GEN_503; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_505 = 8'h19 == total_offset_3 ? phv_data_25 : _GEN_504; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_506 = 8'h1a == total_offset_3 ? phv_data_26 : _GEN_505; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_507 = 8'h1b == total_offset_3 ? phv_data_27 : _GEN_506; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_508 = 8'h1c == total_offset_3 ? phv_data_28 : _GEN_507; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_509 = 8'h1d == total_offset_3 ? phv_data_29 : _GEN_508; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_510 = 8'h1e == total_offset_3 ? phv_data_30 : _GEN_509; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_511 = 8'h1f == total_offset_3 ? phv_data_31 : _GEN_510; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_512 = 8'h20 == total_offset_3 ? phv_data_32 : _GEN_511; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_513 = 8'h21 == total_offset_3 ? phv_data_33 : _GEN_512; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_514 = 8'h22 == total_offset_3 ? phv_data_34 : _GEN_513; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_515 = 8'h23 == total_offset_3 ? phv_data_35 : _GEN_514; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_516 = 8'h24 == total_offset_3 ? phv_data_36 : _GEN_515; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_517 = 8'h25 == total_offset_3 ? phv_data_37 : _GEN_516; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_518 = 8'h26 == total_offset_3 ? phv_data_38 : _GEN_517; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_519 = 8'h27 == total_offset_3 ? phv_data_39 : _GEN_518; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_520 = 8'h28 == total_offset_3 ? phv_data_40 : _GEN_519; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_521 = 8'h29 == total_offset_3 ? phv_data_41 : _GEN_520; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_522 = 8'h2a == total_offset_3 ? phv_data_42 : _GEN_521; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_523 = 8'h2b == total_offset_3 ? phv_data_43 : _GEN_522; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_524 = 8'h2c == total_offset_3 ? phv_data_44 : _GEN_523; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_525 = 8'h2d == total_offset_3 ? phv_data_45 : _GEN_524; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_526 = 8'h2e == total_offset_3 ? phv_data_46 : _GEN_525; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_527 = 8'h2f == total_offset_3 ? phv_data_47 : _GEN_526; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_528 = 8'h30 == total_offset_3 ? phv_data_48 : _GEN_527; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_529 = 8'h31 == total_offset_3 ? phv_data_49 : _GEN_528; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_530 = 8'h32 == total_offset_3 ? phv_data_50 : _GEN_529; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_531 = 8'h33 == total_offset_3 ? phv_data_51 : _GEN_530; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_532 = 8'h34 == total_offset_3 ? phv_data_52 : _GEN_531; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_533 = 8'h35 == total_offset_3 ? phv_data_53 : _GEN_532; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_534 = 8'h36 == total_offset_3 ? phv_data_54 : _GEN_533; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_535 = 8'h37 == total_offset_3 ? phv_data_55 : _GEN_534; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_536 = 8'h38 == total_offset_3 ? phv_data_56 : _GEN_535; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_537 = 8'h39 == total_offset_3 ? phv_data_57 : _GEN_536; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_538 = 8'h3a == total_offset_3 ? phv_data_58 : _GEN_537; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_539 = 8'h3b == total_offset_3 ? phv_data_59 : _GEN_538; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_540 = 8'h3c == total_offset_3 ? phv_data_60 : _GEN_539; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_541 = 8'h3d == total_offset_3 ? phv_data_61 : _GEN_540; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_542 = 8'h3e == total_offset_3 ? phv_data_62 : _GEN_541; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_543 = 8'h3f == total_offset_3 ? phv_data_63 : _GEN_542; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_544 = 8'h40 == total_offset_3 ? phv_data_64 : _GEN_543; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_545 = 8'h41 == total_offset_3 ? phv_data_65 : _GEN_544; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_546 = 8'h42 == total_offset_3 ? phv_data_66 : _GEN_545; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_547 = 8'h43 == total_offset_3 ? phv_data_67 : _GEN_546; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_548 = 8'h44 == total_offset_3 ? phv_data_68 : _GEN_547; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_549 = 8'h45 == total_offset_3 ? phv_data_69 : _GEN_548; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_550 = 8'h46 == total_offset_3 ? phv_data_70 : _GEN_549; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_551 = 8'h47 == total_offset_3 ? phv_data_71 : _GEN_550; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_552 = 8'h48 == total_offset_3 ? phv_data_72 : _GEN_551; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_553 = 8'h49 == total_offset_3 ? phv_data_73 : _GEN_552; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_554 = 8'h4a == total_offset_3 ? phv_data_74 : _GEN_553; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_555 = 8'h4b == total_offset_3 ? phv_data_75 : _GEN_554; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_556 = 8'h4c == total_offset_3 ? phv_data_76 : _GEN_555; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_557 = 8'h4d == total_offset_3 ? phv_data_77 : _GEN_556; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_558 = 8'h4e == total_offset_3 ? phv_data_78 : _GEN_557; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_559 = 8'h4f == total_offset_3 ? phv_data_79 : _GEN_558; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_560 = 8'h50 == total_offset_3 ? phv_data_80 : _GEN_559; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_561 = 8'h51 == total_offset_3 ? phv_data_81 : _GEN_560; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_562 = 8'h52 == total_offset_3 ? phv_data_82 : _GEN_561; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_563 = 8'h53 == total_offset_3 ? phv_data_83 : _GEN_562; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_564 = 8'h54 == total_offset_3 ? phv_data_84 : _GEN_563; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_565 = 8'h55 == total_offset_3 ? phv_data_85 : _GEN_564; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_566 = 8'h56 == total_offset_3 ? phv_data_86 : _GEN_565; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_567 = 8'h57 == total_offset_3 ? phv_data_87 : _GEN_566; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_568 = 8'h58 == total_offset_3 ? phv_data_88 : _GEN_567; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_569 = 8'h59 == total_offset_3 ? phv_data_89 : _GEN_568; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_570 = 8'h5a == total_offset_3 ? phv_data_90 : _GEN_569; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_571 = 8'h5b == total_offset_3 ? phv_data_91 : _GEN_570; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_572 = 8'h5c == total_offset_3 ? phv_data_92 : _GEN_571; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_573 = 8'h5d == total_offset_3 ? phv_data_93 : _GEN_572; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_574 = 8'h5e == total_offset_3 ? phv_data_94 : _GEN_573; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_575 = 8'h5f == total_offset_3 ? phv_data_95 : _GEN_574; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_576 = 8'h60 == total_offset_3 ? phv_data_96 : _GEN_575; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_577 = 8'h61 == total_offset_3 ? phv_data_97 : _GEN_576; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_578 = 8'h62 == total_offset_3 ? phv_data_98 : _GEN_577; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_579 = 8'h63 == total_offset_3 ? phv_data_99 : _GEN_578; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_580 = 8'h64 == total_offset_3 ? phv_data_100 : _GEN_579; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_581 = 8'h65 == total_offset_3 ? phv_data_101 : _GEN_580; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_582 = 8'h66 == total_offset_3 ? phv_data_102 : _GEN_581; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_583 = 8'h67 == total_offset_3 ? phv_data_103 : _GEN_582; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_584 = 8'h68 == total_offset_3 ? phv_data_104 : _GEN_583; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_585 = 8'h69 == total_offset_3 ? phv_data_105 : _GEN_584; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_586 = 8'h6a == total_offset_3 ? phv_data_106 : _GEN_585; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_587 = 8'h6b == total_offset_3 ? phv_data_107 : _GEN_586; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_588 = 8'h6c == total_offset_3 ? phv_data_108 : _GEN_587; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_589 = 8'h6d == total_offset_3 ? phv_data_109 : _GEN_588; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_590 = 8'h6e == total_offset_3 ? phv_data_110 : _GEN_589; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_591 = 8'h6f == total_offset_3 ? phv_data_111 : _GEN_590; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_592 = 8'h70 == total_offset_3 ? phv_data_112 : _GEN_591; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_593 = 8'h71 == total_offset_3 ? phv_data_113 : _GEN_592; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_594 = 8'h72 == total_offset_3 ? phv_data_114 : _GEN_593; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_595 = 8'h73 == total_offset_3 ? phv_data_115 : _GEN_594; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_596 = 8'h74 == total_offset_3 ? phv_data_116 : _GEN_595; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_597 = 8'h75 == total_offset_3 ? phv_data_117 : _GEN_596; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_598 = 8'h76 == total_offset_3 ? phv_data_118 : _GEN_597; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_599 = 8'h77 == total_offset_3 ? phv_data_119 : _GEN_598; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_600 = 8'h78 == total_offset_3 ? phv_data_120 : _GEN_599; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_601 = 8'h79 == total_offset_3 ? phv_data_121 : _GEN_600; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_602 = 8'h7a == total_offset_3 ? phv_data_122 : _GEN_601; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_603 = 8'h7b == total_offset_3 ? phv_data_123 : _GEN_602; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_604 = 8'h7c == total_offset_3 ? phv_data_124 : _GEN_603; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_605 = 8'h7d == total_offset_3 ? phv_data_125 : _GEN_604; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_606 = 8'h7e == total_offset_3 ? phv_data_126 : _GEN_605; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_607 = 8'h7f == total_offset_3 ? phv_data_127 : _GEN_606; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_608 = 8'h80 == total_offset_3 ? phv_data_128 : _GEN_607; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_609 = 8'h81 == total_offset_3 ? phv_data_129 : _GEN_608; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_610 = 8'h82 == total_offset_3 ? phv_data_130 : _GEN_609; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_611 = 8'h83 == total_offset_3 ? phv_data_131 : _GEN_610; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_612 = 8'h84 == total_offset_3 ? phv_data_132 : _GEN_611; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_613 = 8'h85 == total_offset_3 ? phv_data_133 : _GEN_612; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_614 = 8'h86 == total_offset_3 ? phv_data_134 : _GEN_613; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_615 = 8'h87 == total_offset_3 ? phv_data_135 : _GEN_614; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_616 = 8'h88 == total_offset_3 ? phv_data_136 : _GEN_615; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_617 = 8'h89 == total_offset_3 ? phv_data_137 : _GEN_616; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_618 = 8'h8a == total_offset_3 ? phv_data_138 : _GEN_617; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_619 = 8'h8b == total_offset_3 ? phv_data_139 : _GEN_618; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_620 = 8'h8c == total_offset_3 ? phv_data_140 : _GEN_619; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_621 = 8'h8d == total_offset_3 ? phv_data_141 : _GEN_620; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_622 = 8'h8e == total_offset_3 ? phv_data_142 : _GEN_621; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_623 = 8'h8f == total_offset_3 ? phv_data_143 : _GEN_622; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_624 = 8'h90 == total_offset_3 ? phv_data_144 : _GEN_623; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_625 = 8'h91 == total_offset_3 ? phv_data_145 : _GEN_624; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_626 = 8'h92 == total_offset_3 ? phv_data_146 : _GEN_625; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_627 = 8'h93 == total_offset_3 ? phv_data_147 : _GEN_626; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_628 = 8'h94 == total_offset_3 ? phv_data_148 : _GEN_627; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_629 = 8'h95 == total_offset_3 ? phv_data_149 : _GEN_628; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_630 = 8'h96 == total_offset_3 ? phv_data_150 : _GEN_629; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_631 = 8'h97 == total_offset_3 ? phv_data_151 : _GEN_630; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_632 = 8'h98 == total_offset_3 ? phv_data_152 : _GEN_631; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_633 = 8'h99 == total_offset_3 ? phv_data_153 : _GEN_632; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_634 = 8'h9a == total_offset_3 ? phv_data_154 : _GEN_633; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_635 = 8'h9b == total_offset_3 ? phv_data_155 : _GEN_634; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_636 = 8'h9c == total_offset_3 ? phv_data_156 : _GEN_635; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_637 = 8'h9d == total_offset_3 ? phv_data_157 : _GEN_636; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_638 = 8'h9e == total_offset_3 ? phv_data_158 : _GEN_637; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes__0 = 8'h9f == total_offset_3 ? phv_data_159 : _GEN_638; // @[executor.scala 197:66 executor.scala 197:66]
  wire [31:0] _io_field_out_0_T = {bytes__0,bytes__1,bytes__2,bytes__3}; // @[Cat.scala 30:58]
  wire [3:0] _io_mask_out_0_T = {_mask_3_T_3,mask__1,mask__2,mask__3}; // @[Cat.scala 30:58]
  wire [17:0] io_field_out_0_hi_4 = io_field_out_0_lo[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _io_field_out_0_T_4 = {io_field_out_0_hi_4,io_field_out_0_lo}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_865 = 4'hb == opcode ? _io_field_out_0_T_4 : 32'h0; // @[executor.scala 230:56 executor.scala 231:41]
  wire [1:0] _GEN_866 = from_header ? bias : 2'h0; // @[executor.scala 178:36 executor.scala 203:36 executor.scala 174:29]
  wire [31:0] _GEN_867 = from_header ? _io_field_out_0_T : _GEN_865; // @[executor.scala 178:36 executor.scala 204:37]
  wire [3:0] _GEN_868 = from_header ? _io_mask_out_0_T : 4'h0; // @[executor.scala 178:36 executor.scala 205:37 executor.scala 173:29]
  wire [3:0] opcode_1 = vliw_1[31:28]; // @[primitive.scala 9:44]
  wire [13:0] io_field_out_1_lo = vliw_1[13:0]; // @[primitive.scala 11:44]
  wire  from_header_1 = length_1 != 8'h0; // @[executor.scala 177:45]
  wire [5:0] total_offset_hi_1 = offset_1[7:2]; // @[executor.scala 191:57]
  wire [7:0] _ending_T_3 = offset_1 + length_1; // @[executor.scala 193:46]
  wire [1:0] ending_1 = _ending_T_3[1:0]; // @[executor.scala 193:58]
  wire [3:0] _GEN_3495 = {{2'd0}, ending_1}; // @[executor.scala 194:45]
  wire [3:0] _bias_T_3 = 4'h4 - _GEN_3495; // @[executor.scala 194:45]
  wire [1:0] bias_1 = _bias_T_3[1:0]; // @[executor.scala 194:54]
  wire [7:0] total_offset_4 = {total_offset_hi_1,2'h0}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_873 = 8'h1 == total_offset_4 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_874 = 8'h2 == total_offset_4 ? phv_data_2 : _GEN_873; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_875 = 8'h3 == total_offset_4 ? phv_data_3 : _GEN_874; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_876 = 8'h4 == total_offset_4 ? phv_data_4 : _GEN_875; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_877 = 8'h5 == total_offset_4 ? phv_data_5 : _GEN_876; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_878 = 8'h6 == total_offset_4 ? phv_data_6 : _GEN_877; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_879 = 8'h7 == total_offset_4 ? phv_data_7 : _GEN_878; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_880 = 8'h8 == total_offset_4 ? phv_data_8 : _GEN_879; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_881 = 8'h9 == total_offset_4 ? phv_data_9 : _GEN_880; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_882 = 8'ha == total_offset_4 ? phv_data_10 : _GEN_881; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_883 = 8'hb == total_offset_4 ? phv_data_11 : _GEN_882; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_884 = 8'hc == total_offset_4 ? phv_data_12 : _GEN_883; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_885 = 8'hd == total_offset_4 ? phv_data_13 : _GEN_884; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_886 = 8'he == total_offset_4 ? phv_data_14 : _GEN_885; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_887 = 8'hf == total_offset_4 ? phv_data_15 : _GEN_886; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_888 = 8'h10 == total_offset_4 ? phv_data_16 : _GEN_887; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_889 = 8'h11 == total_offset_4 ? phv_data_17 : _GEN_888; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_890 = 8'h12 == total_offset_4 ? phv_data_18 : _GEN_889; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_891 = 8'h13 == total_offset_4 ? phv_data_19 : _GEN_890; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_892 = 8'h14 == total_offset_4 ? phv_data_20 : _GEN_891; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_893 = 8'h15 == total_offset_4 ? phv_data_21 : _GEN_892; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_894 = 8'h16 == total_offset_4 ? phv_data_22 : _GEN_893; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_895 = 8'h17 == total_offset_4 ? phv_data_23 : _GEN_894; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_896 = 8'h18 == total_offset_4 ? phv_data_24 : _GEN_895; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_897 = 8'h19 == total_offset_4 ? phv_data_25 : _GEN_896; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_898 = 8'h1a == total_offset_4 ? phv_data_26 : _GEN_897; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_899 = 8'h1b == total_offset_4 ? phv_data_27 : _GEN_898; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_900 = 8'h1c == total_offset_4 ? phv_data_28 : _GEN_899; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_901 = 8'h1d == total_offset_4 ? phv_data_29 : _GEN_900; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_902 = 8'h1e == total_offset_4 ? phv_data_30 : _GEN_901; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_903 = 8'h1f == total_offset_4 ? phv_data_31 : _GEN_902; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_904 = 8'h20 == total_offset_4 ? phv_data_32 : _GEN_903; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_905 = 8'h21 == total_offset_4 ? phv_data_33 : _GEN_904; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_906 = 8'h22 == total_offset_4 ? phv_data_34 : _GEN_905; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_907 = 8'h23 == total_offset_4 ? phv_data_35 : _GEN_906; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_908 = 8'h24 == total_offset_4 ? phv_data_36 : _GEN_907; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_909 = 8'h25 == total_offset_4 ? phv_data_37 : _GEN_908; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_910 = 8'h26 == total_offset_4 ? phv_data_38 : _GEN_909; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_911 = 8'h27 == total_offset_4 ? phv_data_39 : _GEN_910; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_912 = 8'h28 == total_offset_4 ? phv_data_40 : _GEN_911; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_913 = 8'h29 == total_offset_4 ? phv_data_41 : _GEN_912; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_914 = 8'h2a == total_offset_4 ? phv_data_42 : _GEN_913; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_915 = 8'h2b == total_offset_4 ? phv_data_43 : _GEN_914; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_916 = 8'h2c == total_offset_4 ? phv_data_44 : _GEN_915; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_917 = 8'h2d == total_offset_4 ? phv_data_45 : _GEN_916; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_918 = 8'h2e == total_offset_4 ? phv_data_46 : _GEN_917; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_919 = 8'h2f == total_offset_4 ? phv_data_47 : _GEN_918; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_920 = 8'h30 == total_offset_4 ? phv_data_48 : _GEN_919; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_921 = 8'h31 == total_offset_4 ? phv_data_49 : _GEN_920; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_922 = 8'h32 == total_offset_4 ? phv_data_50 : _GEN_921; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_923 = 8'h33 == total_offset_4 ? phv_data_51 : _GEN_922; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_924 = 8'h34 == total_offset_4 ? phv_data_52 : _GEN_923; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_925 = 8'h35 == total_offset_4 ? phv_data_53 : _GEN_924; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_926 = 8'h36 == total_offset_4 ? phv_data_54 : _GEN_925; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_927 = 8'h37 == total_offset_4 ? phv_data_55 : _GEN_926; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_928 = 8'h38 == total_offset_4 ? phv_data_56 : _GEN_927; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_929 = 8'h39 == total_offset_4 ? phv_data_57 : _GEN_928; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_930 = 8'h3a == total_offset_4 ? phv_data_58 : _GEN_929; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_931 = 8'h3b == total_offset_4 ? phv_data_59 : _GEN_930; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_932 = 8'h3c == total_offset_4 ? phv_data_60 : _GEN_931; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_933 = 8'h3d == total_offset_4 ? phv_data_61 : _GEN_932; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_934 = 8'h3e == total_offset_4 ? phv_data_62 : _GEN_933; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_935 = 8'h3f == total_offset_4 ? phv_data_63 : _GEN_934; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_936 = 8'h40 == total_offset_4 ? phv_data_64 : _GEN_935; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_937 = 8'h41 == total_offset_4 ? phv_data_65 : _GEN_936; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_938 = 8'h42 == total_offset_4 ? phv_data_66 : _GEN_937; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_939 = 8'h43 == total_offset_4 ? phv_data_67 : _GEN_938; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_940 = 8'h44 == total_offset_4 ? phv_data_68 : _GEN_939; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_941 = 8'h45 == total_offset_4 ? phv_data_69 : _GEN_940; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_942 = 8'h46 == total_offset_4 ? phv_data_70 : _GEN_941; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_943 = 8'h47 == total_offset_4 ? phv_data_71 : _GEN_942; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_944 = 8'h48 == total_offset_4 ? phv_data_72 : _GEN_943; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_945 = 8'h49 == total_offset_4 ? phv_data_73 : _GEN_944; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_946 = 8'h4a == total_offset_4 ? phv_data_74 : _GEN_945; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_947 = 8'h4b == total_offset_4 ? phv_data_75 : _GEN_946; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_948 = 8'h4c == total_offset_4 ? phv_data_76 : _GEN_947; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_949 = 8'h4d == total_offset_4 ? phv_data_77 : _GEN_948; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_950 = 8'h4e == total_offset_4 ? phv_data_78 : _GEN_949; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_951 = 8'h4f == total_offset_4 ? phv_data_79 : _GEN_950; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_952 = 8'h50 == total_offset_4 ? phv_data_80 : _GEN_951; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_953 = 8'h51 == total_offset_4 ? phv_data_81 : _GEN_952; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_954 = 8'h52 == total_offset_4 ? phv_data_82 : _GEN_953; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_955 = 8'h53 == total_offset_4 ? phv_data_83 : _GEN_954; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_956 = 8'h54 == total_offset_4 ? phv_data_84 : _GEN_955; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_957 = 8'h55 == total_offset_4 ? phv_data_85 : _GEN_956; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_958 = 8'h56 == total_offset_4 ? phv_data_86 : _GEN_957; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_959 = 8'h57 == total_offset_4 ? phv_data_87 : _GEN_958; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_960 = 8'h58 == total_offset_4 ? phv_data_88 : _GEN_959; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_961 = 8'h59 == total_offset_4 ? phv_data_89 : _GEN_960; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_962 = 8'h5a == total_offset_4 ? phv_data_90 : _GEN_961; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_963 = 8'h5b == total_offset_4 ? phv_data_91 : _GEN_962; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_964 = 8'h5c == total_offset_4 ? phv_data_92 : _GEN_963; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_965 = 8'h5d == total_offset_4 ? phv_data_93 : _GEN_964; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_966 = 8'h5e == total_offset_4 ? phv_data_94 : _GEN_965; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_967 = 8'h5f == total_offset_4 ? phv_data_95 : _GEN_966; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_968 = 8'h60 == total_offset_4 ? phv_data_96 : _GEN_967; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_969 = 8'h61 == total_offset_4 ? phv_data_97 : _GEN_968; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_970 = 8'h62 == total_offset_4 ? phv_data_98 : _GEN_969; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_971 = 8'h63 == total_offset_4 ? phv_data_99 : _GEN_970; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_972 = 8'h64 == total_offset_4 ? phv_data_100 : _GEN_971; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_973 = 8'h65 == total_offset_4 ? phv_data_101 : _GEN_972; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_974 = 8'h66 == total_offset_4 ? phv_data_102 : _GEN_973; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_975 = 8'h67 == total_offset_4 ? phv_data_103 : _GEN_974; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_976 = 8'h68 == total_offset_4 ? phv_data_104 : _GEN_975; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_977 = 8'h69 == total_offset_4 ? phv_data_105 : _GEN_976; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_978 = 8'h6a == total_offset_4 ? phv_data_106 : _GEN_977; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_979 = 8'h6b == total_offset_4 ? phv_data_107 : _GEN_978; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_980 = 8'h6c == total_offset_4 ? phv_data_108 : _GEN_979; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_981 = 8'h6d == total_offset_4 ? phv_data_109 : _GEN_980; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_982 = 8'h6e == total_offset_4 ? phv_data_110 : _GEN_981; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_983 = 8'h6f == total_offset_4 ? phv_data_111 : _GEN_982; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_984 = 8'h70 == total_offset_4 ? phv_data_112 : _GEN_983; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_985 = 8'h71 == total_offset_4 ? phv_data_113 : _GEN_984; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_986 = 8'h72 == total_offset_4 ? phv_data_114 : _GEN_985; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_987 = 8'h73 == total_offset_4 ? phv_data_115 : _GEN_986; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_988 = 8'h74 == total_offset_4 ? phv_data_116 : _GEN_987; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_989 = 8'h75 == total_offset_4 ? phv_data_117 : _GEN_988; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_990 = 8'h76 == total_offset_4 ? phv_data_118 : _GEN_989; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_991 = 8'h77 == total_offset_4 ? phv_data_119 : _GEN_990; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_992 = 8'h78 == total_offset_4 ? phv_data_120 : _GEN_991; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_993 = 8'h79 == total_offset_4 ? phv_data_121 : _GEN_992; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_994 = 8'h7a == total_offset_4 ? phv_data_122 : _GEN_993; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_995 = 8'h7b == total_offset_4 ? phv_data_123 : _GEN_994; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_996 = 8'h7c == total_offset_4 ? phv_data_124 : _GEN_995; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_997 = 8'h7d == total_offset_4 ? phv_data_125 : _GEN_996; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_998 = 8'h7e == total_offset_4 ? phv_data_126 : _GEN_997; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_999 = 8'h7f == total_offset_4 ? phv_data_127 : _GEN_998; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1000 = 8'h80 == total_offset_4 ? phv_data_128 : _GEN_999; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1001 = 8'h81 == total_offset_4 ? phv_data_129 : _GEN_1000; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1002 = 8'h82 == total_offset_4 ? phv_data_130 : _GEN_1001; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1003 = 8'h83 == total_offset_4 ? phv_data_131 : _GEN_1002; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1004 = 8'h84 == total_offset_4 ? phv_data_132 : _GEN_1003; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1005 = 8'h85 == total_offset_4 ? phv_data_133 : _GEN_1004; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1006 = 8'h86 == total_offset_4 ? phv_data_134 : _GEN_1005; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1007 = 8'h87 == total_offset_4 ? phv_data_135 : _GEN_1006; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1008 = 8'h88 == total_offset_4 ? phv_data_136 : _GEN_1007; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1009 = 8'h89 == total_offset_4 ? phv_data_137 : _GEN_1008; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1010 = 8'h8a == total_offset_4 ? phv_data_138 : _GEN_1009; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1011 = 8'h8b == total_offset_4 ? phv_data_139 : _GEN_1010; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1012 = 8'h8c == total_offset_4 ? phv_data_140 : _GEN_1011; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1013 = 8'h8d == total_offset_4 ? phv_data_141 : _GEN_1012; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1014 = 8'h8e == total_offset_4 ? phv_data_142 : _GEN_1013; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1015 = 8'h8f == total_offset_4 ? phv_data_143 : _GEN_1014; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1016 = 8'h90 == total_offset_4 ? phv_data_144 : _GEN_1015; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1017 = 8'h91 == total_offset_4 ? phv_data_145 : _GEN_1016; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1018 = 8'h92 == total_offset_4 ? phv_data_146 : _GEN_1017; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1019 = 8'h93 == total_offset_4 ? phv_data_147 : _GEN_1018; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1020 = 8'h94 == total_offset_4 ? phv_data_148 : _GEN_1019; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1021 = 8'h95 == total_offset_4 ? phv_data_149 : _GEN_1020; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1022 = 8'h96 == total_offset_4 ? phv_data_150 : _GEN_1021; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1023 = 8'h97 == total_offset_4 ? phv_data_151 : _GEN_1022; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1024 = 8'h98 == total_offset_4 ? phv_data_152 : _GEN_1023; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1025 = 8'h99 == total_offset_4 ? phv_data_153 : _GEN_1024; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1026 = 8'h9a == total_offset_4 ? phv_data_154 : _GEN_1025; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1027 = 8'h9b == total_offset_4 ? phv_data_155 : _GEN_1026; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1028 = 8'h9c == total_offset_4 ? phv_data_156 : _GEN_1027; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1029 = 8'h9d == total_offset_4 ? phv_data_157 : _GEN_1028; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1030 = 8'h9e == total_offset_4 ? phv_data_158 : _GEN_1029; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes_1_3 = 8'h9f == total_offset_4 ? phv_data_159 : _GEN_1030; // @[executor.scala 197:66 executor.scala 197:66]
  wire  _mask_3_T_10 = ending_1 == 2'h0; // @[executor.scala 199:88]
  wire  mask_1_3 = 2'h0 >= offset_1[1:0] & (2'h0 < ending_1 | ending_1 == 2'h0); // @[executor.scala 199:56]
  wire [7:0] total_offset_5 = {total_offset_hi_1,2'h1}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_1033 = 8'h1 == total_offset_5 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1034 = 8'h2 == total_offset_5 ? phv_data_2 : _GEN_1033; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1035 = 8'h3 == total_offset_5 ? phv_data_3 : _GEN_1034; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1036 = 8'h4 == total_offset_5 ? phv_data_4 : _GEN_1035; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1037 = 8'h5 == total_offset_5 ? phv_data_5 : _GEN_1036; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1038 = 8'h6 == total_offset_5 ? phv_data_6 : _GEN_1037; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1039 = 8'h7 == total_offset_5 ? phv_data_7 : _GEN_1038; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1040 = 8'h8 == total_offset_5 ? phv_data_8 : _GEN_1039; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1041 = 8'h9 == total_offset_5 ? phv_data_9 : _GEN_1040; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1042 = 8'ha == total_offset_5 ? phv_data_10 : _GEN_1041; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1043 = 8'hb == total_offset_5 ? phv_data_11 : _GEN_1042; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1044 = 8'hc == total_offset_5 ? phv_data_12 : _GEN_1043; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1045 = 8'hd == total_offset_5 ? phv_data_13 : _GEN_1044; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1046 = 8'he == total_offset_5 ? phv_data_14 : _GEN_1045; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1047 = 8'hf == total_offset_5 ? phv_data_15 : _GEN_1046; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1048 = 8'h10 == total_offset_5 ? phv_data_16 : _GEN_1047; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1049 = 8'h11 == total_offset_5 ? phv_data_17 : _GEN_1048; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1050 = 8'h12 == total_offset_5 ? phv_data_18 : _GEN_1049; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1051 = 8'h13 == total_offset_5 ? phv_data_19 : _GEN_1050; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1052 = 8'h14 == total_offset_5 ? phv_data_20 : _GEN_1051; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1053 = 8'h15 == total_offset_5 ? phv_data_21 : _GEN_1052; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1054 = 8'h16 == total_offset_5 ? phv_data_22 : _GEN_1053; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1055 = 8'h17 == total_offset_5 ? phv_data_23 : _GEN_1054; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1056 = 8'h18 == total_offset_5 ? phv_data_24 : _GEN_1055; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1057 = 8'h19 == total_offset_5 ? phv_data_25 : _GEN_1056; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1058 = 8'h1a == total_offset_5 ? phv_data_26 : _GEN_1057; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1059 = 8'h1b == total_offset_5 ? phv_data_27 : _GEN_1058; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1060 = 8'h1c == total_offset_5 ? phv_data_28 : _GEN_1059; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1061 = 8'h1d == total_offset_5 ? phv_data_29 : _GEN_1060; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1062 = 8'h1e == total_offset_5 ? phv_data_30 : _GEN_1061; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1063 = 8'h1f == total_offset_5 ? phv_data_31 : _GEN_1062; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1064 = 8'h20 == total_offset_5 ? phv_data_32 : _GEN_1063; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1065 = 8'h21 == total_offset_5 ? phv_data_33 : _GEN_1064; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1066 = 8'h22 == total_offset_5 ? phv_data_34 : _GEN_1065; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1067 = 8'h23 == total_offset_5 ? phv_data_35 : _GEN_1066; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1068 = 8'h24 == total_offset_5 ? phv_data_36 : _GEN_1067; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1069 = 8'h25 == total_offset_5 ? phv_data_37 : _GEN_1068; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1070 = 8'h26 == total_offset_5 ? phv_data_38 : _GEN_1069; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1071 = 8'h27 == total_offset_5 ? phv_data_39 : _GEN_1070; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1072 = 8'h28 == total_offset_5 ? phv_data_40 : _GEN_1071; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1073 = 8'h29 == total_offset_5 ? phv_data_41 : _GEN_1072; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1074 = 8'h2a == total_offset_5 ? phv_data_42 : _GEN_1073; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1075 = 8'h2b == total_offset_5 ? phv_data_43 : _GEN_1074; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1076 = 8'h2c == total_offset_5 ? phv_data_44 : _GEN_1075; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1077 = 8'h2d == total_offset_5 ? phv_data_45 : _GEN_1076; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1078 = 8'h2e == total_offset_5 ? phv_data_46 : _GEN_1077; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1079 = 8'h2f == total_offset_5 ? phv_data_47 : _GEN_1078; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1080 = 8'h30 == total_offset_5 ? phv_data_48 : _GEN_1079; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1081 = 8'h31 == total_offset_5 ? phv_data_49 : _GEN_1080; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1082 = 8'h32 == total_offset_5 ? phv_data_50 : _GEN_1081; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1083 = 8'h33 == total_offset_5 ? phv_data_51 : _GEN_1082; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1084 = 8'h34 == total_offset_5 ? phv_data_52 : _GEN_1083; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1085 = 8'h35 == total_offset_5 ? phv_data_53 : _GEN_1084; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1086 = 8'h36 == total_offset_5 ? phv_data_54 : _GEN_1085; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1087 = 8'h37 == total_offset_5 ? phv_data_55 : _GEN_1086; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1088 = 8'h38 == total_offset_5 ? phv_data_56 : _GEN_1087; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1089 = 8'h39 == total_offset_5 ? phv_data_57 : _GEN_1088; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1090 = 8'h3a == total_offset_5 ? phv_data_58 : _GEN_1089; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1091 = 8'h3b == total_offset_5 ? phv_data_59 : _GEN_1090; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1092 = 8'h3c == total_offset_5 ? phv_data_60 : _GEN_1091; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1093 = 8'h3d == total_offset_5 ? phv_data_61 : _GEN_1092; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1094 = 8'h3e == total_offset_5 ? phv_data_62 : _GEN_1093; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1095 = 8'h3f == total_offset_5 ? phv_data_63 : _GEN_1094; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1096 = 8'h40 == total_offset_5 ? phv_data_64 : _GEN_1095; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1097 = 8'h41 == total_offset_5 ? phv_data_65 : _GEN_1096; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1098 = 8'h42 == total_offset_5 ? phv_data_66 : _GEN_1097; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1099 = 8'h43 == total_offset_5 ? phv_data_67 : _GEN_1098; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1100 = 8'h44 == total_offset_5 ? phv_data_68 : _GEN_1099; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1101 = 8'h45 == total_offset_5 ? phv_data_69 : _GEN_1100; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1102 = 8'h46 == total_offset_5 ? phv_data_70 : _GEN_1101; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1103 = 8'h47 == total_offset_5 ? phv_data_71 : _GEN_1102; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1104 = 8'h48 == total_offset_5 ? phv_data_72 : _GEN_1103; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1105 = 8'h49 == total_offset_5 ? phv_data_73 : _GEN_1104; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1106 = 8'h4a == total_offset_5 ? phv_data_74 : _GEN_1105; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1107 = 8'h4b == total_offset_5 ? phv_data_75 : _GEN_1106; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1108 = 8'h4c == total_offset_5 ? phv_data_76 : _GEN_1107; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1109 = 8'h4d == total_offset_5 ? phv_data_77 : _GEN_1108; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1110 = 8'h4e == total_offset_5 ? phv_data_78 : _GEN_1109; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1111 = 8'h4f == total_offset_5 ? phv_data_79 : _GEN_1110; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1112 = 8'h50 == total_offset_5 ? phv_data_80 : _GEN_1111; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1113 = 8'h51 == total_offset_5 ? phv_data_81 : _GEN_1112; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1114 = 8'h52 == total_offset_5 ? phv_data_82 : _GEN_1113; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1115 = 8'h53 == total_offset_5 ? phv_data_83 : _GEN_1114; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1116 = 8'h54 == total_offset_5 ? phv_data_84 : _GEN_1115; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1117 = 8'h55 == total_offset_5 ? phv_data_85 : _GEN_1116; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1118 = 8'h56 == total_offset_5 ? phv_data_86 : _GEN_1117; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1119 = 8'h57 == total_offset_5 ? phv_data_87 : _GEN_1118; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1120 = 8'h58 == total_offset_5 ? phv_data_88 : _GEN_1119; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1121 = 8'h59 == total_offset_5 ? phv_data_89 : _GEN_1120; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1122 = 8'h5a == total_offset_5 ? phv_data_90 : _GEN_1121; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1123 = 8'h5b == total_offset_5 ? phv_data_91 : _GEN_1122; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1124 = 8'h5c == total_offset_5 ? phv_data_92 : _GEN_1123; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1125 = 8'h5d == total_offset_5 ? phv_data_93 : _GEN_1124; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1126 = 8'h5e == total_offset_5 ? phv_data_94 : _GEN_1125; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1127 = 8'h5f == total_offset_5 ? phv_data_95 : _GEN_1126; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1128 = 8'h60 == total_offset_5 ? phv_data_96 : _GEN_1127; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1129 = 8'h61 == total_offset_5 ? phv_data_97 : _GEN_1128; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1130 = 8'h62 == total_offset_5 ? phv_data_98 : _GEN_1129; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1131 = 8'h63 == total_offset_5 ? phv_data_99 : _GEN_1130; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1132 = 8'h64 == total_offset_5 ? phv_data_100 : _GEN_1131; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1133 = 8'h65 == total_offset_5 ? phv_data_101 : _GEN_1132; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1134 = 8'h66 == total_offset_5 ? phv_data_102 : _GEN_1133; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1135 = 8'h67 == total_offset_5 ? phv_data_103 : _GEN_1134; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1136 = 8'h68 == total_offset_5 ? phv_data_104 : _GEN_1135; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1137 = 8'h69 == total_offset_5 ? phv_data_105 : _GEN_1136; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1138 = 8'h6a == total_offset_5 ? phv_data_106 : _GEN_1137; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1139 = 8'h6b == total_offset_5 ? phv_data_107 : _GEN_1138; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1140 = 8'h6c == total_offset_5 ? phv_data_108 : _GEN_1139; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1141 = 8'h6d == total_offset_5 ? phv_data_109 : _GEN_1140; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1142 = 8'h6e == total_offset_5 ? phv_data_110 : _GEN_1141; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1143 = 8'h6f == total_offset_5 ? phv_data_111 : _GEN_1142; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1144 = 8'h70 == total_offset_5 ? phv_data_112 : _GEN_1143; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1145 = 8'h71 == total_offset_5 ? phv_data_113 : _GEN_1144; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1146 = 8'h72 == total_offset_5 ? phv_data_114 : _GEN_1145; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1147 = 8'h73 == total_offset_5 ? phv_data_115 : _GEN_1146; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1148 = 8'h74 == total_offset_5 ? phv_data_116 : _GEN_1147; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1149 = 8'h75 == total_offset_5 ? phv_data_117 : _GEN_1148; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1150 = 8'h76 == total_offset_5 ? phv_data_118 : _GEN_1149; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1151 = 8'h77 == total_offset_5 ? phv_data_119 : _GEN_1150; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1152 = 8'h78 == total_offset_5 ? phv_data_120 : _GEN_1151; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1153 = 8'h79 == total_offset_5 ? phv_data_121 : _GEN_1152; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1154 = 8'h7a == total_offset_5 ? phv_data_122 : _GEN_1153; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1155 = 8'h7b == total_offset_5 ? phv_data_123 : _GEN_1154; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1156 = 8'h7c == total_offset_5 ? phv_data_124 : _GEN_1155; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1157 = 8'h7d == total_offset_5 ? phv_data_125 : _GEN_1156; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1158 = 8'h7e == total_offset_5 ? phv_data_126 : _GEN_1157; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1159 = 8'h7f == total_offset_5 ? phv_data_127 : _GEN_1158; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1160 = 8'h80 == total_offset_5 ? phv_data_128 : _GEN_1159; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1161 = 8'h81 == total_offset_5 ? phv_data_129 : _GEN_1160; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1162 = 8'h82 == total_offset_5 ? phv_data_130 : _GEN_1161; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1163 = 8'h83 == total_offset_5 ? phv_data_131 : _GEN_1162; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1164 = 8'h84 == total_offset_5 ? phv_data_132 : _GEN_1163; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1165 = 8'h85 == total_offset_5 ? phv_data_133 : _GEN_1164; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1166 = 8'h86 == total_offset_5 ? phv_data_134 : _GEN_1165; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1167 = 8'h87 == total_offset_5 ? phv_data_135 : _GEN_1166; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1168 = 8'h88 == total_offset_5 ? phv_data_136 : _GEN_1167; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1169 = 8'h89 == total_offset_5 ? phv_data_137 : _GEN_1168; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1170 = 8'h8a == total_offset_5 ? phv_data_138 : _GEN_1169; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1171 = 8'h8b == total_offset_5 ? phv_data_139 : _GEN_1170; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1172 = 8'h8c == total_offset_5 ? phv_data_140 : _GEN_1171; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1173 = 8'h8d == total_offset_5 ? phv_data_141 : _GEN_1172; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1174 = 8'h8e == total_offset_5 ? phv_data_142 : _GEN_1173; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1175 = 8'h8f == total_offset_5 ? phv_data_143 : _GEN_1174; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1176 = 8'h90 == total_offset_5 ? phv_data_144 : _GEN_1175; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1177 = 8'h91 == total_offset_5 ? phv_data_145 : _GEN_1176; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1178 = 8'h92 == total_offset_5 ? phv_data_146 : _GEN_1177; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1179 = 8'h93 == total_offset_5 ? phv_data_147 : _GEN_1178; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1180 = 8'h94 == total_offset_5 ? phv_data_148 : _GEN_1179; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1181 = 8'h95 == total_offset_5 ? phv_data_149 : _GEN_1180; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1182 = 8'h96 == total_offset_5 ? phv_data_150 : _GEN_1181; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1183 = 8'h97 == total_offset_5 ? phv_data_151 : _GEN_1182; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1184 = 8'h98 == total_offset_5 ? phv_data_152 : _GEN_1183; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1185 = 8'h99 == total_offset_5 ? phv_data_153 : _GEN_1184; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1186 = 8'h9a == total_offset_5 ? phv_data_154 : _GEN_1185; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1187 = 8'h9b == total_offset_5 ? phv_data_155 : _GEN_1186; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1188 = 8'h9c == total_offset_5 ? phv_data_156 : _GEN_1187; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1189 = 8'h9d == total_offset_5 ? phv_data_157 : _GEN_1188; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1190 = 8'h9e == total_offset_5 ? phv_data_158 : _GEN_1189; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes_1_2 = 8'h9f == total_offset_5 ? phv_data_159 : _GEN_1190; // @[executor.scala 197:66 executor.scala 197:66]
  wire  mask_1_2 = 2'h1 >= offset_1[1:0] & (2'h1 < ending_1 | ending_1 == 2'h0); // @[executor.scala 199:56]
  wire [7:0] total_offset_6 = {total_offset_hi_1,2'h2}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_1193 = 8'h1 == total_offset_6 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1194 = 8'h2 == total_offset_6 ? phv_data_2 : _GEN_1193; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1195 = 8'h3 == total_offset_6 ? phv_data_3 : _GEN_1194; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1196 = 8'h4 == total_offset_6 ? phv_data_4 : _GEN_1195; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1197 = 8'h5 == total_offset_6 ? phv_data_5 : _GEN_1196; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1198 = 8'h6 == total_offset_6 ? phv_data_6 : _GEN_1197; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1199 = 8'h7 == total_offset_6 ? phv_data_7 : _GEN_1198; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1200 = 8'h8 == total_offset_6 ? phv_data_8 : _GEN_1199; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1201 = 8'h9 == total_offset_6 ? phv_data_9 : _GEN_1200; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1202 = 8'ha == total_offset_6 ? phv_data_10 : _GEN_1201; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1203 = 8'hb == total_offset_6 ? phv_data_11 : _GEN_1202; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1204 = 8'hc == total_offset_6 ? phv_data_12 : _GEN_1203; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1205 = 8'hd == total_offset_6 ? phv_data_13 : _GEN_1204; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1206 = 8'he == total_offset_6 ? phv_data_14 : _GEN_1205; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1207 = 8'hf == total_offset_6 ? phv_data_15 : _GEN_1206; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1208 = 8'h10 == total_offset_6 ? phv_data_16 : _GEN_1207; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1209 = 8'h11 == total_offset_6 ? phv_data_17 : _GEN_1208; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1210 = 8'h12 == total_offset_6 ? phv_data_18 : _GEN_1209; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1211 = 8'h13 == total_offset_6 ? phv_data_19 : _GEN_1210; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1212 = 8'h14 == total_offset_6 ? phv_data_20 : _GEN_1211; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1213 = 8'h15 == total_offset_6 ? phv_data_21 : _GEN_1212; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1214 = 8'h16 == total_offset_6 ? phv_data_22 : _GEN_1213; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1215 = 8'h17 == total_offset_6 ? phv_data_23 : _GEN_1214; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1216 = 8'h18 == total_offset_6 ? phv_data_24 : _GEN_1215; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1217 = 8'h19 == total_offset_6 ? phv_data_25 : _GEN_1216; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1218 = 8'h1a == total_offset_6 ? phv_data_26 : _GEN_1217; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1219 = 8'h1b == total_offset_6 ? phv_data_27 : _GEN_1218; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1220 = 8'h1c == total_offset_6 ? phv_data_28 : _GEN_1219; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1221 = 8'h1d == total_offset_6 ? phv_data_29 : _GEN_1220; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1222 = 8'h1e == total_offset_6 ? phv_data_30 : _GEN_1221; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1223 = 8'h1f == total_offset_6 ? phv_data_31 : _GEN_1222; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1224 = 8'h20 == total_offset_6 ? phv_data_32 : _GEN_1223; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1225 = 8'h21 == total_offset_6 ? phv_data_33 : _GEN_1224; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1226 = 8'h22 == total_offset_6 ? phv_data_34 : _GEN_1225; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1227 = 8'h23 == total_offset_6 ? phv_data_35 : _GEN_1226; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1228 = 8'h24 == total_offset_6 ? phv_data_36 : _GEN_1227; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1229 = 8'h25 == total_offset_6 ? phv_data_37 : _GEN_1228; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1230 = 8'h26 == total_offset_6 ? phv_data_38 : _GEN_1229; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1231 = 8'h27 == total_offset_6 ? phv_data_39 : _GEN_1230; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1232 = 8'h28 == total_offset_6 ? phv_data_40 : _GEN_1231; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1233 = 8'h29 == total_offset_6 ? phv_data_41 : _GEN_1232; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1234 = 8'h2a == total_offset_6 ? phv_data_42 : _GEN_1233; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1235 = 8'h2b == total_offset_6 ? phv_data_43 : _GEN_1234; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1236 = 8'h2c == total_offset_6 ? phv_data_44 : _GEN_1235; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1237 = 8'h2d == total_offset_6 ? phv_data_45 : _GEN_1236; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1238 = 8'h2e == total_offset_6 ? phv_data_46 : _GEN_1237; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1239 = 8'h2f == total_offset_6 ? phv_data_47 : _GEN_1238; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1240 = 8'h30 == total_offset_6 ? phv_data_48 : _GEN_1239; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1241 = 8'h31 == total_offset_6 ? phv_data_49 : _GEN_1240; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1242 = 8'h32 == total_offset_6 ? phv_data_50 : _GEN_1241; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1243 = 8'h33 == total_offset_6 ? phv_data_51 : _GEN_1242; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1244 = 8'h34 == total_offset_6 ? phv_data_52 : _GEN_1243; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1245 = 8'h35 == total_offset_6 ? phv_data_53 : _GEN_1244; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1246 = 8'h36 == total_offset_6 ? phv_data_54 : _GEN_1245; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1247 = 8'h37 == total_offset_6 ? phv_data_55 : _GEN_1246; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1248 = 8'h38 == total_offset_6 ? phv_data_56 : _GEN_1247; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1249 = 8'h39 == total_offset_6 ? phv_data_57 : _GEN_1248; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1250 = 8'h3a == total_offset_6 ? phv_data_58 : _GEN_1249; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1251 = 8'h3b == total_offset_6 ? phv_data_59 : _GEN_1250; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1252 = 8'h3c == total_offset_6 ? phv_data_60 : _GEN_1251; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1253 = 8'h3d == total_offset_6 ? phv_data_61 : _GEN_1252; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1254 = 8'h3e == total_offset_6 ? phv_data_62 : _GEN_1253; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1255 = 8'h3f == total_offset_6 ? phv_data_63 : _GEN_1254; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1256 = 8'h40 == total_offset_6 ? phv_data_64 : _GEN_1255; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1257 = 8'h41 == total_offset_6 ? phv_data_65 : _GEN_1256; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1258 = 8'h42 == total_offset_6 ? phv_data_66 : _GEN_1257; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1259 = 8'h43 == total_offset_6 ? phv_data_67 : _GEN_1258; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1260 = 8'h44 == total_offset_6 ? phv_data_68 : _GEN_1259; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1261 = 8'h45 == total_offset_6 ? phv_data_69 : _GEN_1260; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1262 = 8'h46 == total_offset_6 ? phv_data_70 : _GEN_1261; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1263 = 8'h47 == total_offset_6 ? phv_data_71 : _GEN_1262; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1264 = 8'h48 == total_offset_6 ? phv_data_72 : _GEN_1263; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1265 = 8'h49 == total_offset_6 ? phv_data_73 : _GEN_1264; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1266 = 8'h4a == total_offset_6 ? phv_data_74 : _GEN_1265; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1267 = 8'h4b == total_offset_6 ? phv_data_75 : _GEN_1266; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1268 = 8'h4c == total_offset_6 ? phv_data_76 : _GEN_1267; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1269 = 8'h4d == total_offset_6 ? phv_data_77 : _GEN_1268; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1270 = 8'h4e == total_offset_6 ? phv_data_78 : _GEN_1269; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1271 = 8'h4f == total_offset_6 ? phv_data_79 : _GEN_1270; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1272 = 8'h50 == total_offset_6 ? phv_data_80 : _GEN_1271; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1273 = 8'h51 == total_offset_6 ? phv_data_81 : _GEN_1272; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1274 = 8'h52 == total_offset_6 ? phv_data_82 : _GEN_1273; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1275 = 8'h53 == total_offset_6 ? phv_data_83 : _GEN_1274; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1276 = 8'h54 == total_offset_6 ? phv_data_84 : _GEN_1275; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1277 = 8'h55 == total_offset_6 ? phv_data_85 : _GEN_1276; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1278 = 8'h56 == total_offset_6 ? phv_data_86 : _GEN_1277; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1279 = 8'h57 == total_offset_6 ? phv_data_87 : _GEN_1278; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1280 = 8'h58 == total_offset_6 ? phv_data_88 : _GEN_1279; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1281 = 8'h59 == total_offset_6 ? phv_data_89 : _GEN_1280; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1282 = 8'h5a == total_offset_6 ? phv_data_90 : _GEN_1281; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1283 = 8'h5b == total_offset_6 ? phv_data_91 : _GEN_1282; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1284 = 8'h5c == total_offset_6 ? phv_data_92 : _GEN_1283; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1285 = 8'h5d == total_offset_6 ? phv_data_93 : _GEN_1284; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1286 = 8'h5e == total_offset_6 ? phv_data_94 : _GEN_1285; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1287 = 8'h5f == total_offset_6 ? phv_data_95 : _GEN_1286; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1288 = 8'h60 == total_offset_6 ? phv_data_96 : _GEN_1287; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1289 = 8'h61 == total_offset_6 ? phv_data_97 : _GEN_1288; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1290 = 8'h62 == total_offset_6 ? phv_data_98 : _GEN_1289; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1291 = 8'h63 == total_offset_6 ? phv_data_99 : _GEN_1290; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1292 = 8'h64 == total_offset_6 ? phv_data_100 : _GEN_1291; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1293 = 8'h65 == total_offset_6 ? phv_data_101 : _GEN_1292; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1294 = 8'h66 == total_offset_6 ? phv_data_102 : _GEN_1293; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1295 = 8'h67 == total_offset_6 ? phv_data_103 : _GEN_1294; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1296 = 8'h68 == total_offset_6 ? phv_data_104 : _GEN_1295; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1297 = 8'h69 == total_offset_6 ? phv_data_105 : _GEN_1296; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1298 = 8'h6a == total_offset_6 ? phv_data_106 : _GEN_1297; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1299 = 8'h6b == total_offset_6 ? phv_data_107 : _GEN_1298; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1300 = 8'h6c == total_offset_6 ? phv_data_108 : _GEN_1299; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1301 = 8'h6d == total_offset_6 ? phv_data_109 : _GEN_1300; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1302 = 8'h6e == total_offset_6 ? phv_data_110 : _GEN_1301; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1303 = 8'h6f == total_offset_6 ? phv_data_111 : _GEN_1302; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1304 = 8'h70 == total_offset_6 ? phv_data_112 : _GEN_1303; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1305 = 8'h71 == total_offset_6 ? phv_data_113 : _GEN_1304; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1306 = 8'h72 == total_offset_6 ? phv_data_114 : _GEN_1305; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1307 = 8'h73 == total_offset_6 ? phv_data_115 : _GEN_1306; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1308 = 8'h74 == total_offset_6 ? phv_data_116 : _GEN_1307; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1309 = 8'h75 == total_offset_6 ? phv_data_117 : _GEN_1308; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1310 = 8'h76 == total_offset_6 ? phv_data_118 : _GEN_1309; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1311 = 8'h77 == total_offset_6 ? phv_data_119 : _GEN_1310; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1312 = 8'h78 == total_offset_6 ? phv_data_120 : _GEN_1311; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1313 = 8'h79 == total_offset_6 ? phv_data_121 : _GEN_1312; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1314 = 8'h7a == total_offset_6 ? phv_data_122 : _GEN_1313; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1315 = 8'h7b == total_offset_6 ? phv_data_123 : _GEN_1314; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1316 = 8'h7c == total_offset_6 ? phv_data_124 : _GEN_1315; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1317 = 8'h7d == total_offset_6 ? phv_data_125 : _GEN_1316; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1318 = 8'h7e == total_offset_6 ? phv_data_126 : _GEN_1317; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1319 = 8'h7f == total_offset_6 ? phv_data_127 : _GEN_1318; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1320 = 8'h80 == total_offset_6 ? phv_data_128 : _GEN_1319; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1321 = 8'h81 == total_offset_6 ? phv_data_129 : _GEN_1320; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1322 = 8'h82 == total_offset_6 ? phv_data_130 : _GEN_1321; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1323 = 8'h83 == total_offset_6 ? phv_data_131 : _GEN_1322; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1324 = 8'h84 == total_offset_6 ? phv_data_132 : _GEN_1323; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1325 = 8'h85 == total_offset_6 ? phv_data_133 : _GEN_1324; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1326 = 8'h86 == total_offset_6 ? phv_data_134 : _GEN_1325; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1327 = 8'h87 == total_offset_6 ? phv_data_135 : _GEN_1326; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1328 = 8'h88 == total_offset_6 ? phv_data_136 : _GEN_1327; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1329 = 8'h89 == total_offset_6 ? phv_data_137 : _GEN_1328; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1330 = 8'h8a == total_offset_6 ? phv_data_138 : _GEN_1329; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1331 = 8'h8b == total_offset_6 ? phv_data_139 : _GEN_1330; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1332 = 8'h8c == total_offset_6 ? phv_data_140 : _GEN_1331; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1333 = 8'h8d == total_offset_6 ? phv_data_141 : _GEN_1332; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1334 = 8'h8e == total_offset_6 ? phv_data_142 : _GEN_1333; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1335 = 8'h8f == total_offset_6 ? phv_data_143 : _GEN_1334; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1336 = 8'h90 == total_offset_6 ? phv_data_144 : _GEN_1335; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1337 = 8'h91 == total_offset_6 ? phv_data_145 : _GEN_1336; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1338 = 8'h92 == total_offset_6 ? phv_data_146 : _GEN_1337; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1339 = 8'h93 == total_offset_6 ? phv_data_147 : _GEN_1338; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1340 = 8'h94 == total_offset_6 ? phv_data_148 : _GEN_1339; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1341 = 8'h95 == total_offset_6 ? phv_data_149 : _GEN_1340; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1342 = 8'h96 == total_offset_6 ? phv_data_150 : _GEN_1341; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1343 = 8'h97 == total_offset_6 ? phv_data_151 : _GEN_1342; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1344 = 8'h98 == total_offset_6 ? phv_data_152 : _GEN_1343; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1345 = 8'h99 == total_offset_6 ? phv_data_153 : _GEN_1344; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1346 = 8'h9a == total_offset_6 ? phv_data_154 : _GEN_1345; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1347 = 8'h9b == total_offset_6 ? phv_data_155 : _GEN_1346; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1348 = 8'h9c == total_offset_6 ? phv_data_156 : _GEN_1347; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1349 = 8'h9d == total_offset_6 ? phv_data_157 : _GEN_1348; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1350 = 8'h9e == total_offset_6 ? phv_data_158 : _GEN_1349; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes_1_1 = 8'h9f == total_offset_6 ? phv_data_159 : _GEN_1350; // @[executor.scala 197:66 executor.scala 197:66]
  wire  mask_1_1 = 2'h2 >= offset_1[1:0] & (2'h2 < ending_1 | ending_1 == 2'h0); // @[executor.scala 199:56]
  wire [7:0] total_offset_7 = {total_offset_hi_1,2'h3}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_1353 = 8'h1 == total_offset_7 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1354 = 8'h2 == total_offset_7 ? phv_data_2 : _GEN_1353; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1355 = 8'h3 == total_offset_7 ? phv_data_3 : _GEN_1354; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1356 = 8'h4 == total_offset_7 ? phv_data_4 : _GEN_1355; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1357 = 8'h5 == total_offset_7 ? phv_data_5 : _GEN_1356; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1358 = 8'h6 == total_offset_7 ? phv_data_6 : _GEN_1357; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1359 = 8'h7 == total_offset_7 ? phv_data_7 : _GEN_1358; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1360 = 8'h8 == total_offset_7 ? phv_data_8 : _GEN_1359; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1361 = 8'h9 == total_offset_7 ? phv_data_9 : _GEN_1360; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1362 = 8'ha == total_offset_7 ? phv_data_10 : _GEN_1361; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1363 = 8'hb == total_offset_7 ? phv_data_11 : _GEN_1362; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1364 = 8'hc == total_offset_7 ? phv_data_12 : _GEN_1363; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1365 = 8'hd == total_offset_7 ? phv_data_13 : _GEN_1364; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1366 = 8'he == total_offset_7 ? phv_data_14 : _GEN_1365; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1367 = 8'hf == total_offset_7 ? phv_data_15 : _GEN_1366; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1368 = 8'h10 == total_offset_7 ? phv_data_16 : _GEN_1367; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1369 = 8'h11 == total_offset_7 ? phv_data_17 : _GEN_1368; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1370 = 8'h12 == total_offset_7 ? phv_data_18 : _GEN_1369; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1371 = 8'h13 == total_offset_7 ? phv_data_19 : _GEN_1370; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1372 = 8'h14 == total_offset_7 ? phv_data_20 : _GEN_1371; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1373 = 8'h15 == total_offset_7 ? phv_data_21 : _GEN_1372; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1374 = 8'h16 == total_offset_7 ? phv_data_22 : _GEN_1373; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1375 = 8'h17 == total_offset_7 ? phv_data_23 : _GEN_1374; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1376 = 8'h18 == total_offset_7 ? phv_data_24 : _GEN_1375; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1377 = 8'h19 == total_offset_7 ? phv_data_25 : _GEN_1376; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1378 = 8'h1a == total_offset_7 ? phv_data_26 : _GEN_1377; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1379 = 8'h1b == total_offset_7 ? phv_data_27 : _GEN_1378; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1380 = 8'h1c == total_offset_7 ? phv_data_28 : _GEN_1379; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1381 = 8'h1d == total_offset_7 ? phv_data_29 : _GEN_1380; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1382 = 8'h1e == total_offset_7 ? phv_data_30 : _GEN_1381; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1383 = 8'h1f == total_offset_7 ? phv_data_31 : _GEN_1382; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1384 = 8'h20 == total_offset_7 ? phv_data_32 : _GEN_1383; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1385 = 8'h21 == total_offset_7 ? phv_data_33 : _GEN_1384; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1386 = 8'h22 == total_offset_7 ? phv_data_34 : _GEN_1385; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1387 = 8'h23 == total_offset_7 ? phv_data_35 : _GEN_1386; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1388 = 8'h24 == total_offset_7 ? phv_data_36 : _GEN_1387; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1389 = 8'h25 == total_offset_7 ? phv_data_37 : _GEN_1388; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1390 = 8'h26 == total_offset_7 ? phv_data_38 : _GEN_1389; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1391 = 8'h27 == total_offset_7 ? phv_data_39 : _GEN_1390; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1392 = 8'h28 == total_offset_7 ? phv_data_40 : _GEN_1391; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1393 = 8'h29 == total_offset_7 ? phv_data_41 : _GEN_1392; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1394 = 8'h2a == total_offset_7 ? phv_data_42 : _GEN_1393; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1395 = 8'h2b == total_offset_7 ? phv_data_43 : _GEN_1394; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1396 = 8'h2c == total_offset_7 ? phv_data_44 : _GEN_1395; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1397 = 8'h2d == total_offset_7 ? phv_data_45 : _GEN_1396; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1398 = 8'h2e == total_offset_7 ? phv_data_46 : _GEN_1397; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1399 = 8'h2f == total_offset_7 ? phv_data_47 : _GEN_1398; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1400 = 8'h30 == total_offset_7 ? phv_data_48 : _GEN_1399; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1401 = 8'h31 == total_offset_7 ? phv_data_49 : _GEN_1400; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1402 = 8'h32 == total_offset_7 ? phv_data_50 : _GEN_1401; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1403 = 8'h33 == total_offset_7 ? phv_data_51 : _GEN_1402; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1404 = 8'h34 == total_offset_7 ? phv_data_52 : _GEN_1403; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1405 = 8'h35 == total_offset_7 ? phv_data_53 : _GEN_1404; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1406 = 8'h36 == total_offset_7 ? phv_data_54 : _GEN_1405; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1407 = 8'h37 == total_offset_7 ? phv_data_55 : _GEN_1406; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1408 = 8'h38 == total_offset_7 ? phv_data_56 : _GEN_1407; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1409 = 8'h39 == total_offset_7 ? phv_data_57 : _GEN_1408; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1410 = 8'h3a == total_offset_7 ? phv_data_58 : _GEN_1409; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1411 = 8'h3b == total_offset_7 ? phv_data_59 : _GEN_1410; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1412 = 8'h3c == total_offset_7 ? phv_data_60 : _GEN_1411; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1413 = 8'h3d == total_offset_7 ? phv_data_61 : _GEN_1412; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1414 = 8'h3e == total_offset_7 ? phv_data_62 : _GEN_1413; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1415 = 8'h3f == total_offset_7 ? phv_data_63 : _GEN_1414; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1416 = 8'h40 == total_offset_7 ? phv_data_64 : _GEN_1415; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1417 = 8'h41 == total_offset_7 ? phv_data_65 : _GEN_1416; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1418 = 8'h42 == total_offset_7 ? phv_data_66 : _GEN_1417; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1419 = 8'h43 == total_offset_7 ? phv_data_67 : _GEN_1418; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1420 = 8'h44 == total_offset_7 ? phv_data_68 : _GEN_1419; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1421 = 8'h45 == total_offset_7 ? phv_data_69 : _GEN_1420; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1422 = 8'h46 == total_offset_7 ? phv_data_70 : _GEN_1421; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1423 = 8'h47 == total_offset_7 ? phv_data_71 : _GEN_1422; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1424 = 8'h48 == total_offset_7 ? phv_data_72 : _GEN_1423; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1425 = 8'h49 == total_offset_7 ? phv_data_73 : _GEN_1424; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1426 = 8'h4a == total_offset_7 ? phv_data_74 : _GEN_1425; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1427 = 8'h4b == total_offset_7 ? phv_data_75 : _GEN_1426; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1428 = 8'h4c == total_offset_7 ? phv_data_76 : _GEN_1427; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1429 = 8'h4d == total_offset_7 ? phv_data_77 : _GEN_1428; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1430 = 8'h4e == total_offset_7 ? phv_data_78 : _GEN_1429; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1431 = 8'h4f == total_offset_7 ? phv_data_79 : _GEN_1430; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1432 = 8'h50 == total_offset_7 ? phv_data_80 : _GEN_1431; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1433 = 8'h51 == total_offset_7 ? phv_data_81 : _GEN_1432; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1434 = 8'h52 == total_offset_7 ? phv_data_82 : _GEN_1433; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1435 = 8'h53 == total_offset_7 ? phv_data_83 : _GEN_1434; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1436 = 8'h54 == total_offset_7 ? phv_data_84 : _GEN_1435; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1437 = 8'h55 == total_offset_7 ? phv_data_85 : _GEN_1436; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1438 = 8'h56 == total_offset_7 ? phv_data_86 : _GEN_1437; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1439 = 8'h57 == total_offset_7 ? phv_data_87 : _GEN_1438; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1440 = 8'h58 == total_offset_7 ? phv_data_88 : _GEN_1439; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1441 = 8'h59 == total_offset_7 ? phv_data_89 : _GEN_1440; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1442 = 8'h5a == total_offset_7 ? phv_data_90 : _GEN_1441; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1443 = 8'h5b == total_offset_7 ? phv_data_91 : _GEN_1442; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1444 = 8'h5c == total_offset_7 ? phv_data_92 : _GEN_1443; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1445 = 8'h5d == total_offset_7 ? phv_data_93 : _GEN_1444; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1446 = 8'h5e == total_offset_7 ? phv_data_94 : _GEN_1445; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1447 = 8'h5f == total_offset_7 ? phv_data_95 : _GEN_1446; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1448 = 8'h60 == total_offset_7 ? phv_data_96 : _GEN_1447; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1449 = 8'h61 == total_offset_7 ? phv_data_97 : _GEN_1448; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1450 = 8'h62 == total_offset_7 ? phv_data_98 : _GEN_1449; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1451 = 8'h63 == total_offset_7 ? phv_data_99 : _GEN_1450; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1452 = 8'h64 == total_offset_7 ? phv_data_100 : _GEN_1451; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1453 = 8'h65 == total_offset_7 ? phv_data_101 : _GEN_1452; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1454 = 8'h66 == total_offset_7 ? phv_data_102 : _GEN_1453; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1455 = 8'h67 == total_offset_7 ? phv_data_103 : _GEN_1454; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1456 = 8'h68 == total_offset_7 ? phv_data_104 : _GEN_1455; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1457 = 8'h69 == total_offset_7 ? phv_data_105 : _GEN_1456; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1458 = 8'h6a == total_offset_7 ? phv_data_106 : _GEN_1457; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1459 = 8'h6b == total_offset_7 ? phv_data_107 : _GEN_1458; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1460 = 8'h6c == total_offset_7 ? phv_data_108 : _GEN_1459; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1461 = 8'h6d == total_offset_7 ? phv_data_109 : _GEN_1460; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1462 = 8'h6e == total_offset_7 ? phv_data_110 : _GEN_1461; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1463 = 8'h6f == total_offset_7 ? phv_data_111 : _GEN_1462; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1464 = 8'h70 == total_offset_7 ? phv_data_112 : _GEN_1463; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1465 = 8'h71 == total_offset_7 ? phv_data_113 : _GEN_1464; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1466 = 8'h72 == total_offset_7 ? phv_data_114 : _GEN_1465; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1467 = 8'h73 == total_offset_7 ? phv_data_115 : _GEN_1466; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1468 = 8'h74 == total_offset_7 ? phv_data_116 : _GEN_1467; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1469 = 8'h75 == total_offset_7 ? phv_data_117 : _GEN_1468; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1470 = 8'h76 == total_offset_7 ? phv_data_118 : _GEN_1469; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1471 = 8'h77 == total_offset_7 ? phv_data_119 : _GEN_1470; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1472 = 8'h78 == total_offset_7 ? phv_data_120 : _GEN_1471; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1473 = 8'h79 == total_offset_7 ? phv_data_121 : _GEN_1472; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1474 = 8'h7a == total_offset_7 ? phv_data_122 : _GEN_1473; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1475 = 8'h7b == total_offset_7 ? phv_data_123 : _GEN_1474; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1476 = 8'h7c == total_offset_7 ? phv_data_124 : _GEN_1475; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1477 = 8'h7d == total_offset_7 ? phv_data_125 : _GEN_1476; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1478 = 8'h7e == total_offset_7 ? phv_data_126 : _GEN_1477; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1479 = 8'h7f == total_offset_7 ? phv_data_127 : _GEN_1478; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1480 = 8'h80 == total_offset_7 ? phv_data_128 : _GEN_1479; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1481 = 8'h81 == total_offset_7 ? phv_data_129 : _GEN_1480; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1482 = 8'h82 == total_offset_7 ? phv_data_130 : _GEN_1481; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1483 = 8'h83 == total_offset_7 ? phv_data_131 : _GEN_1482; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1484 = 8'h84 == total_offset_7 ? phv_data_132 : _GEN_1483; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1485 = 8'h85 == total_offset_7 ? phv_data_133 : _GEN_1484; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1486 = 8'h86 == total_offset_7 ? phv_data_134 : _GEN_1485; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1487 = 8'h87 == total_offset_7 ? phv_data_135 : _GEN_1486; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1488 = 8'h88 == total_offset_7 ? phv_data_136 : _GEN_1487; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1489 = 8'h89 == total_offset_7 ? phv_data_137 : _GEN_1488; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1490 = 8'h8a == total_offset_7 ? phv_data_138 : _GEN_1489; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1491 = 8'h8b == total_offset_7 ? phv_data_139 : _GEN_1490; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1492 = 8'h8c == total_offset_7 ? phv_data_140 : _GEN_1491; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1493 = 8'h8d == total_offset_7 ? phv_data_141 : _GEN_1492; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1494 = 8'h8e == total_offset_7 ? phv_data_142 : _GEN_1493; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1495 = 8'h8f == total_offset_7 ? phv_data_143 : _GEN_1494; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1496 = 8'h90 == total_offset_7 ? phv_data_144 : _GEN_1495; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1497 = 8'h91 == total_offset_7 ? phv_data_145 : _GEN_1496; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1498 = 8'h92 == total_offset_7 ? phv_data_146 : _GEN_1497; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1499 = 8'h93 == total_offset_7 ? phv_data_147 : _GEN_1498; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1500 = 8'h94 == total_offset_7 ? phv_data_148 : _GEN_1499; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1501 = 8'h95 == total_offset_7 ? phv_data_149 : _GEN_1500; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1502 = 8'h96 == total_offset_7 ? phv_data_150 : _GEN_1501; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1503 = 8'h97 == total_offset_7 ? phv_data_151 : _GEN_1502; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1504 = 8'h98 == total_offset_7 ? phv_data_152 : _GEN_1503; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1505 = 8'h99 == total_offset_7 ? phv_data_153 : _GEN_1504; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1506 = 8'h9a == total_offset_7 ? phv_data_154 : _GEN_1505; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1507 = 8'h9b == total_offset_7 ? phv_data_155 : _GEN_1506; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1508 = 8'h9c == total_offset_7 ? phv_data_156 : _GEN_1507; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1509 = 8'h9d == total_offset_7 ? phv_data_157 : _GEN_1508; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1510 = 8'h9e == total_offset_7 ? phv_data_158 : _GEN_1509; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes_1_0 = 8'h9f == total_offset_7 ? phv_data_159 : _GEN_1510; // @[executor.scala 197:66 executor.scala 197:66]
  wire [31:0] _io_field_out_1_T = {bytes_1_0,bytes_1_1,bytes_1_2,bytes_1_3}; // @[Cat.scala 30:58]
  wire [3:0] _io_mask_out_1_T = {_mask_3_T_10,mask_1_1,mask_1_2,mask_1_3}; // @[Cat.scala 30:58]
  wire [17:0] io_field_out_1_hi_4 = io_field_out_1_lo[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _io_field_out_1_T_4 = {io_field_out_1_hi_4,io_field_out_1_lo}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_1737 = 4'hb == opcode_1 ? _io_field_out_1_T_4 : 32'h0; // @[executor.scala 230:56 executor.scala 231:41]
  wire [1:0] _GEN_1738 = from_header_1 ? bias_1 : 2'h0; // @[executor.scala 178:36 executor.scala 203:36 executor.scala 174:29]
  wire [31:0] _GEN_1739 = from_header_1 ? _io_field_out_1_T : _GEN_1737; // @[executor.scala 178:36 executor.scala 204:37]
  wire [3:0] _GEN_1740 = from_header_1 ? _io_mask_out_1_T : 4'h0; // @[executor.scala 178:36 executor.scala 205:37 executor.scala 173:29]
  wire [3:0] opcode_2 = vliw_2[31:28]; // @[primitive.scala 9:44]
  wire [13:0] io_field_out_2_lo = vliw_2[13:0]; // @[primitive.scala 11:44]
  wire  from_header_2 = length_2 != 8'h0; // @[executor.scala 177:45]
  wire [5:0] total_offset_hi_2 = offset_2[7:2]; // @[executor.scala 191:57]
  wire [7:0] _ending_T_5 = offset_2 + length_2; // @[executor.scala 193:46]
  wire [1:0] ending_2 = _ending_T_5[1:0]; // @[executor.scala 193:58]
  wire [3:0] _GEN_3502 = {{2'd0}, ending_2}; // @[executor.scala 194:45]
  wire [3:0] _bias_T_5 = 4'h4 - _GEN_3502; // @[executor.scala 194:45]
  wire [1:0] bias_2 = _bias_T_5[1:0]; // @[executor.scala 194:54]
  wire [7:0] total_offset_8 = {total_offset_hi_2,2'h0}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_1745 = 8'h1 == total_offset_8 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1746 = 8'h2 == total_offset_8 ? phv_data_2 : _GEN_1745; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1747 = 8'h3 == total_offset_8 ? phv_data_3 : _GEN_1746; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1748 = 8'h4 == total_offset_8 ? phv_data_4 : _GEN_1747; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1749 = 8'h5 == total_offset_8 ? phv_data_5 : _GEN_1748; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1750 = 8'h6 == total_offset_8 ? phv_data_6 : _GEN_1749; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1751 = 8'h7 == total_offset_8 ? phv_data_7 : _GEN_1750; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1752 = 8'h8 == total_offset_8 ? phv_data_8 : _GEN_1751; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1753 = 8'h9 == total_offset_8 ? phv_data_9 : _GEN_1752; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1754 = 8'ha == total_offset_8 ? phv_data_10 : _GEN_1753; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1755 = 8'hb == total_offset_8 ? phv_data_11 : _GEN_1754; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1756 = 8'hc == total_offset_8 ? phv_data_12 : _GEN_1755; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1757 = 8'hd == total_offset_8 ? phv_data_13 : _GEN_1756; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1758 = 8'he == total_offset_8 ? phv_data_14 : _GEN_1757; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1759 = 8'hf == total_offset_8 ? phv_data_15 : _GEN_1758; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1760 = 8'h10 == total_offset_8 ? phv_data_16 : _GEN_1759; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1761 = 8'h11 == total_offset_8 ? phv_data_17 : _GEN_1760; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1762 = 8'h12 == total_offset_8 ? phv_data_18 : _GEN_1761; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1763 = 8'h13 == total_offset_8 ? phv_data_19 : _GEN_1762; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1764 = 8'h14 == total_offset_8 ? phv_data_20 : _GEN_1763; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1765 = 8'h15 == total_offset_8 ? phv_data_21 : _GEN_1764; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1766 = 8'h16 == total_offset_8 ? phv_data_22 : _GEN_1765; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1767 = 8'h17 == total_offset_8 ? phv_data_23 : _GEN_1766; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1768 = 8'h18 == total_offset_8 ? phv_data_24 : _GEN_1767; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1769 = 8'h19 == total_offset_8 ? phv_data_25 : _GEN_1768; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1770 = 8'h1a == total_offset_8 ? phv_data_26 : _GEN_1769; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1771 = 8'h1b == total_offset_8 ? phv_data_27 : _GEN_1770; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1772 = 8'h1c == total_offset_8 ? phv_data_28 : _GEN_1771; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1773 = 8'h1d == total_offset_8 ? phv_data_29 : _GEN_1772; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1774 = 8'h1e == total_offset_8 ? phv_data_30 : _GEN_1773; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1775 = 8'h1f == total_offset_8 ? phv_data_31 : _GEN_1774; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1776 = 8'h20 == total_offset_8 ? phv_data_32 : _GEN_1775; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1777 = 8'h21 == total_offset_8 ? phv_data_33 : _GEN_1776; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1778 = 8'h22 == total_offset_8 ? phv_data_34 : _GEN_1777; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1779 = 8'h23 == total_offset_8 ? phv_data_35 : _GEN_1778; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1780 = 8'h24 == total_offset_8 ? phv_data_36 : _GEN_1779; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1781 = 8'h25 == total_offset_8 ? phv_data_37 : _GEN_1780; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1782 = 8'h26 == total_offset_8 ? phv_data_38 : _GEN_1781; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1783 = 8'h27 == total_offset_8 ? phv_data_39 : _GEN_1782; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1784 = 8'h28 == total_offset_8 ? phv_data_40 : _GEN_1783; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1785 = 8'h29 == total_offset_8 ? phv_data_41 : _GEN_1784; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1786 = 8'h2a == total_offset_8 ? phv_data_42 : _GEN_1785; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1787 = 8'h2b == total_offset_8 ? phv_data_43 : _GEN_1786; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1788 = 8'h2c == total_offset_8 ? phv_data_44 : _GEN_1787; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1789 = 8'h2d == total_offset_8 ? phv_data_45 : _GEN_1788; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1790 = 8'h2e == total_offset_8 ? phv_data_46 : _GEN_1789; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1791 = 8'h2f == total_offset_8 ? phv_data_47 : _GEN_1790; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1792 = 8'h30 == total_offset_8 ? phv_data_48 : _GEN_1791; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1793 = 8'h31 == total_offset_8 ? phv_data_49 : _GEN_1792; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1794 = 8'h32 == total_offset_8 ? phv_data_50 : _GEN_1793; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1795 = 8'h33 == total_offset_8 ? phv_data_51 : _GEN_1794; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1796 = 8'h34 == total_offset_8 ? phv_data_52 : _GEN_1795; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1797 = 8'h35 == total_offset_8 ? phv_data_53 : _GEN_1796; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1798 = 8'h36 == total_offset_8 ? phv_data_54 : _GEN_1797; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1799 = 8'h37 == total_offset_8 ? phv_data_55 : _GEN_1798; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1800 = 8'h38 == total_offset_8 ? phv_data_56 : _GEN_1799; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1801 = 8'h39 == total_offset_8 ? phv_data_57 : _GEN_1800; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1802 = 8'h3a == total_offset_8 ? phv_data_58 : _GEN_1801; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1803 = 8'h3b == total_offset_8 ? phv_data_59 : _GEN_1802; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1804 = 8'h3c == total_offset_8 ? phv_data_60 : _GEN_1803; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1805 = 8'h3d == total_offset_8 ? phv_data_61 : _GEN_1804; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1806 = 8'h3e == total_offset_8 ? phv_data_62 : _GEN_1805; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1807 = 8'h3f == total_offset_8 ? phv_data_63 : _GEN_1806; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1808 = 8'h40 == total_offset_8 ? phv_data_64 : _GEN_1807; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1809 = 8'h41 == total_offset_8 ? phv_data_65 : _GEN_1808; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1810 = 8'h42 == total_offset_8 ? phv_data_66 : _GEN_1809; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1811 = 8'h43 == total_offset_8 ? phv_data_67 : _GEN_1810; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1812 = 8'h44 == total_offset_8 ? phv_data_68 : _GEN_1811; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1813 = 8'h45 == total_offset_8 ? phv_data_69 : _GEN_1812; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1814 = 8'h46 == total_offset_8 ? phv_data_70 : _GEN_1813; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1815 = 8'h47 == total_offset_8 ? phv_data_71 : _GEN_1814; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1816 = 8'h48 == total_offset_8 ? phv_data_72 : _GEN_1815; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1817 = 8'h49 == total_offset_8 ? phv_data_73 : _GEN_1816; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1818 = 8'h4a == total_offset_8 ? phv_data_74 : _GEN_1817; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1819 = 8'h4b == total_offset_8 ? phv_data_75 : _GEN_1818; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1820 = 8'h4c == total_offset_8 ? phv_data_76 : _GEN_1819; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1821 = 8'h4d == total_offset_8 ? phv_data_77 : _GEN_1820; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1822 = 8'h4e == total_offset_8 ? phv_data_78 : _GEN_1821; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1823 = 8'h4f == total_offset_8 ? phv_data_79 : _GEN_1822; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1824 = 8'h50 == total_offset_8 ? phv_data_80 : _GEN_1823; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1825 = 8'h51 == total_offset_8 ? phv_data_81 : _GEN_1824; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1826 = 8'h52 == total_offset_8 ? phv_data_82 : _GEN_1825; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1827 = 8'h53 == total_offset_8 ? phv_data_83 : _GEN_1826; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1828 = 8'h54 == total_offset_8 ? phv_data_84 : _GEN_1827; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1829 = 8'h55 == total_offset_8 ? phv_data_85 : _GEN_1828; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1830 = 8'h56 == total_offset_8 ? phv_data_86 : _GEN_1829; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1831 = 8'h57 == total_offset_8 ? phv_data_87 : _GEN_1830; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1832 = 8'h58 == total_offset_8 ? phv_data_88 : _GEN_1831; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1833 = 8'h59 == total_offset_8 ? phv_data_89 : _GEN_1832; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1834 = 8'h5a == total_offset_8 ? phv_data_90 : _GEN_1833; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1835 = 8'h5b == total_offset_8 ? phv_data_91 : _GEN_1834; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1836 = 8'h5c == total_offset_8 ? phv_data_92 : _GEN_1835; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1837 = 8'h5d == total_offset_8 ? phv_data_93 : _GEN_1836; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1838 = 8'h5e == total_offset_8 ? phv_data_94 : _GEN_1837; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1839 = 8'h5f == total_offset_8 ? phv_data_95 : _GEN_1838; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1840 = 8'h60 == total_offset_8 ? phv_data_96 : _GEN_1839; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1841 = 8'h61 == total_offset_8 ? phv_data_97 : _GEN_1840; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1842 = 8'h62 == total_offset_8 ? phv_data_98 : _GEN_1841; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1843 = 8'h63 == total_offset_8 ? phv_data_99 : _GEN_1842; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1844 = 8'h64 == total_offset_8 ? phv_data_100 : _GEN_1843; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1845 = 8'h65 == total_offset_8 ? phv_data_101 : _GEN_1844; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1846 = 8'h66 == total_offset_8 ? phv_data_102 : _GEN_1845; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1847 = 8'h67 == total_offset_8 ? phv_data_103 : _GEN_1846; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1848 = 8'h68 == total_offset_8 ? phv_data_104 : _GEN_1847; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1849 = 8'h69 == total_offset_8 ? phv_data_105 : _GEN_1848; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1850 = 8'h6a == total_offset_8 ? phv_data_106 : _GEN_1849; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1851 = 8'h6b == total_offset_8 ? phv_data_107 : _GEN_1850; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1852 = 8'h6c == total_offset_8 ? phv_data_108 : _GEN_1851; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1853 = 8'h6d == total_offset_8 ? phv_data_109 : _GEN_1852; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1854 = 8'h6e == total_offset_8 ? phv_data_110 : _GEN_1853; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1855 = 8'h6f == total_offset_8 ? phv_data_111 : _GEN_1854; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1856 = 8'h70 == total_offset_8 ? phv_data_112 : _GEN_1855; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1857 = 8'h71 == total_offset_8 ? phv_data_113 : _GEN_1856; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1858 = 8'h72 == total_offset_8 ? phv_data_114 : _GEN_1857; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1859 = 8'h73 == total_offset_8 ? phv_data_115 : _GEN_1858; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1860 = 8'h74 == total_offset_8 ? phv_data_116 : _GEN_1859; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1861 = 8'h75 == total_offset_8 ? phv_data_117 : _GEN_1860; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1862 = 8'h76 == total_offset_8 ? phv_data_118 : _GEN_1861; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1863 = 8'h77 == total_offset_8 ? phv_data_119 : _GEN_1862; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1864 = 8'h78 == total_offset_8 ? phv_data_120 : _GEN_1863; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1865 = 8'h79 == total_offset_8 ? phv_data_121 : _GEN_1864; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1866 = 8'h7a == total_offset_8 ? phv_data_122 : _GEN_1865; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1867 = 8'h7b == total_offset_8 ? phv_data_123 : _GEN_1866; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1868 = 8'h7c == total_offset_8 ? phv_data_124 : _GEN_1867; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1869 = 8'h7d == total_offset_8 ? phv_data_125 : _GEN_1868; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1870 = 8'h7e == total_offset_8 ? phv_data_126 : _GEN_1869; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1871 = 8'h7f == total_offset_8 ? phv_data_127 : _GEN_1870; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1872 = 8'h80 == total_offset_8 ? phv_data_128 : _GEN_1871; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1873 = 8'h81 == total_offset_8 ? phv_data_129 : _GEN_1872; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1874 = 8'h82 == total_offset_8 ? phv_data_130 : _GEN_1873; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1875 = 8'h83 == total_offset_8 ? phv_data_131 : _GEN_1874; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1876 = 8'h84 == total_offset_8 ? phv_data_132 : _GEN_1875; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1877 = 8'h85 == total_offset_8 ? phv_data_133 : _GEN_1876; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1878 = 8'h86 == total_offset_8 ? phv_data_134 : _GEN_1877; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1879 = 8'h87 == total_offset_8 ? phv_data_135 : _GEN_1878; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1880 = 8'h88 == total_offset_8 ? phv_data_136 : _GEN_1879; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1881 = 8'h89 == total_offset_8 ? phv_data_137 : _GEN_1880; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1882 = 8'h8a == total_offset_8 ? phv_data_138 : _GEN_1881; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1883 = 8'h8b == total_offset_8 ? phv_data_139 : _GEN_1882; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1884 = 8'h8c == total_offset_8 ? phv_data_140 : _GEN_1883; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1885 = 8'h8d == total_offset_8 ? phv_data_141 : _GEN_1884; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1886 = 8'h8e == total_offset_8 ? phv_data_142 : _GEN_1885; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1887 = 8'h8f == total_offset_8 ? phv_data_143 : _GEN_1886; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1888 = 8'h90 == total_offset_8 ? phv_data_144 : _GEN_1887; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1889 = 8'h91 == total_offset_8 ? phv_data_145 : _GEN_1888; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1890 = 8'h92 == total_offset_8 ? phv_data_146 : _GEN_1889; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1891 = 8'h93 == total_offset_8 ? phv_data_147 : _GEN_1890; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1892 = 8'h94 == total_offset_8 ? phv_data_148 : _GEN_1891; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1893 = 8'h95 == total_offset_8 ? phv_data_149 : _GEN_1892; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1894 = 8'h96 == total_offset_8 ? phv_data_150 : _GEN_1893; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1895 = 8'h97 == total_offset_8 ? phv_data_151 : _GEN_1894; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1896 = 8'h98 == total_offset_8 ? phv_data_152 : _GEN_1895; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1897 = 8'h99 == total_offset_8 ? phv_data_153 : _GEN_1896; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1898 = 8'h9a == total_offset_8 ? phv_data_154 : _GEN_1897; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1899 = 8'h9b == total_offset_8 ? phv_data_155 : _GEN_1898; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1900 = 8'h9c == total_offset_8 ? phv_data_156 : _GEN_1899; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1901 = 8'h9d == total_offset_8 ? phv_data_157 : _GEN_1900; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1902 = 8'h9e == total_offset_8 ? phv_data_158 : _GEN_1901; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes_2_3 = 8'h9f == total_offset_8 ? phv_data_159 : _GEN_1902; // @[executor.scala 197:66 executor.scala 197:66]
  wire  _mask_3_T_17 = ending_2 == 2'h0; // @[executor.scala 199:88]
  wire  mask_2_3 = 2'h0 >= offset_2[1:0] & (2'h0 < ending_2 | ending_2 == 2'h0); // @[executor.scala 199:56]
  wire [7:0] total_offset_9 = {total_offset_hi_2,2'h1}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_1905 = 8'h1 == total_offset_9 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1906 = 8'h2 == total_offset_9 ? phv_data_2 : _GEN_1905; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1907 = 8'h3 == total_offset_9 ? phv_data_3 : _GEN_1906; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1908 = 8'h4 == total_offset_9 ? phv_data_4 : _GEN_1907; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1909 = 8'h5 == total_offset_9 ? phv_data_5 : _GEN_1908; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1910 = 8'h6 == total_offset_9 ? phv_data_6 : _GEN_1909; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1911 = 8'h7 == total_offset_9 ? phv_data_7 : _GEN_1910; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1912 = 8'h8 == total_offset_9 ? phv_data_8 : _GEN_1911; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1913 = 8'h9 == total_offset_9 ? phv_data_9 : _GEN_1912; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1914 = 8'ha == total_offset_9 ? phv_data_10 : _GEN_1913; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1915 = 8'hb == total_offset_9 ? phv_data_11 : _GEN_1914; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1916 = 8'hc == total_offset_9 ? phv_data_12 : _GEN_1915; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1917 = 8'hd == total_offset_9 ? phv_data_13 : _GEN_1916; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1918 = 8'he == total_offset_9 ? phv_data_14 : _GEN_1917; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1919 = 8'hf == total_offset_9 ? phv_data_15 : _GEN_1918; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1920 = 8'h10 == total_offset_9 ? phv_data_16 : _GEN_1919; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1921 = 8'h11 == total_offset_9 ? phv_data_17 : _GEN_1920; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1922 = 8'h12 == total_offset_9 ? phv_data_18 : _GEN_1921; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1923 = 8'h13 == total_offset_9 ? phv_data_19 : _GEN_1922; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1924 = 8'h14 == total_offset_9 ? phv_data_20 : _GEN_1923; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1925 = 8'h15 == total_offset_9 ? phv_data_21 : _GEN_1924; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1926 = 8'h16 == total_offset_9 ? phv_data_22 : _GEN_1925; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1927 = 8'h17 == total_offset_9 ? phv_data_23 : _GEN_1926; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1928 = 8'h18 == total_offset_9 ? phv_data_24 : _GEN_1927; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1929 = 8'h19 == total_offset_9 ? phv_data_25 : _GEN_1928; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1930 = 8'h1a == total_offset_9 ? phv_data_26 : _GEN_1929; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1931 = 8'h1b == total_offset_9 ? phv_data_27 : _GEN_1930; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1932 = 8'h1c == total_offset_9 ? phv_data_28 : _GEN_1931; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1933 = 8'h1d == total_offset_9 ? phv_data_29 : _GEN_1932; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1934 = 8'h1e == total_offset_9 ? phv_data_30 : _GEN_1933; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1935 = 8'h1f == total_offset_9 ? phv_data_31 : _GEN_1934; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1936 = 8'h20 == total_offset_9 ? phv_data_32 : _GEN_1935; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1937 = 8'h21 == total_offset_9 ? phv_data_33 : _GEN_1936; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1938 = 8'h22 == total_offset_9 ? phv_data_34 : _GEN_1937; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1939 = 8'h23 == total_offset_9 ? phv_data_35 : _GEN_1938; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1940 = 8'h24 == total_offset_9 ? phv_data_36 : _GEN_1939; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1941 = 8'h25 == total_offset_9 ? phv_data_37 : _GEN_1940; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1942 = 8'h26 == total_offset_9 ? phv_data_38 : _GEN_1941; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1943 = 8'h27 == total_offset_9 ? phv_data_39 : _GEN_1942; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1944 = 8'h28 == total_offset_9 ? phv_data_40 : _GEN_1943; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1945 = 8'h29 == total_offset_9 ? phv_data_41 : _GEN_1944; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1946 = 8'h2a == total_offset_9 ? phv_data_42 : _GEN_1945; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1947 = 8'h2b == total_offset_9 ? phv_data_43 : _GEN_1946; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1948 = 8'h2c == total_offset_9 ? phv_data_44 : _GEN_1947; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1949 = 8'h2d == total_offset_9 ? phv_data_45 : _GEN_1948; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1950 = 8'h2e == total_offset_9 ? phv_data_46 : _GEN_1949; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1951 = 8'h2f == total_offset_9 ? phv_data_47 : _GEN_1950; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1952 = 8'h30 == total_offset_9 ? phv_data_48 : _GEN_1951; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1953 = 8'h31 == total_offset_9 ? phv_data_49 : _GEN_1952; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1954 = 8'h32 == total_offset_9 ? phv_data_50 : _GEN_1953; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1955 = 8'h33 == total_offset_9 ? phv_data_51 : _GEN_1954; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1956 = 8'h34 == total_offset_9 ? phv_data_52 : _GEN_1955; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1957 = 8'h35 == total_offset_9 ? phv_data_53 : _GEN_1956; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1958 = 8'h36 == total_offset_9 ? phv_data_54 : _GEN_1957; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1959 = 8'h37 == total_offset_9 ? phv_data_55 : _GEN_1958; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1960 = 8'h38 == total_offset_9 ? phv_data_56 : _GEN_1959; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1961 = 8'h39 == total_offset_9 ? phv_data_57 : _GEN_1960; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1962 = 8'h3a == total_offset_9 ? phv_data_58 : _GEN_1961; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1963 = 8'h3b == total_offset_9 ? phv_data_59 : _GEN_1962; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1964 = 8'h3c == total_offset_9 ? phv_data_60 : _GEN_1963; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1965 = 8'h3d == total_offset_9 ? phv_data_61 : _GEN_1964; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1966 = 8'h3e == total_offset_9 ? phv_data_62 : _GEN_1965; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1967 = 8'h3f == total_offset_9 ? phv_data_63 : _GEN_1966; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1968 = 8'h40 == total_offset_9 ? phv_data_64 : _GEN_1967; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1969 = 8'h41 == total_offset_9 ? phv_data_65 : _GEN_1968; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1970 = 8'h42 == total_offset_9 ? phv_data_66 : _GEN_1969; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1971 = 8'h43 == total_offset_9 ? phv_data_67 : _GEN_1970; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1972 = 8'h44 == total_offset_9 ? phv_data_68 : _GEN_1971; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1973 = 8'h45 == total_offset_9 ? phv_data_69 : _GEN_1972; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1974 = 8'h46 == total_offset_9 ? phv_data_70 : _GEN_1973; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1975 = 8'h47 == total_offset_9 ? phv_data_71 : _GEN_1974; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1976 = 8'h48 == total_offset_9 ? phv_data_72 : _GEN_1975; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1977 = 8'h49 == total_offset_9 ? phv_data_73 : _GEN_1976; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1978 = 8'h4a == total_offset_9 ? phv_data_74 : _GEN_1977; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1979 = 8'h4b == total_offset_9 ? phv_data_75 : _GEN_1978; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1980 = 8'h4c == total_offset_9 ? phv_data_76 : _GEN_1979; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1981 = 8'h4d == total_offset_9 ? phv_data_77 : _GEN_1980; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1982 = 8'h4e == total_offset_9 ? phv_data_78 : _GEN_1981; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1983 = 8'h4f == total_offset_9 ? phv_data_79 : _GEN_1982; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1984 = 8'h50 == total_offset_9 ? phv_data_80 : _GEN_1983; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1985 = 8'h51 == total_offset_9 ? phv_data_81 : _GEN_1984; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1986 = 8'h52 == total_offset_9 ? phv_data_82 : _GEN_1985; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1987 = 8'h53 == total_offset_9 ? phv_data_83 : _GEN_1986; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1988 = 8'h54 == total_offset_9 ? phv_data_84 : _GEN_1987; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1989 = 8'h55 == total_offset_9 ? phv_data_85 : _GEN_1988; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1990 = 8'h56 == total_offset_9 ? phv_data_86 : _GEN_1989; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1991 = 8'h57 == total_offset_9 ? phv_data_87 : _GEN_1990; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1992 = 8'h58 == total_offset_9 ? phv_data_88 : _GEN_1991; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1993 = 8'h59 == total_offset_9 ? phv_data_89 : _GEN_1992; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1994 = 8'h5a == total_offset_9 ? phv_data_90 : _GEN_1993; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1995 = 8'h5b == total_offset_9 ? phv_data_91 : _GEN_1994; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1996 = 8'h5c == total_offset_9 ? phv_data_92 : _GEN_1995; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1997 = 8'h5d == total_offset_9 ? phv_data_93 : _GEN_1996; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1998 = 8'h5e == total_offset_9 ? phv_data_94 : _GEN_1997; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1999 = 8'h5f == total_offset_9 ? phv_data_95 : _GEN_1998; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2000 = 8'h60 == total_offset_9 ? phv_data_96 : _GEN_1999; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2001 = 8'h61 == total_offset_9 ? phv_data_97 : _GEN_2000; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2002 = 8'h62 == total_offset_9 ? phv_data_98 : _GEN_2001; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2003 = 8'h63 == total_offset_9 ? phv_data_99 : _GEN_2002; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2004 = 8'h64 == total_offset_9 ? phv_data_100 : _GEN_2003; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2005 = 8'h65 == total_offset_9 ? phv_data_101 : _GEN_2004; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2006 = 8'h66 == total_offset_9 ? phv_data_102 : _GEN_2005; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2007 = 8'h67 == total_offset_9 ? phv_data_103 : _GEN_2006; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2008 = 8'h68 == total_offset_9 ? phv_data_104 : _GEN_2007; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2009 = 8'h69 == total_offset_9 ? phv_data_105 : _GEN_2008; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2010 = 8'h6a == total_offset_9 ? phv_data_106 : _GEN_2009; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2011 = 8'h6b == total_offset_9 ? phv_data_107 : _GEN_2010; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2012 = 8'h6c == total_offset_9 ? phv_data_108 : _GEN_2011; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2013 = 8'h6d == total_offset_9 ? phv_data_109 : _GEN_2012; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2014 = 8'h6e == total_offset_9 ? phv_data_110 : _GEN_2013; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2015 = 8'h6f == total_offset_9 ? phv_data_111 : _GEN_2014; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2016 = 8'h70 == total_offset_9 ? phv_data_112 : _GEN_2015; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2017 = 8'h71 == total_offset_9 ? phv_data_113 : _GEN_2016; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2018 = 8'h72 == total_offset_9 ? phv_data_114 : _GEN_2017; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2019 = 8'h73 == total_offset_9 ? phv_data_115 : _GEN_2018; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2020 = 8'h74 == total_offset_9 ? phv_data_116 : _GEN_2019; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2021 = 8'h75 == total_offset_9 ? phv_data_117 : _GEN_2020; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2022 = 8'h76 == total_offset_9 ? phv_data_118 : _GEN_2021; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2023 = 8'h77 == total_offset_9 ? phv_data_119 : _GEN_2022; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2024 = 8'h78 == total_offset_9 ? phv_data_120 : _GEN_2023; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2025 = 8'h79 == total_offset_9 ? phv_data_121 : _GEN_2024; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2026 = 8'h7a == total_offset_9 ? phv_data_122 : _GEN_2025; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2027 = 8'h7b == total_offset_9 ? phv_data_123 : _GEN_2026; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2028 = 8'h7c == total_offset_9 ? phv_data_124 : _GEN_2027; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2029 = 8'h7d == total_offset_9 ? phv_data_125 : _GEN_2028; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2030 = 8'h7e == total_offset_9 ? phv_data_126 : _GEN_2029; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2031 = 8'h7f == total_offset_9 ? phv_data_127 : _GEN_2030; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2032 = 8'h80 == total_offset_9 ? phv_data_128 : _GEN_2031; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2033 = 8'h81 == total_offset_9 ? phv_data_129 : _GEN_2032; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2034 = 8'h82 == total_offset_9 ? phv_data_130 : _GEN_2033; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2035 = 8'h83 == total_offset_9 ? phv_data_131 : _GEN_2034; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2036 = 8'h84 == total_offset_9 ? phv_data_132 : _GEN_2035; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2037 = 8'h85 == total_offset_9 ? phv_data_133 : _GEN_2036; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2038 = 8'h86 == total_offset_9 ? phv_data_134 : _GEN_2037; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2039 = 8'h87 == total_offset_9 ? phv_data_135 : _GEN_2038; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2040 = 8'h88 == total_offset_9 ? phv_data_136 : _GEN_2039; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2041 = 8'h89 == total_offset_9 ? phv_data_137 : _GEN_2040; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2042 = 8'h8a == total_offset_9 ? phv_data_138 : _GEN_2041; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2043 = 8'h8b == total_offset_9 ? phv_data_139 : _GEN_2042; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2044 = 8'h8c == total_offset_9 ? phv_data_140 : _GEN_2043; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2045 = 8'h8d == total_offset_9 ? phv_data_141 : _GEN_2044; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2046 = 8'h8e == total_offset_9 ? phv_data_142 : _GEN_2045; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2047 = 8'h8f == total_offset_9 ? phv_data_143 : _GEN_2046; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2048 = 8'h90 == total_offset_9 ? phv_data_144 : _GEN_2047; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2049 = 8'h91 == total_offset_9 ? phv_data_145 : _GEN_2048; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2050 = 8'h92 == total_offset_9 ? phv_data_146 : _GEN_2049; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2051 = 8'h93 == total_offset_9 ? phv_data_147 : _GEN_2050; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2052 = 8'h94 == total_offset_9 ? phv_data_148 : _GEN_2051; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2053 = 8'h95 == total_offset_9 ? phv_data_149 : _GEN_2052; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2054 = 8'h96 == total_offset_9 ? phv_data_150 : _GEN_2053; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2055 = 8'h97 == total_offset_9 ? phv_data_151 : _GEN_2054; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2056 = 8'h98 == total_offset_9 ? phv_data_152 : _GEN_2055; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2057 = 8'h99 == total_offset_9 ? phv_data_153 : _GEN_2056; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2058 = 8'h9a == total_offset_9 ? phv_data_154 : _GEN_2057; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2059 = 8'h9b == total_offset_9 ? phv_data_155 : _GEN_2058; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2060 = 8'h9c == total_offset_9 ? phv_data_156 : _GEN_2059; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2061 = 8'h9d == total_offset_9 ? phv_data_157 : _GEN_2060; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2062 = 8'h9e == total_offset_9 ? phv_data_158 : _GEN_2061; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes_2_2 = 8'h9f == total_offset_9 ? phv_data_159 : _GEN_2062; // @[executor.scala 197:66 executor.scala 197:66]
  wire  mask_2_2 = 2'h1 >= offset_2[1:0] & (2'h1 < ending_2 | ending_2 == 2'h0); // @[executor.scala 199:56]
  wire [7:0] total_offset_10 = {total_offset_hi_2,2'h2}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_2065 = 8'h1 == total_offset_10 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2066 = 8'h2 == total_offset_10 ? phv_data_2 : _GEN_2065; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2067 = 8'h3 == total_offset_10 ? phv_data_3 : _GEN_2066; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2068 = 8'h4 == total_offset_10 ? phv_data_4 : _GEN_2067; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2069 = 8'h5 == total_offset_10 ? phv_data_5 : _GEN_2068; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2070 = 8'h6 == total_offset_10 ? phv_data_6 : _GEN_2069; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2071 = 8'h7 == total_offset_10 ? phv_data_7 : _GEN_2070; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2072 = 8'h8 == total_offset_10 ? phv_data_8 : _GEN_2071; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2073 = 8'h9 == total_offset_10 ? phv_data_9 : _GEN_2072; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2074 = 8'ha == total_offset_10 ? phv_data_10 : _GEN_2073; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2075 = 8'hb == total_offset_10 ? phv_data_11 : _GEN_2074; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2076 = 8'hc == total_offset_10 ? phv_data_12 : _GEN_2075; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2077 = 8'hd == total_offset_10 ? phv_data_13 : _GEN_2076; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2078 = 8'he == total_offset_10 ? phv_data_14 : _GEN_2077; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2079 = 8'hf == total_offset_10 ? phv_data_15 : _GEN_2078; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2080 = 8'h10 == total_offset_10 ? phv_data_16 : _GEN_2079; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2081 = 8'h11 == total_offset_10 ? phv_data_17 : _GEN_2080; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2082 = 8'h12 == total_offset_10 ? phv_data_18 : _GEN_2081; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2083 = 8'h13 == total_offset_10 ? phv_data_19 : _GEN_2082; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2084 = 8'h14 == total_offset_10 ? phv_data_20 : _GEN_2083; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2085 = 8'h15 == total_offset_10 ? phv_data_21 : _GEN_2084; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2086 = 8'h16 == total_offset_10 ? phv_data_22 : _GEN_2085; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2087 = 8'h17 == total_offset_10 ? phv_data_23 : _GEN_2086; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2088 = 8'h18 == total_offset_10 ? phv_data_24 : _GEN_2087; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2089 = 8'h19 == total_offset_10 ? phv_data_25 : _GEN_2088; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2090 = 8'h1a == total_offset_10 ? phv_data_26 : _GEN_2089; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2091 = 8'h1b == total_offset_10 ? phv_data_27 : _GEN_2090; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2092 = 8'h1c == total_offset_10 ? phv_data_28 : _GEN_2091; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2093 = 8'h1d == total_offset_10 ? phv_data_29 : _GEN_2092; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2094 = 8'h1e == total_offset_10 ? phv_data_30 : _GEN_2093; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2095 = 8'h1f == total_offset_10 ? phv_data_31 : _GEN_2094; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2096 = 8'h20 == total_offset_10 ? phv_data_32 : _GEN_2095; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2097 = 8'h21 == total_offset_10 ? phv_data_33 : _GEN_2096; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2098 = 8'h22 == total_offset_10 ? phv_data_34 : _GEN_2097; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2099 = 8'h23 == total_offset_10 ? phv_data_35 : _GEN_2098; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2100 = 8'h24 == total_offset_10 ? phv_data_36 : _GEN_2099; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2101 = 8'h25 == total_offset_10 ? phv_data_37 : _GEN_2100; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2102 = 8'h26 == total_offset_10 ? phv_data_38 : _GEN_2101; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2103 = 8'h27 == total_offset_10 ? phv_data_39 : _GEN_2102; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2104 = 8'h28 == total_offset_10 ? phv_data_40 : _GEN_2103; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2105 = 8'h29 == total_offset_10 ? phv_data_41 : _GEN_2104; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2106 = 8'h2a == total_offset_10 ? phv_data_42 : _GEN_2105; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2107 = 8'h2b == total_offset_10 ? phv_data_43 : _GEN_2106; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2108 = 8'h2c == total_offset_10 ? phv_data_44 : _GEN_2107; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2109 = 8'h2d == total_offset_10 ? phv_data_45 : _GEN_2108; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2110 = 8'h2e == total_offset_10 ? phv_data_46 : _GEN_2109; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2111 = 8'h2f == total_offset_10 ? phv_data_47 : _GEN_2110; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2112 = 8'h30 == total_offset_10 ? phv_data_48 : _GEN_2111; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2113 = 8'h31 == total_offset_10 ? phv_data_49 : _GEN_2112; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2114 = 8'h32 == total_offset_10 ? phv_data_50 : _GEN_2113; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2115 = 8'h33 == total_offset_10 ? phv_data_51 : _GEN_2114; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2116 = 8'h34 == total_offset_10 ? phv_data_52 : _GEN_2115; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2117 = 8'h35 == total_offset_10 ? phv_data_53 : _GEN_2116; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2118 = 8'h36 == total_offset_10 ? phv_data_54 : _GEN_2117; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2119 = 8'h37 == total_offset_10 ? phv_data_55 : _GEN_2118; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2120 = 8'h38 == total_offset_10 ? phv_data_56 : _GEN_2119; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2121 = 8'h39 == total_offset_10 ? phv_data_57 : _GEN_2120; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2122 = 8'h3a == total_offset_10 ? phv_data_58 : _GEN_2121; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2123 = 8'h3b == total_offset_10 ? phv_data_59 : _GEN_2122; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2124 = 8'h3c == total_offset_10 ? phv_data_60 : _GEN_2123; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2125 = 8'h3d == total_offset_10 ? phv_data_61 : _GEN_2124; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2126 = 8'h3e == total_offset_10 ? phv_data_62 : _GEN_2125; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2127 = 8'h3f == total_offset_10 ? phv_data_63 : _GEN_2126; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2128 = 8'h40 == total_offset_10 ? phv_data_64 : _GEN_2127; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2129 = 8'h41 == total_offset_10 ? phv_data_65 : _GEN_2128; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2130 = 8'h42 == total_offset_10 ? phv_data_66 : _GEN_2129; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2131 = 8'h43 == total_offset_10 ? phv_data_67 : _GEN_2130; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2132 = 8'h44 == total_offset_10 ? phv_data_68 : _GEN_2131; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2133 = 8'h45 == total_offset_10 ? phv_data_69 : _GEN_2132; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2134 = 8'h46 == total_offset_10 ? phv_data_70 : _GEN_2133; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2135 = 8'h47 == total_offset_10 ? phv_data_71 : _GEN_2134; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2136 = 8'h48 == total_offset_10 ? phv_data_72 : _GEN_2135; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2137 = 8'h49 == total_offset_10 ? phv_data_73 : _GEN_2136; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2138 = 8'h4a == total_offset_10 ? phv_data_74 : _GEN_2137; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2139 = 8'h4b == total_offset_10 ? phv_data_75 : _GEN_2138; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2140 = 8'h4c == total_offset_10 ? phv_data_76 : _GEN_2139; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2141 = 8'h4d == total_offset_10 ? phv_data_77 : _GEN_2140; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2142 = 8'h4e == total_offset_10 ? phv_data_78 : _GEN_2141; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2143 = 8'h4f == total_offset_10 ? phv_data_79 : _GEN_2142; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2144 = 8'h50 == total_offset_10 ? phv_data_80 : _GEN_2143; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2145 = 8'h51 == total_offset_10 ? phv_data_81 : _GEN_2144; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2146 = 8'h52 == total_offset_10 ? phv_data_82 : _GEN_2145; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2147 = 8'h53 == total_offset_10 ? phv_data_83 : _GEN_2146; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2148 = 8'h54 == total_offset_10 ? phv_data_84 : _GEN_2147; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2149 = 8'h55 == total_offset_10 ? phv_data_85 : _GEN_2148; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2150 = 8'h56 == total_offset_10 ? phv_data_86 : _GEN_2149; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2151 = 8'h57 == total_offset_10 ? phv_data_87 : _GEN_2150; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2152 = 8'h58 == total_offset_10 ? phv_data_88 : _GEN_2151; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2153 = 8'h59 == total_offset_10 ? phv_data_89 : _GEN_2152; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2154 = 8'h5a == total_offset_10 ? phv_data_90 : _GEN_2153; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2155 = 8'h5b == total_offset_10 ? phv_data_91 : _GEN_2154; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2156 = 8'h5c == total_offset_10 ? phv_data_92 : _GEN_2155; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2157 = 8'h5d == total_offset_10 ? phv_data_93 : _GEN_2156; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2158 = 8'h5e == total_offset_10 ? phv_data_94 : _GEN_2157; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2159 = 8'h5f == total_offset_10 ? phv_data_95 : _GEN_2158; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2160 = 8'h60 == total_offset_10 ? phv_data_96 : _GEN_2159; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2161 = 8'h61 == total_offset_10 ? phv_data_97 : _GEN_2160; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2162 = 8'h62 == total_offset_10 ? phv_data_98 : _GEN_2161; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2163 = 8'h63 == total_offset_10 ? phv_data_99 : _GEN_2162; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2164 = 8'h64 == total_offset_10 ? phv_data_100 : _GEN_2163; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2165 = 8'h65 == total_offset_10 ? phv_data_101 : _GEN_2164; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2166 = 8'h66 == total_offset_10 ? phv_data_102 : _GEN_2165; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2167 = 8'h67 == total_offset_10 ? phv_data_103 : _GEN_2166; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2168 = 8'h68 == total_offset_10 ? phv_data_104 : _GEN_2167; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2169 = 8'h69 == total_offset_10 ? phv_data_105 : _GEN_2168; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2170 = 8'h6a == total_offset_10 ? phv_data_106 : _GEN_2169; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2171 = 8'h6b == total_offset_10 ? phv_data_107 : _GEN_2170; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2172 = 8'h6c == total_offset_10 ? phv_data_108 : _GEN_2171; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2173 = 8'h6d == total_offset_10 ? phv_data_109 : _GEN_2172; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2174 = 8'h6e == total_offset_10 ? phv_data_110 : _GEN_2173; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2175 = 8'h6f == total_offset_10 ? phv_data_111 : _GEN_2174; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2176 = 8'h70 == total_offset_10 ? phv_data_112 : _GEN_2175; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2177 = 8'h71 == total_offset_10 ? phv_data_113 : _GEN_2176; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2178 = 8'h72 == total_offset_10 ? phv_data_114 : _GEN_2177; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2179 = 8'h73 == total_offset_10 ? phv_data_115 : _GEN_2178; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2180 = 8'h74 == total_offset_10 ? phv_data_116 : _GEN_2179; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2181 = 8'h75 == total_offset_10 ? phv_data_117 : _GEN_2180; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2182 = 8'h76 == total_offset_10 ? phv_data_118 : _GEN_2181; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2183 = 8'h77 == total_offset_10 ? phv_data_119 : _GEN_2182; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2184 = 8'h78 == total_offset_10 ? phv_data_120 : _GEN_2183; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2185 = 8'h79 == total_offset_10 ? phv_data_121 : _GEN_2184; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2186 = 8'h7a == total_offset_10 ? phv_data_122 : _GEN_2185; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2187 = 8'h7b == total_offset_10 ? phv_data_123 : _GEN_2186; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2188 = 8'h7c == total_offset_10 ? phv_data_124 : _GEN_2187; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2189 = 8'h7d == total_offset_10 ? phv_data_125 : _GEN_2188; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2190 = 8'h7e == total_offset_10 ? phv_data_126 : _GEN_2189; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2191 = 8'h7f == total_offset_10 ? phv_data_127 : _GEN_2190; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2192 = 8'h80 == total_offset_10 ? phv_data_128 : _GEN_2191; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2193 = 8'h81 == total_offset_10 ? phv_data_129 : _GEN_2192; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2194 = 8'h82 == total_offset_10 ? phv_data_130 : _GEN_2193; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2195 = 8'h83 == total_offset_10 ? phv_data_131 : _GEN_2194; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2196 = 8'h84 == total_offset_10 ? phv_data_132 : _GEN_2195; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2197 = 8'h85 == total_offset_10 ? phv_data_133 : _GEN_2196; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2198 = 8'h86 == total_offset_10 ? phv_data_134 : _GEN_2197; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2199 = 8'h87 == total_offset_10 ? phv_data_135 : _GEN_2198; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2200 = 8'h88 == total_offset_10 ? phv_data_136 : _GEN_2199; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2201 = 8'h89 == total_offset_10 ? phv_data_137 : _GEN_2200; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2202 = 8'h8a == total_offset_10 ? phv_data_138 : _GEN_2201; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2203 = 8'h8b == total_offset_10 ? phv_data_139 : _GEN_2202; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2204 = 8'h8c == total_offset_10 ? phv_data_140 : _GEN_2203; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2205 = 8'h8d == total_offset_10 ? phv_data_141 : _GEN_2204; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2206 = 8'h8e == total_offset_10 ? phv_data_142 : _GEN_2205; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2207 = 8'h8f == total_offset_10 ? phv_data_143 : _GEN_2206; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2208 = 8'h90 == total_offset_10 ? phv_data_144 : _GEN_2207; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2209 = 8'h91 == total_offset_10 ? phv_data_145 : _GEN_2208; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2210 = 8'h92 == total_offset_10 ? phv_data_146 : _GEN_2209; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2211 = 8'h93 == total_offset_10 ? phv_data_147 : _GEN_2210; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2212 = 8'h94 == total_offset_10 ? phv_data_148 : _GEN_2211; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2213 = 8'h95 == total_offset_10 ? phv_data_149 : _GEN_2212; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2214 = 8'h96 == total_offset_10 ? phv_data_150 : _GEN_2213; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2215 = 8'h97 == total_offset_10 ? phv_data_151 : _GEN_2214; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2216 = 8'h98 == total_offset_10 ? phv_data_152 : _GEN_2215; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2217 = 8'h99 == total_offset_10 ? phv_data_153 : _GEN_2216; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2218 = 8'h9a == total_offset_10 ? phv_data_154 : _GEN_2217; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2219 = 8'h9b == total_offset_10 ? phv_data_155 : _GEN_2218; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2220 = 8'h9c == total_offset_10 ? phv_data_156 : _GEN_2219; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2221 = 8'h9d == total_offset_10 ? phv_data_157 : _GEN_2220; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2222 = 8'h9e == total_offset_10 ? phv_data_158 : _GEN_2221; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes_2_1 = 8'h9f == total_offset_10 ? phv_data_159 : _GEN_2222; // @[executor.scala 197:66 executor.scala 197:66]
  wire  mask_2_1 = 2'h2 >= offset_2[1:0] & (2'h2 < ending_2 | ending_2 == 2'h0); // @[executor.scala 199:56]
  wire [7:0] total_offset_11 = {total_offset_hi_2,2'h3}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_2225 = 8'h1 == total_offset_11 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2226 = 8'h2 == total_offset_11 ? phv_data_2 : _GEN_2225; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2227 = 8'h3 == total_offset_11 ? phv_data_3 : _GEN_2226; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2228 = 8'h4 == total_offset_11 ? phv_data_4 : _GEN_2227; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2229 = 8'h5 == total_offset_11 ? phv_data_5 : _GEN_2228; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2230 = 8'h6 == total_offset_11 ? phv_data_6 : _GEN_2229; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2231 = 8'h7 == total_offset_11 ? phv_data_7 : _GEN_2230; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2232 = 8'h8 == total_offset_11 ? phv_data_8 : _GEN_2231; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2233 = 8'h9 == total_offset_11 ? phv_data_9 : _GEN_2232; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2234 = 8'ha == total_offset_11 ? phv_data_10 : _GEN_2233; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2235 = 8'hb == total_offset_11 ? phv_data_11 : _GEN_2234; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2236 = 8'hc == total_offset_11 ? phv_data_12 : _GEN_2235; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2237 = 8'hd == total_offset_11 ? phv_data_13 : _GEN_2236; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2238 = 8'he == total_offset_11 ? phv_data_14 : _GEN_2237; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2239 = 8'hf == total_offset_11 ? phv_data_15 : _GEN_2238; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2240 = 8'h10 == total_offset_11 ? phv_data_16 : _GEN_2239; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2241 = 8'h11 == total_offset_11 ? phv_data_17 : _GEN_2240; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2242 = 8'h12 == total_offset_11 ? phv_data_18 : _GEN_2241; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2243 = 8'h13 == total_offset_11 ? phv_data_19 : _GEN_2242; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2244 = 8'h14 == total_offset_11 ? phv_data_20 : _GEN_2243; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2245 = 8'h15 == total_offset_11 ? phv_data_21 : _GEN_2244; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2246 = 8'h16 == total_offset_11 ? phv_data_22 : _GEN_2245; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2247 = 8'h17 == total_offset_11 ? phv_data_23 : _GEN_2246; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2248 = 8'h18 == total_offset_11 ? phv_data_24 : _GEN_2247; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2249 = 8'h19 == total_offset_11 ? phv_data_25 : _GEN_2248; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2250 = 8'h1a == total_offset_11 ? phv_data_26 : _GEN_2249; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2251 = 8'h1b == total_offset_11 ? phv_data_27 : _GEN_2250; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2252 = 8'h1c == total_offset_11 ? phv_data_28 : _GEN_2251; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2253 = 8'h1d == total_offset_11 ? phv_data_29 : _GEN_2252; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2254 = 8'h1e == total_offset_11 ? phv_data_30 : _GEN_2253; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2255 = 8'h1f == total_offset_11 ? phv_data_31 : _GEN_2254; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2256 = 8'h20 == total_offset_11 ? phv_data_32 : _GEN_2255; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2257 = 8'h21 == total_offset_11 ? phv_data_33 : _GEN_2256; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2258 = 8'h22 == total_offset_11 ? phv_data_34 : _GEN_2257; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2259 = 8'h23 == total_offset_11 ? phv_data_35 : _GEN_2258; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2260 = 8'h24 == total_offset_11 ? phv_data_36 : _GEN_2259; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2261 = 8'h25 == total_offset_11 ? phv_data_37 : _GEN_2260; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2262 = 8'h26 == total_offset_11 ? phv_data_38 : _GEN_2261; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2263 = 8'h27 == total_offset_11 ? phv_data_39 : _GEN_2262; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2264 = 8'h28 == total_offset_11 ? phv_data_40 : _GEN_2263; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2265 = 8'h29 == total_offset_11 ? phv_data_41 : _GEN_2264; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2266 = 8'h2a == total_offset_11 ? phv_data_42 : _GEN_2265; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2267 = 8'h2b == total_offset_11 ? phv_data_43 : _GEN_2266; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2268 = 8'h2c == total_offset_11 ? phv_data_44 : _GEN_2267; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2269 = 8'h2d == total_offset_11 ? phv_data_45 : _GEN_2268; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2270 = 8'h2e == total_offset_11 ? phv_data_46 : _GEN_2269; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2271 = 8'h2f == total_offset_11 ? phv_data_47 : _GEN_2270; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2272 = 8'h30 == total_offset_11 ? phv_data_48 : _GEN_2271; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2273 = 8'h31 == total_offset_11 ? phv_data_49 : _GEN_2272; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2274 = 8'h32 == total_offset_11 ? phv_data_50 : _GEN_2273; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2275 = 8'h33 == total_offset_11 ? phv_data_51 : _GEN_2274; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2276 = 8'h34 == total_offset_11 ? phv_data_52 : _GEN_2275; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2277 = 8'h35 == total_offset_11 ? phv_data_53 : _GEN_2276; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2278 = 8'h36 == total_offset_11 ? phv_data_54 : _GEN_2277; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2279 = 8'h37 == total_offset_11 ? phv_data_55 : _GEN_2278; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2280 = 8'h38 == total_offset_11 ? phv_data_56 : _GEN_2279; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2281 = 8'h39 == total_offset_11 ? phv_data_57 : _GEN_2280; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2282 = 8'h3a == total_offset_11 ? phv_data_58 : _GEN_2281; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2283 = 8'h3b == total_offset_11 ? phv_data_59 : _GEN_2282; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2284 = 8'h3c == total_offset_11 ? phv_data_60 : _GEN_2283; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2285 = 8'h3d == total_offset_11 ? phv_data_61 : _GEN_2284; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2286 = 8'h3e == total_offset_11 ? phv_data_62 : _GEN_2285; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2287 = 8'h3f == total_offset_11 ? phv_data_63 : _GEN_2286; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2288 = 8'h40 == total_offset_11 ? phv_data_64 : _GEN_2287; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2289 = 8'h41 == total_offset_11 ? phv_data_65 : _GEN_2288; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2290 = 8'h42 == total_offset_11 ? phv_data_66 : _GEN_2289; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2291 = 8'h43 == total_offset_11 ? phv_data_67 : _GEN_2290; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2292 = 8'h44 == total_offset_11 ? phv_data_68 : _GEN_2291; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2293 = 8'h45 == total_offset_11 ? phv_data_69 : _GEN_2292; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2294 = 8'h46 == total_offset_11 ? phv_data_70 : _GEN_2293; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2295 = 8'h47 == total_offset_11 ? phv_data_71 : _GEN_2294; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2296 = 8'h48 == total_offset_11 ? phv_data_72 : _GEN_2295; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2297 = 8'h49 == total_offset_11 ? phv_data_73 : _GEN_2296; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2298 = 8'h4a == total_offset_11 ? phv_data_74 : _GEN_2297; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2299 = 8'h4b == total_offset_11 ? phv_data_75 : _GEN_2298; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2300 = 8'h4c == total_offset_11 ? phv_data_76 : _GEN_2299; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2301 = 8'h4d == total_offset_11 ? phv_data_77 : _GEN_2300; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2302 = 8'h4e == total_offset_11 ? phv_data_78 : _GEN_2301; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2303 = 8'h4f == total_offset_11 ? phv_data_79 : _GEN_2302; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2304 = 8'h50 == total_offset_11 ? phv_data_80 : _GEN_2303; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2305 = 8'h51 == total_offset_11 ? phv_data_81 : _GEN_2304; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2306 = 8'h52 == total_offset_11 ? phv_data_82 : _GEN_2305; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2307 = 8'h53 == total_offset_11 ? phv_data_83 : _GEN_2306; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2308 = 8'h54 == total_offset_11 ? phv_data_84 : _GEN_2307; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2309 = 8'h55 == total_offset_11 ? phv_data_85 : _GEN_2308; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2310 = 8'h56 == total_offset_11 ? phv_data_86 : _GEN_2309; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2311 = 8'h57 == total_offset_11 ? phv_data_87 : _GEN_2310; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2312 = 8'h58 == total_offset_11 ? phv_data_88 : _GEN_2311; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2313 = 8'h59 == total_offset_11 ? phv_data_89 : _GEN_2312; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2314 = 8'h5a == total_offset_11 ? phv_data_90 : _GEN_2313; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2315 = 8'h5b == total_offset_11 ? phv_data_91 : _GEN_2314; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2316 = 8'h5c == total_offset_11 ? phv_data_92 : _GEN_2315; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2317 = 8'h5d == total_offset_11 ? phv_data_93 : _GEN_2316; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2318 = 8'h5e == total_offset_11 ? phv_data_94 : _GEN_2317; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2319 = 8'h5f == total_offset_11 ? phv_data_95 : _GEN_2318; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2320 = 8'h60 == total_offset_11 ? phv_data_96 : _GEN_2319; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2321 = 8'h61 == total_offset_11 ? phv_data_97 : _GEN_2320; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2322 = 8'h62 == total_offset_11 ? phv_data_98 : _GEN_2321; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2323 = 8'h63 == total_offset_11 ? phv_data_99 : _GEN_2322; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2324 = 8'h64 == total_offset_11 ? phv_data_100 : _GEN_2323; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2325 = 8'h65 == total_offset_11 ? phv_data_101 : _GEN_2324; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2326 = 8'h66 == total_offset_11 ? phv_data_102 : _GEN_2325; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2327 = 8'h67 == total_offset_11 ? phv_data_103 : _GEN_2326; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2328 = 8'h68 == total_offset_11 ? phv_data_104 : _GEN_2327; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2329 = 8'h69 == total_offset_11 ? phv_data_105 : _GEN_2328; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2330 = 8'h6a == total_offset_11 ? phv_data_106 : _GEN_2329; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2331 = 8'h6b == total_offset_11 ? phv_data_107 : _GEN_2330; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2332 = 8'h6c == total_offset_11 ? phv_data_108 : _GEN_2331; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2333 = 8'h6d == total_offset_11 ? phv_data_109 : _GEN_2332; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2334 = 8'h6e == total_offset_11 ? phv_data_110 : _GEN_2333; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2335 = 8'h6f == total_offset_11 ? phv_data_111 : _GEN_2334; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2336 = 8'h70 == total_offset_11 ? phv_data_112 : _GEN_2335; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2337 = 8'h71 == total_offset_11 ? phv_data_113 : _GEN_2336; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2338 = 8'h72 == total_offset_11 ? phv_data_114 : _GEN_2337; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2339 = 8'h73 == total_offset_11 ? phv_data_115 : _GEN_2338; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2340 = 8'h74 == total_offset_11 ? phv_data_116 : _GEN_2339; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2341 = 8'h75 == total_offset_11 ? phv_data_117 : _GEN_2340; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2342 = 8'h76 == total_offset_11 ? phv_data_118 : _GEN_2341; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2343 = 8'h77 == total_offset_11 ? phv_data_119 : _GEN_2342; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2344 = 8'h78 == total_offset_11 ? phv_data_120 : _GEN_2343; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2345 = 8'h79 == total_offset_11 ? phv_data_121 : _GEN_2344; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2346 = 8'h7a == total_offset_11 ? phv_data_122 : _GEN_2345; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2347 = 8'h7b == total_offset_11 ? phv_data_123 : _GEN_2346; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2348 = 8'h7c == total_offset_11 ? phv_data_124 : _GEN_2347; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2349 = 8'h7d == total_offset_11 ? phv_data_125 : _GEN_2348; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2350 = 8'h7e == total_offset_11 ? phv_data_126 : _GEN_2349; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2351 = 8'h7f == total_offset_11 ? phv_data_127 : _GEN_2350; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2352 = 8'h80 == total_offset_11 ? phv_data_128 : _GEN_2351; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2353 = 8'h81 == total_offset_11 ? phv_data_129 : _GEN_2352; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2354 = 8'h82 == total_offset_11 ? phv_data_130 : _GEN_2353; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2355 = 8'h83 == total_offset_11 ? phv_data_131 : _GEN_2354; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2356 = 8'h84 == total_offset_11 ? phv_data_132 : _GEN_2355; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2357 = 8'h85 == total_offset_11 ? phv_data_133 : _GEN_2356; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2358 = 8'h86 == total_offset_11 ? phv_data_134 : _GEN_2357; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2359 = 8'h87 == total_offset_11 ? phv_data_135 : _GEN_2358; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2360 = 8'h88 == total_offset_11 ? phv_data_136 : _GEN_2359; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2361 = 8'h89 == total_offset_11 ? phv_data_137 : _GEN_2360; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2362 = 8'h8a == total_offset_11 ? phv_data_138 : _GEN_2361; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2363 = 8'h8b == total_offset_11 ? phv_data_139 : _GEN_2362; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2364 = 8'h8c == total_offset_11 ? phv_data_140 : _GEN_2363; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2365 = 8'h8d == total_offset_11 ? phv_data_141 : _GEN_2364; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2366 = 8'h8e == total_offset_11 ? phv_data_142 : _GEN_2365; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2367 = 8'h8f == total_offset_11 ? phv_data_143 : _GEN_2366; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2368 = 8'h90 == total_offset_11 ? phv_data_144 : _GEN_2367; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2369 = 8'h91 == total_offset_11 ? phv_data_145 : _GEN_2368; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2370 = 8'h92 == total_offset_11 ? phv_data_146 : _GEN_2369; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2371 = 8'h93 == total_offset_11 ? phv_data_147 : _GEN_2370; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2372 = 8'h94 == total_offset_11 ? phv_data_148 : _GEN_2371; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2373 = 8'h95 == total_offset_11 ? phv_data_149 : _GEN_2372; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2374 = 8'h96 == total_offset_11 ? phv_data_150 : _GEN_2373; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2375 = 8'h97 == total_offset_11 ? phv_data_151 : _GEN_2374; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2376 = 8'h98 == total_offset_11 ? phv_data_152 : _GEN_2375; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2377 = 8'h99 == total_offset_11 ? phv_data_153 : _GEN_2376; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2378 = 8'h9a == total_offset_11 ? phv_data_154 : _GEN_2377; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2379 = 8'h9b == total_offset_11 ? phv_data_155 : _GEN_2378; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2380 = 8'h9c == total_offset_11 ? phv_data_156 : _GEN_2379; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2381 = 8'h9d == total_offset_11 ? phv_data_157 : _GEN_2380; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2382 = 8'h9e == total_offset_11 ? phv_data_158 : _GEN_2381; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes_2_0 = 8'h9f == total_offset_11 ? phv_data_159 : _GEN_2382; // @[executor.scala 197:66 executor.scala 197:66]
  wire [31:0] _io_field_out_2_T = {bytes_2_0,bytes_2_1,bytes_2_2,bytes_2_3}; // @[Cat.scala 30:58]
  wire [3:0] _io_mask_out_2_T = {_mask_3_T_17,mask_2_1,mask_2_2,mask_2_3}; // @[Cat.scala 30:58]
  wire [17:0] io_field_out_2_hi_4 = io_field_out_2_lo[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _io_field_out_2_T_4 = {io_field_out_2_hi_4,io_field_out_2_lo}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2609 = 4'hb == opcode_2 ? _io_field_out_2_T_4 : 32'h0; // @[executor.scala 230:56 executor.scala 231:41]
  wire [1:0] _GEN_2610 = from_header_2 ? bias_2 : 2'h0; // @[executor.scala 178:36 executor.scala 203:36 executor.scala 174:29]
  wire [31:0] _GEN_2611 = from_header_2 ? _io_field_out_2_T : _GEN_2609; // @[executor.scala 178:36 executor.scala 204:37]
  wire [3:0] _GEN_2612 = from_header_2 ? _io_mask_out_2_T : 4'h0; // @[executor.scala 178:36 executor.scala 205:37 executor.scala 173:29]
  wire [3:0] opcode_3 = vliw_3[31:28]; // @[primitive.scala 9:44]
  wire [13:0] io_field_out_3_lo = vliw_3[13:0]; // @[primitive.scala 11:44]
  wire  from_header_3 = length_3 != 8'h0; // @[executor.scala 177:45]
  wire [5:0] total_offset_hi_3 = offset_3[7:2]; // @[executor.scala 191:57]
  wire [7:0] _ending_T_7 = offset_3 + length_3; // @[executor.scala 193:46]
  wire [1:0] ending_3 = _ending_T_7[1:0]; // @[executor.scala 193:58]
  wire [3:0] _GEN_3509 = {{2'd0}, ending_3}; // @[executor.scala 194:45]
  wire [3:0] _bias_T_7 = 4'h4 - _GEN_3509; // @[executor.scala 194:45]
  wire [1:0] bias_3 = _bias_T_7[1:0]; // @[executor.scala 194:54]
  wire [7:0] total_offset_12 = {total_offset_hi_3,2'h0}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_2617 = 8'h1 == total_offset_12 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2618 = 8'h2 == total_offset_12 ? phv_data_2 : _GEN_2617; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2619 = 8'h3 == total_offset_12 ? phv_data_3 : _GEN_2618; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2620 = 8'h4 == total_offset_12 ? phv_data_4 : _GEN_2619; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2621 = 8'h5 == total_offset_12 ? phv_data_5 : _GEN_2620; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2622 = 8'h6 == total_offset_12 ? phv_data_6 : _GEN_2621; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2623 = 8'h7 == total_offset_12 ? phv_data_7 : _GEN_2622; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2624 = 8'h8 == total_offset_12 ? phv_data_8 : _GEN_2623; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2625 = 8'h9 == total_offset_12 ? phv_data_9 : _GEN_2624; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2626 = 8'ha == total_offset_12 ? phv_data_10 : _GEN_2625; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2627 = 8'hb == total_offset_12 ? phv_data_11 : _GEN_2626; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2628 = 8'hc == total_offset_12 ? phv_data_12 : _GEN_2627; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2629 = 8'hd == total_offset_12 ? phv_data_13 : _GEN_2628; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2630 = 8'he == total_offset_12 ? phv_data_14 : _GEN_2629; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2631 = 8'hf == total_offset_12 ? phv_data_15 : _GEN_2630; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2632 = 8'h10 == total_offset_12 ? phv_data_16 : _GEN_2631; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2633 = 8'h11 == total_offset_12 ? phv_data_17 : _GEN_2632; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2634 = 8'h12 == total_offset_12 ? phv_data_18 : _GEN_2633; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2635 = 8'h13 == total_offset_12 ? phv_data_19 : _GEN_2634; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2636 = 8'h14 == total_offset_12 ? phv_data_20 : _GEN_2635; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2637 = 8'h15 == total_offset_12 ? phv_data_21 : _GEN_2636; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2638 = 8'h16 == total_offset_12 ? phv_data_22 : _GEN_2637; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2639 = 8'h17 == total_offset_12 ? phv_data_23 : _GEN_2638; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2640 = 8'h18 == total_offset_12 ? phv_data_24 : _GEN_2639; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2641 = 8'h19 == total_offset_12 ? phv_data_25 : _GEN_2640; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2642 = 8'h1a == total_offset_12 ? phv_data_26 : _GEN_2641; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2643 = 8'h1b == total_offset_12 ? phv_data_27 : _GEN_2642; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2644 = 8'h1c == total_offset_12 ? phv_data_28 : _GEN_2643; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2645 = 8'h1d == total_offset_12 ? phv_data_29 : _GEN_2644; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2646 = 8'h1e == total_offset_12 ? phv_data_30 : _GEN_2645; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2647 = 8'h1f == total_offset_12 ? phv_data_31 : _GEN_2646; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2648 = 8'h20 == total_offset_12 ? phv_data_32 : _GEN_2647; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2649 = 8'h21 == total_offset_12 ? phv_data_33 : _GEN_2648; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2650 = 8'h22 == total_offset_12 ? phv_data_34 : _GEN_2649; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2651 = 8'h23 == total_offset_12 ? phv_data_35 : _GEN_2650; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2652 = 8'h24 == total_offset_12 ? phv_data_36 : _GEN_2651; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2653 = 8'h25 == total_offset_12 ? phv_data_37 : _GEN_2652; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2654 = 8'h26 == total_offset_12 ? phv_data_38 : _GEN_2653; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2655 = 8'h27 == total_offset_12 ? phv_data_39 : _GEN_2654; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2656 = 8'h28 == total_offset_12 ? phv_data_40 : _GEN_2655; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2657 = 8'h29 == total_offset_12 ? phv_data_41 : _GEN_2656; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2658 = 8'h2a == total_offset_12 ? phv_data_42 : _GEN_2657; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2659 = 8'h2b == total_offset_12 ? phv_data_43 : _GEN_2658; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2660 = 8'h2c == total_offset_12 ? phv_data_44 : _GEN_2659; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2661 = 8'h2d == total_offset_12 ? phv_data_45 : _GEN_2660; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2662 = 8'h2e == total_offset_12 ? phv_data_46 : _GEN_2661; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2663 = 8'h2f == total_offset_12 ? phv_data_47 : _GEN_2662; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2664 = 8'h30 == total_offset_12 ? phv_data_48 : _GEN_2663; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2665 = 8'h31 == total_offset_12 ? phv_data_49 : _GEN_2664; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2666 = 8'h32 == total_offset_12 ? phv_data_50 : _GEN_2665; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2667 = 8'h33 == total_offset_12 ? phv_data_51 : _GEN_2666; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2668 = 8'h34 == total_offset_12 ? phv_data_52 : _GEN_2667; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2669 = 8'h35 == total_offset_12 ? phv_data_53 : _GEN_2668; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2670 = 8'h36 == total_offset_12 ? phv_data_54 : _GEN_2669; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2671 = 8'h37 == total_offset_12 ? phv_data_55 : _GEN_2670; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2672 = 8'h38 == total_offset_12 ? phv_data_56 : _GEN_2671; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2673 = 8'h39 == total_offset_12 ? phv_data_57 : _GEN_2672; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2674 = 8'h3a == total_offset_12 ? phv_data_58 : _GEN_2673; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2675 = 8'h3b == total_offset_12 ? phv_data_59 : _GEN_2674; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2676 = 8'h3c == total_offset_12 ? phv_data_60 : _GEN_2675; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2677 = 8'h3d == total_offset_12 ? phv_data_61 : _GEN_2676; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2678 = 8'h3e == total_offset_12 ? phv_data_62 : _GEN_2677; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2679 = 8'h3f == total_offset_12 ? phv_data_63 : _GEN_2678; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2680 = 8'h40 == total_offset_12 ? phv_data_64 : _GEN_2679; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2681 = 8'h41 == total_offset_12 ? phv_data_65 : _GEN_2680; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2682 = 8'h42 == total_offset_12 ? phv_data_66 : _GEN_2681; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2683 = 8'h43 == total_offset_12 ? phv_data_67 : _GEN_2682; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2684 = 8'h44 == total_offset_12 ? phv_data_68 : _GEN_2683; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2685 = 8'h45 == total_offset_12 ? phv_data_69 : _GEN_2684; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2686 = 8'h46 == total_offset_12 ? phv_data_70 : _GEN_2685; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2687 = 8'h47 == total_offset_12 ? phv_data_71 : _GEN_2686; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2688 = 8'h48 == total_offset_12 ? phv_data_72 : _GEN_2687; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2689 = 8'h49 == total_offset_12 ? phv_data_73 : _GEN_2688; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2690 = 8'h4a == total_offset_12 ? phv_data_74 : _GEN_2689; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2691 = 8'h4b == total_offset_12 ? phv_data_75 : _GEN_2690; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2692 = 8'h4c == total_offset_12 ? phv_data_76 : _GEN_2691; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2693 = 8'h4d == total_offset_12 ? phv_data_77 : _GEN_2692; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2694 = 8'h4e == total_offset_12 ? phv_data_78 : _GEN_2693; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2695 = 8'h4f == total_offset_12 ? phv_data_79 : _GEN_2694; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2696 = 8'h50 == total_offset_12 ? phv_data_80 : _GEN_2695; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2697 = 8'h51 == total_offset_12 ? phv_data_81 : _GEN_2696; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2698 = 8'h52 == total_offset_12 ? phv_data_82 : _GEN_2697; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2699 = 8'h53 == total_offset_12 ? phv_data_83 : _GEN_2698; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2700 = 8'h54 == total_offset_12 ? phv_data_84 : _GEN_2699; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2701 = 8'h55 == total_offset_12 ? phv_data_85 : _GEN_2700; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2702 = 8'h56 == total_offset_12 ? phv_data_86 : _GEN_2701; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2703 = 8'h57 == total_offset_12 ? phv_data_87 : _GEN_2702; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2704 = 8'h58 == total_offset_12 ? phv_data_88 : _GEN_2703; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2705 = 8'h59 == total_offset_12 ? phv_data_89 : _GEN_2704; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2706 = 8'h5a == total_offset_12 ? phv_data_90 : _GEN_2705; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2707 = 8'h5b == total_offset_12 ? phv_data_91 : _GEN_2706; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2708 = 8'h5c == total_offset_12 ? phv_data_92 : _GEN_2707; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2709 = 8'h5d == total_offset_12 ? phv_data_93 : _GEN_2708; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2710 = 8'h5e == total_offset_12 ? phv_data_94 : _GEN_2709; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2711 = 8'h5f == total_offset_12 ? phv_data_95 : _GEN_2710; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2712 = 8'h60 == total_offset_12 ? phv_data_96 : _GEN_2711; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2713 = 8'h61 == total_offset_12 ? phv_data_97 : _GEN_2712; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2714 = 8'h62 == total_offset_12 ? phv_data_98 : _GEN_2713; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2715 = 8'h63 == total_offset_12 ? phv_data_99 : _GEN_2714; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2716 = 8'h64 == total_offset_12 ? phv_data_100 : _GEN_2715; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2717 = 8'h65 == total_offset_12 ? phv_data_101 : _GEN_2716; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2718 = 8'h66 == total_offset_12 ? phv_data_102 : _GEN_2717; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2719 = 8'h67 == total_offset_12 ? phv_data_103 : _GEN_2718; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2720 = 8'h68 == total_offset_12 ? phv_data_104 : _GEN_2719; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2721 = 8'h69 == total_offset_12 ? phv_data_105 : _GEN_2720; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2722 = 8'h6a == total_offset_12 ? phv_data_106 : _GEN_2721; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2723 = 8'h6b == total_offset_12 ? phv_data_107 : _GEN_2722; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2724 = 8'h6c == total_offset_12 ? phv_data_108 : _GEN_2723; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2725 = 8'h6d == total_offset_12 ? phv_data_109 : _GEN_2724; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2726 = 8'h6e == total_offset_12 ? phv_data_110 : _GEN_2725; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2727 = 8'h6f == total_offset_12 ? phv_data_111 : _GEN_2726; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2728 = 8'h70 == total_offset_12 ? phv_data_112 : _GEN_2727; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2729 = 8'h71 == total_offset_12 ? phv_data_113 : _GEN_2728; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2730 = 8'h72 == total_offset_12 ? phv_data_114 : _GEN_2729; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2731 = 8'h73 == total_offset_12 ? phv_data_115 : _GEN_2730; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2732 = 8'h74 == total_offset_12 ? phv_data_116 : _GEN_2731; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2733 = 8'h75 == total_offset_12 ? phv_data_117 : _GEN_2732; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2734 = 8'h76 == total_offset_12 ? phv_data_118 : _GEN_2733; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2735 = 8'h77 == total_offset_12 ? phv_data_119 : _GEN_2734; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2736 = 8'h78 == total_offset_12 ? phv_data_120 : _GEN_2735; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2737 = 8'h79 == total_offset_12 ? phv_data_121 : _GEN_2736; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2738 = 8'h7a == total_offset_12 ? phv_data_122 : _GEN_2737; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2739 = 8'h7b == total_offset_12 ? phv_data_123 : _GEN_2738; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2740 = 8'h7c == total_offset_12 ? phv_data_124 : _GEN_2739; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2741 = 8'h7d == total_offset_12 ? phv_data_125 : _GEN_2740; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2742 = 8'h7e == total_offset_12 ? phv_data_126 : _GEN_2741; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2743 = 8'h7f == total_offset_12 ? phv_data_127 : _GEN_2742; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2744 = 8'h80 == total_offset_12 ? phv_data_128 : _GEN_2743; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2745 = 8'h81 == total_offset_12 ? phv_data_129 : _GEN_2744; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2746 = 8'h82 == total_offset_12 ? phv_data_130 : _GEN_2745; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2747 = 8'h83 == total_offset_12 ? phv_data_131 : _GEN_2746; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2748 = 8'h84 == total_offset_12 ? phv_data_132 : _GEN_2747; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2749 = 8'h85 == total_offset_12 ? phv_data_133 : _GEN_2748; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2750 = 8'h86 == total_offset_12 ? phv_data_134 : _GEN_2749; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2751 = 8'h87 == total_offset_12 ? phv_data_135 : _GEN_2750; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2752 = 8'h88 == total_offset_12 ? phv_data_136 : _GEN_2751; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2753 = 8'h89 == total_offset_12 ? phv_data_137 : _GEN_2752; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2754 = 8'h8a == total_offset_12 ? phv_data_138 : _GEN_2753; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2755 = 8'h8b == total_offset_12 ? phv_data_139 : _GEN_2754; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2756 = 8'h8c == total_offset_12 ? phv_data_140 : _GEN_2755; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2757 = 8'h8d == total_offset_12 ? phv_data_141 : _GEN_2756; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2758 = 8'h8e == total_offset_12 ? phv_data_142 : _GEN_2757; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2759 = 8'h8f == total_offset_12 ? phv_data_143 : _GEN_2758; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2760 = 8'h90 == total_offset_12 ? phv_data_144 : _GEN_2759; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2761 = 8'h91 == total_offset_12 ? phv_data_145 : _GEN_2760; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2762 = 8'h92 == total_offset_12 ? phv_data_146 : _GEN_2761; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2763 = 8'h93 == total_offset_12 ? phv_data_147 : _GEN_2762; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2764 = 8'h94 == total_offset_12 ? phv_data_148 : _GEN_2763; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2765 = 8'h95 == total_offset_12 ? phv_data_149 : _GEN_2764; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2766 = 8'h96 == total_offset_12 ? phv_data_150 : _GEN_2765; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2767 = 8'h97 == total_offset_12 ? phv_data_151 : _GEN_2766; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2768 = 8'h98 == total_offset_12 ? phv_data_152 : _GEN_2767; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2769 = 8'h99 == total_offset_12 ? phv_data_153 : _GEN_2768; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2770 = 8'h9a == total_offset_12 ? phv_data_154 : _GEN_2769; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2771 = 8'h9b == total_offset_12 ? phv_data_155 : _GEN_2770; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2772 = 8'h9c == total_offset_12 ? phv_data_156 : _GEN_2771; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2773 = 8'h9d == total_offset_12 ? phv_data_157 : _GEN_2772; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2774 = 8'h9e == total_offset_12 ? phv_data_158 : _GEN_2773; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes_3_3 = 8'h9f == total_offset_12 ? phv_data_159 : _GEN_2774; // @[executor.scala 197:66 executor.scala 197:66]
  wire  _mask_3_T_24 = ending_3 == 2'h0; // @[executor.scala 199:88]
  wire  mask_3_3 = 2'h0 >= offset_3[1:0] & (2'h0 < ending_3 | ending_3 == 2'h0); // @[executor.scala 199:56]
  wire [7:0] total_offset_13 = {total_offset_hi_3,2'h1}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_2777 = 8'h1 == total_offset_13 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2778 = 8'h2 == total_offset_13 ? phv_data_2 : _GEN_2777; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2779 = 8'h3 == total_offset_13 ? phv_data_3 : _GEN_2778; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2780 = 8'h4 == total_offset_13 ? phv_data_4 : _GEN_2779; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2781 = 8'h5 == total_offset_13 ? phv_data_5 : _GEN_2780; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2782 = 8'h6 == total_offset_13 ? phv_data_6 : _GEN_2781; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2783 = 8'h7 == total_offset_13 ? phv_data_7 : _GEN_2782; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2784 = 8'h8 == total_offset_13 ? phv_data_8 : _GEN_2783; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2785 = 8'h9 == total_offset_13 ? phv_data_9 : _GEN_2784; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2786 = 8'ha == total_offset_13 ? phv_data_10 : _GEN_2785; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2787 = 8'hb == total_offset_13 ? phv_data_11 : _GEN_2786; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2788 = 8'hc == total_offset_13 ? phv_data_12 : _GEN_2787; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2789 = 8'hd == total_offset_13 ? phv_data_13 : _GEN_2788; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2790 = 8'he == total_offset_13 ? phv_data_14 : _GEN_2789; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2791 = 8'hf == total_offset_13 ? phv_data_15 : _GEN_2790; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2792 = 8'h10 == total_offset_13 ? phv_data_16 : _GEN_2791; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2793 = 8'h11 == total_offset_13 ? phv_data_17 : _GEN_2792; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2794 = 8'h12 == total_offset_13 ? phv_data_18 : _GEN_2793; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2795 = 8'h13 == total_offset_13 ? phv_data_19 : _GEN_2794; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2796 = 8'h14 == total_offset_13 ? phv_data_20 : _GEN_2795; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2797 = 8'h15 == total_offset_13 ? phv_data_21 : _GEN_2796; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2798 = 8'h16 == total_offset_13 ? phv_data_22 : _GEN_2797; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2799 = 8'h17 == total_offset_13 ? phv_data_23 : _GEN_2798; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2800 = 8'h18 == total_offset_13 ? phv_data_24 : _GEN_2799; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2801 = 8'h19 == total_offset_13 ? phv_data_25 : _GEN_2800; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2802 = 8'h1a == total_offset_13 ? phv_data_26 : _GEN_2801; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2803 = 8'h1b == total_offset_13 ? phv_data_27 : _GEN_2802; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2804 = 8'h1c == total_offset_13 ? phv_data_28 : _GEN_2803; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2805 = 8'h1d == total_offset_13 ? phv_data_29 : _GEN_2804; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2806 = 8'h1e == total_offset_13 ? phv_data_30 : _GEN_2805; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2807 = 8'h1f == total_offset_13 ? phv_data_31 : _GEN_2806; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2808 = 8'h20 == total_offset_13 ? phv_data_32 : _GEN_2807; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2809 = 8'h21 == total_offset_13 ? phv_data_33 : _GEN_2808; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2810 = 8'h22 == total_offset_13 ? phv_data_34 : _GEN_2809; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2811 = 8'h23 == total_offset_13 ? phv_data_35 : _GEN_2810; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2812 = 8'h24 == total_offset_13 ? phv_data_36 : _GEN_2811; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2813 = 8'h25 == total_offset_13 ? phv_data_37 : _GEN_2812; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2814 = 8'h26 == total_offset_13 ? phv_data_38 : _GEN_2813; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2815 = 8'h27 == total_offset_13 ? phv_data_39 : _GEN_2814; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2816 = 8'h28 == total_offset_13 ? phv_data_40 : _GEN_2815; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2817 = 8'h29 == total_offset_13 ? phv_data_41 : _GEN_2816; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2818 = 8'h2a == total_offset_13 ? phv_data_42 : _GEN_2817; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2819 = 8'h2b == total_offset_13 ? phv_data_43 : _GEN_2818; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2820 = 8'h2c == total_offset_13 ? phv_data_44 : _GEN_2819; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2821 = 8'h2d == total_offset_13 ? phv_data_45 : _GEN_2820; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2822 = 8'h2e == total_offset_13 ? phv_data_46 : _GEN_2821; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2823 = 8'h2f == total_offset_13 ? phv_data_47 : _GEN_2822; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2824 = 8'h30 == total_offset_13 ? phv_data_48 : _GEN_2823; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2825 = 8'h31 == total_offset_13 ? phv_data_49 : _GEN_2824; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2826 = 8'h32 == total_offset_13 ? phv_data_50 : _GEN_2825; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2827 = 8'h33 == total_offset_13 ? phv_data_51 : _GEN_2826; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2828 = 8'h34 == total_offset_13 ? phv_data_52 : _GEN_2827; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2829 = 8'h35 == total_offset_13 ? phv_data_53 : _GEN_2828; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2830 = 8'h36 == total_offset_13 ? phv_data_54 : _GEN_2829; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2831 = 8'h37 == total_offset_13 ? phv_data_55 : _GEN_2830; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2832 = 8'h38 == total_offset_13 ? phv_data_56 : _GEN_2831; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2833 = 8'h39 == total_offset_13 ? phv_data_57 : _GEN_2832; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2834 = 8'h3a == total_offset_13 ? phv_data_58 : _GEN_2833; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2835 = 8'h3b == total_offset_13 ? phv_data_59 : _GEN_2834; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2836 = 8'h3c == total_offset_13 ? phv_data_60 : _GEN_2835; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2837 = 8'h3d == total_offset_13 ? phv_data_61 : _GEN_2836; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2838 = 8'h3e == total_offset_13 ? phv_data_62 : _GEN_2837; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2839 = 8'h3f == total_offset_13 ? phv_data_63 : _GEN_2838; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2840 = 8'h40 == total_offset_13 ? phv_data_64 : _GEN_2839; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2841 = 8'h41 == total_offset_13 ? phv_data_65 : _GEN_2840; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2842 = 8'h42 == total_offset_13 ? phv_data_66 : _GEN_2841; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2843 = 8'h43 == total_offset_13 ? phv_data_67 : _GEN_2842; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2844 = 8'h44 == total_offset_13 ? phv_data_68 : _GEN_2843; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2845 = 8'h45 == total_offset_13 ? phv_data_69 : _GEN_2844; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2846 = 8'h46 == total_offset_13 ? phv_data_70 : _GEN_2845; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2847 = 8'h47 == total_offset_13 ? phv_data_71 : _GEN_2846; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2848 = 8'h48 == total_offset_13 ? phv_data_72 : _GEN_2847; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2849 = 8'h49 == total_offset_13 ? phv_data_73 : _GEN_2848; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2850 = 8'h4a == total_offset_13 ? phv_data_74 : _GEN_2849; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2851 = 8'h4b == total_offset_13 ? phv_data_75 : _GEN_2850; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2852 = 8'h4c == total_offset_13 ? phv_data_76 : _GEN_2851; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2853 = 8'h4d == total_offset_13 ? phv_data_77 : _GEN_2852; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2854 = 8'h4e == total_offset_13 ? phv_data_78 : _GEN_2853; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2855 = 8'h4f == total_offset_13 ? phv_data_79 : _GEN_2854; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2856 = 8'h50 == total_offset_13 ? phv_data_80 : _GEN_2855; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2857 = 8'h51 == total_offset_13 ? phv_data_81 : _GEN_2856; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2858 = 8'h52 == total_offset_13 ? phv_data_82 : _GEN_2857; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2859 = 8'h53 == total_offset_13 ? phv_data_83 : _GEN_2858; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2860 = 8'h54 == total_offset_13 ? phv_data_84 : _GEN_2859; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2861 = 8'h55 == total_offset_13 ? phv_data_85 : _GEN_2860; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2862 = 8'h56 == total_offset_13 ? phv_data_86 : _GEN_2861; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2863 = 8'h57 == total_offset_13 ? phv_data_87 : _GEN_2862; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2864 = 8'h58 == total_offset_13 ? phv_data_88 : _GEN_2863; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2865 = 8'h59 == total_offset_13 ? phv_data_89 : _GEN_2864; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2866 = 8'h5a == total_offset_13 ? phv_data_90 : _GEN_2865; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2867 = 8'h5b == total_offset_13 ? phv_data_91 : _GEN_2866; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2868 = 8'h5c == total_offset_13 ? phv_data_92 : _GEN_2867; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2869 = 8'h5d == total_offset_13 ? phv_data_93 : _GEN_2868; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2870 = 8'h5e == total_offset_13 ? phv_data_94 : _GEN_2869; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2871 = 8'h5f == total_offset_13 ? phv_data_95 : _GEN_2870; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2872 = 8'h60 == total_offset_13 ? phv_data_96 : _GEN_2871; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2873 = 8'h61 == total_offset_13 ? phv_data_97 : _GEN_2872; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2874 = 8'h62 == total_offset_13 ? phv_data_98 : _GEN_2873; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2875 = 8'h63 == total_offset_13 ? phv_data_99 : _GEN_2874; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2876 = 8'h64 == total_offset_13 ? phv_data_100 : _GEN_2875; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2877 = 8'h65 == total_offset_13 ? phv_data_101 : _GEN_2876; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2878 = 8'h66 == total_offset_13 ? phv_data_102 : _GEN_2877; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2879 = 8'h67 == total_offset_13 ? phv_data_103 : _GEN_2878; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2880 = 8'h68 == total_offset_13 ? phv_data_104 : _GEN_2879; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2881 = 8'h69 == total_offset_13 ? phv_data_105 : _GEN_2880; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2882 = 8'h6a == total_offset_13 ? phv_data_106 : _GEN_2881; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2883 = 8'h6b == total_offset_13 ? phv_data_107 : _GEN_2882; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2884 = 8'h6c == total_offset_13 ? phv_data_108 : _GEN_2883; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2885 = 8'h6d == total_offset_13 ? phv_data_109 : _GEN_2884; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2886 = 8'h6e == total_offset_13 ? phv_data_110 : _GEN_2885; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2887 = 8'h6f == total_offset_13 ? phv_data_111 : _GEN_2886; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2888 = 8'h70 == total_offset_13 ? phv_data_112 : _GEN_2887; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2889 = 8'h71 == total_offset_13 ? phv_data_113 : _GEN_2888; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2890 = 8'h72 == total_offset_13 ? phv_data_114 : _GEN_2889; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2891 = 8'h73 == total_offset_13 ? phv_data_115 : _GEN_2890; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2892 = 8'h74 == total_offset_13 ? phv_data_116 : _GEN_2891; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2893 = 8'h75 == total_offset_13 ? phv_data_117 : _GEN_2892; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2894 = 8'h76 == total_offset_13 ? phv_data_118 : _GEN_2893; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2895 = 8'h77 == total_offset_13 ? phv_data_119 : _GEN_2894; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2896 = 8'h78 == total_offset_13 ? phv_data_120 : _GEN_2895; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2897 = 8'h79 == total_offset_13 ? phv_data_121 : _GEN_2896; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2898 = 8'h7a == total_offset_13 ? phv_data_122 : _GEN_2897; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2899 = 8'h7b == total_offset_13 ? phv_data_123 : _GEN_2898; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2900 = 8'h7c == total_offset_13 ? phv_data_124 : _GEN_2899; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2901 = 8'h7d == total_offset_13 ? phv_data_125 : _GEN_2900; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2902 = 8'h7e == total_offset_13 ? phv_data_126 : _GEN_2901; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2903 = 8'h7f == total_offset_13 ? phv_data_127 : _GEN_2902; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2904 = 8'h80 == total_offset_13 ? phv_data_128 : _GEN_2903; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2905 = 8'h81 == total_offset_13 ? phv_data_129 : _GEN_2904; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2906 = 8'h82 == total_offset_13 ? phv_data_130 : _GEN_2905; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2907 = 8'h83 == total_offset_13 ? phv_data_131 : _GEN_2906; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2908 = 8'h84 == total_offset_13 ? phv_data_132 : _GEN_2907; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2909 = 8'h85 == total_offset_13 ? phv_data_133 : _GEN_2908; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2910 = 8'h86 == total_offset_13 ? phv_data_134 : _GEN_2909; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2911 = 8'h87 == total_offset_13 ? phv_data_135 : _GEN_2910; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2912 = 8'h88 == total_offset_13 ? phv_data_136 : _GEN_2911; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2913 = 8'h89 == total_offset_13 ? phv_data_137 : _GEN_2912; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2914 = 8'h8a == total_offset_13 ? phv_data_138 : _GEN_2913; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2915 = 8'h8b == total_offset_13 ? phv_data_139 : _GEN_2914; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2916 = 8'h8c == total_offset_13 ? phv_data_140 : _GEN_2915; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2917 = 8'h8d == total_offset_13 ? phv_data_141 : _GEN_2916; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2918 = 8'h8e == total_offset_13 ? phv_data_142 : _GEN_2917; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2919 = 8'h8f == total_offset_13 ? phv_data_143 : _GEN_2918; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2920 = 8'h90 == total_offset_13 ? phv_data_144 : _GEN_2919; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2921 = 8'h91 == total_offset_13 ? phv_data_145 : _GEN_2920; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2922 = 8'h92 == total_offset_13 ? phv_data_146 : _GEN_2921; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2923 = 8'h93 == total_offset_13 ? phv_data_147 : _GEN_2922; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2924 = 8'h94 == total_offset_13 ? phv_data_148 : _GEN_2923; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2925 = 8'h95 == total_offset_13 ? phv_data_149 : _GEN_2924; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2926 = 8'h96 == total_offset_13 ? phv_data_150 : _GEN_2925; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2927 = 8'h97 == total_offset_13 ? phv_data_151 : _GEN_2926; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2928 = 8'h98 == total_offset_13 ? phv_data_152 : _GEN_2927; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2929 = 8'h99 == total_offset_13 ? phv_data_153 : _GEN_2928; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2930 = 8'h9a == total_offset_13 ? phv_data_154 : _GEN_2929; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2931 = 8'h9b == total_offset_13 ? phv_data_155 : _GEN_2930; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2932 = 8'h9c == total_offset_13 ? phv_data_156 : _GEN_2931; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2933 = 8'h9d == total_offset_13 ? phv_data_157 : _GEN_2932; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2934 = 8'h9e == total_offset_13 ? phv_data_158 : _GEN_2933; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes_3_2 = 8'h9f == total_offset_13 ? phv_data_159 : _GEN_2934; // @[executor.scala 197:66 executor.scala 197:66]
  wire  mask_3_2 = 2'h1 >= offset_3[1:0] & (2'h1 < ending_3 | ending_3 == 2'h0); // @[executor.scala 199:56]
  wire [7:0] total_offset_14 = {total_offset_hi_3,2'h2}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_2937 = 8'h1 == total_offset_14 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2938 = 8'h2 == total_offset_14 ? phv_data_2 : _GEN_2937; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2939 = 8'h3 == total_offset_14 ? phv_data_3 : _GEN_2938; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2940 = 8'h4 == total_offset_14 ? phv_data_4 : _GEN_2939; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2941 = 8'h5 == total_offset_14 ? phv_data_5 : _GEN_2940; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2942 = 8'h6 == total_offset_14 ? phv_data_6 : _GEN_2941; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2943 = 8'h7 == total_offset_14 ? phv_data_7 : _GEN_2942; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2944 = 8'h8 == total_offset_14 ? phv_data_8 : _GEN_2943; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2945 = 8'h9 == total_offset_14 ? phv_data_9 : _GEN_2944; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2946 = 8'ha == total_offset_14 ? phv_data_10 : _GEN_2945; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2947 = 8'hb == total_offset_14 ? phv_data_11 : _GEN_2946; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2948 = 8'hc == total_offset_14 ? phv_data_12 : _GEN_2947; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2949 = 8'hd == total_offset_14 ? phv_data_13 : _GEN_2948; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2950 = 8'he == total_offset_14 ? phv_data_14 : _GEN_2949; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2951 = 8'hf == total_offset_14 ? phv_data_15 : _GEN_2950; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2952 = 8'h10 == total_offset_14 ? phv_data_16 : _GEN_2951; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2953 = 8'h11 == total_offset_14 ? phv_data_17 : _GEN_2952; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2954 = 8'h12 == total_offset_14 ? phv_data_18 : _GEN_2953; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2955 = 8'h13 == total_offset_14 ? phv_data_19 : _GEN_2954; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2956 = 8'h14 == total_offset_14 ? phv_data_20 : _GEN_2955; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2957 = 8'h15 == total_offset_14 ? phv_data_21 : _GEN_2956; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2958 = 8'h16 == total_offset_14 ? phv_data_22 : _GEN_2957; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2959 = 8'h17 == total_offset_14 ? phv_data_23 : _GEN_2958; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2960 = 8'h18 == total_offset_14 ? phv_data_24 : _GEN_2959; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2961 = 8'h19 == total_offset_14 ? phv_data_25 : _GEN_2960; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2962 = 8'h1a == total_offset_14 ? phv_data_26 : _GEN_2961; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2963 = 8'h1b == total_offset_14 ? phv_data_27 : _GEN_2962; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2964 = 8'h1c == total_offset_14 ? phv_data_28 : _GEN_2963; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2965 = 8'h1d == total_offset_14 ? phv_data_29 : _GEN_2964; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2966 = 8'h1e == total_offset_14 ? phv_data_30 : _GEN_2965; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2967 = 8'h1f == total_offset_14 ? phv_data_31 : _GEN_2966; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2968 = 8'h20 == total_offset_14 ? phv_data_32 : _GEN_2967; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2969 = 8'h21 == total_offset_14 ? phv_data_33 : _GEN_2968; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2970 = 8'h22 == total_offset_14 ? phv_data_34 : _GEN_2969; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2971 = 8'h23 == total_offset_14 ? phv_data_35 : _GEN_2970; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2972 = 8'h24 == total_offset_14 ? phv_data_36 : _GEN_2971; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2973 = 8'h25 == total_offset_14 ? phv_data_37 : _GEN_2972; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2974 = 8'h26 == total_offset_14 ? phv_data_38 : _GEN_2973; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2975 = 8'h27 == total_offset_14 ? phv_data_39 : _GEN_2974; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2976 = 8'h28 == total_offset_14 ? phv_data_40 : _GEN_2975; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2977 = 8'h29 == total_offset_14 ? phv_data_41 : _GEN_2976; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2978 = 8'h2a == total_offset_14 ? phv_data_42 : _GEN_2977; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2979 = 8'h2b == total_offset_14 ? phv_data_43 : _GEN_2978; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2980 = 8'h2c == total_offset_14 ? phv_data_44 : _GEN_2979; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2981 = 8'h2d == total_offset_14 ? phv_data_45 : _GEN_2980; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2982 = 8'h2e == total_offset_14 ? phv_data_46 : _GEN_2981; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2983 = 8'h2f == total_offset_14 ? phv_data_47 : _GEN_2982; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2984 = 8'h30 == total_offset_14 ? phv_data_48 : _GEN_2983; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2985 = 8'h31 == total_offset_14 ? phv_data_49 : _GEN_2984; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2986 = 8'h32 == total_offset_14 ? phv_data_50 : _GEN_2985; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2987 = 8'h33 == total_offset_14 ? phv_data_51 : _GEN_2986; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2988 = 8'h34 == total_offset_14 ? phv_data_52 : _GEN_2987; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2989 = 8'h35 == total_offset_14 ? phv_data_53 : _GEN_2988; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2990 = 8'h36 == total_offset_14 ? phv_data_54 : _GEN_2989; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2991 = 8'h37 == total_offset_14 ? phv_data_55 : _GEN_2990; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2992 = 8'h38 == total_offset_14 ? phv_data_56 : _GEN_2991; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2993 = 8'h39 == total_offset_14 ? phv_data_57 : _GEN_2992; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2994 = 8'h3a == total_offset_14 ? phv_data_58 : _GEN_2993; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2995 = 8'h3b == total_offset_14 ? phv_data_59 : _GEN_2994; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2996 = 8'h3c == total_offset_14 ? phv_data_60 : _GEN_2995; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2997 = 8'h3d == total_offset_14 ? phv_data_61 : _GEN_2996; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2998 = 8'h3e == total_offset_14 ? phv_data_62 : _GEN_2997; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2999 = 8'h3f == total_offset_14 ? phv_data_63 : _GEN_2998; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3000 = 8'h40 == total_offset_14 ? phv_data_64 : _GEN_2999; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3001 = 8'h41 == total_offset_14 ? phv_data_65 : _GEN_3000; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3002 = 8'h42 == total_offset_14 ? phv_data_66 : _GEN_3001; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3003 = 8'h43 == total_offset_14 ? phv_data_67 : _GEN_3002; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3004 = 8'h44 == total_offset_14 ? phv_data_68 : _GEN_3003; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3005 = 8'h45 == total_offset_14 ? phv_data_69 : _GEN_3004; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3006 = 8'h46 == total_offset_14 ? phv_data_70 : _GEN_3005; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3007 = 8'h47 == total_offset_14 ? phv_data_71 : _GEN_3006; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3008 = 8'h48 == total_offset_14 ? phv_data_72 : _GEN_3007; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3009 = 8'h49 == total_offset_14 ? phv_data_73 : _GEN_3008; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3010 = 8'h4a == total_offset_14 ? phv_data_74 : _GEN_3009; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3011 = 8'h4b == total_offset_14 ? phv_data_75 : _GEN_3010; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3012 = 8'h4c == total_offset_14 ? phv_data_76 : _GEN_3011; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3013 = 8'h4d == total_offset_14 ? phv_data_77 : _GEN_3012; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3014 = 8'h4e == total_offset_14 ? phv_data_78 : _GEN_3013; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3015 = 8'h4f == total_offset_14 ? phv_data_79 : _GEN_3014; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3016 = 8'h50 == total_offset_14 ? phv_data_80 : _GEN_3015; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3017 = 8'h51 == total_offset_14 ? phv_data_81 : _GEN_3016; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3018 = 8'h52 == total_offset_14 ? phv_data_82 : _GEN_3017; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3019 = 8'h53 == total_offset_14 ? phv_data_83 : _GEN_3018; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3020 = 8'h54 == total_offset_14 ? phv_data_84 : _GEN_3019; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3021 = 8'h55 == total_offset_14 ? phv_data_85 : _GEN_3020; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3022 = 8'h56 == total_offset_14 ? phv_data_86 : _GEN_3021; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3023 = 8'h57 == total_offset_14 ? phv_data_87 : _GEN_3022; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3024 = 8'h58 == total_offset_14 ? phv_data_88 : _GEN_3023; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3025 = 8'h59 == total_offset_14 ? phv_data_89 : _GEN_3024; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3026 = 8'h5a == total_offset_14 ? phv_data_90 : _GEN_3025; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3027 = 8'h5b == total_offset_14 ? phv_data_91 : _GEN_3026; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3028 = 8'h5c == total_offset_14 ? phv_data_92 : _GEN_3027; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3029 = 8'h5d == total_offset_14 ? phv_data_93 : _GEN_3028; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3030 = 8'h5e == total_offset_14 ? phv_data_94 : _GEN_3029; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3031 = 8'h5f == total_offset_14 ? phv_data_95 : _GEN_3030; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3032 = 8'h60 == total_offset_14 ? phv_data_96 : _GEN_3031; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3033 = 8'h61 == total_offset_14 ? phv_data_97 : _GEN_3032; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3034 = 8'h62 == total_offset_14 ? phv_data_98 : _GEN_3033; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3035 = 8'h63 == total_offset_14 ? phv_data_99 : _GEN_3034; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3036 = 8'h64 == total_offset_14 ? phv_data_100 : _GEN_3035; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3037 = 8'h65 == total_offset_14 ? phv_data_101 : _GEN_3036; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3038 = 8'h66 == total_offset_14 ? phv_data_102 : _GEN_3037; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3039 = 8'h67 == total_offset_14 ? phv_data_103 : _GEN_3038; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3040 = 8'h68 == total_offset_14 ? phv_data_104 : _GEN_3039; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3041 = 8'h69 == total_offset_14 ? phv_data_105 : _GEN_3040; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3042 = 8'h6a == total_offset_14 ? phv_data_106 : _GEN_3041; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3043 = 8'h6b == total_offset_14 ? phv_data_107 : _GEN_3042; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3044 = 8'h6c == total_offset_14 ? phv_data_108 : _GEN_3043; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3045 = 8'h6d == total_offset_14 ? phv_data_109 : _GEN_3044; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3046 = 8'h6e == total_offset_14 ? phv_data_110 : _GEN_3045; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3047 = 8'h6f == total_offset_14 ? phv_data_111 : _GEN_3046; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3048 = 8'h70 == total_offset_14 ? phv_data_112 : _GEN_3047; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3049 = 8'h71 == total_offset_14 ? phv_data_113 : _GEN_3048; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3050 = 8'h72 == total_offset_14 ? phv_data_114 : _GEN_3049; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3051 = 8'h73 == total_offset_14 ? phv_data_115 : _GEN_3050; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3052 = 8'h74 == total_offset_14 ? phv_data_116 : _GEN_3051; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3053 = 8'h75 == total_offset_14 ? phv_data_117 : _GEN_3052; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3054 = 8'h76 == total_offset_14 ? phv_data_118 : _GEN_3053; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3055 = 8'h77 == total_offset_14 ? phv_data_119 : _GEN_3054; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3056 = 8'h78 == total_offset_14 ? phv_data_120 : _GEN_3055; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3057 = 8'h79 == total_offset_14 ? phv_data_121 : _GEN_3056; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3058 = 8'h7a == total_offset_14 ? phv_data_122 : _GEN_3057; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3059 = 8'h7b == total_offset_14 ? phv_data_123 : _GEN_3058; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3060 = 8'h7c == total_offset_14 ? phv_data_124 : _GEN_3059; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3061 = 8'h7d == total_offset_14 ? phv_data_125 : _GEN_3060; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3062 = 8'h7e == total_offset_14 ? phv_data_126 : _GEN_3061; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3063 = 8'h7f == total_offset_14 ? phv_data_127 : _GEN_3062; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3064 = 8'h80 == total_offset_14 ? phv_data_128 : _GEN_3063; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3065 = 8'h81 == total_offset_14 ? phv_data_129 : _GEN_3064; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3066 = 8'h82 == total_offset_14 ? phv_data_130 : _GEN_3065; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3067 = 8'h83 == total_offset_14 ? phv_data_131 : _GEN_3066; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3068 = 8'h84 == total_offset_14 ? phv_data_132 : _GEN_3067; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3069 = 8'h85 == total_offset_14 ? phv_data_133 : _GEN_3068; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3070 = 8'h86 == total_offset_14 ? phv_data_134 : _GEN_3069; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3071 = 8'h87 == total_offset_14 ? phv_data_135 : _GEN_3070; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3072 = 8'h88 == total_offset_14 ? phv_data_136 : _GEN_3071; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3073 = 8'h89 == total_offset_14 ? phv_data_137 : _GEN_3072; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3074 = 8'h8a == total_offset_14 ? phv_data_138 : _GEN_3073; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3075 = 8'h8b == total_offset_14 ? phv_data_139 : _GEN_3074; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3076 = 8'h8c == total_offset_14 ? phv_data_140 : _GEN_3075; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3077 = 8'h8d == total_offset_14 ? phv_data_141 : _GEN_3076; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3078 = 8'h8e == total_offset_14 ? phv_data_142 : _GEN_3077; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3079 = 8'h8f == total_offset_14 ? phv_data_143 : _GEN_3078; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3080 = 8'h90 == total_offset_14 ? phv_data_144 : _GEN_3079; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3081 = 8'h91 == total_offset_14 ? phv_data_145 : _GEN_3080; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3082 = 8'h92 == total_offset_14 ? phv_data_146 : _GEN_3081; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3083 = 8'h93 == total_offset_14 ? phv_data_147 : _GEN_3082; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3084 = 8'h94 == total_offset_14 ? phv_data_148 : _GEN_3083; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3085 = 8'h95 == total_offset_14 ? phv_data_149 : _GEN_3084; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3086 = 8'h96 == total_offset_14 ? phv_data_150 : _GEN_3085; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3087 = 8'h97 == total_offset_14 ? phv_data_151 : _GEN_3086; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3088 = 8'h98 == total_offset_14 ? phv_data_152 : _GEN_3087; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3089 = 8'h99 == total_offset_14 ? phv_data_153 : _GEN_3088; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3090 = 8'h9a == total_offset_14 ? phv_data_154 : _GEN_3089; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3091 = 8'h9b == total_offset_14 ? phv_data_155 : _GEN_3090; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3092 = 8'h9c == total_offset_14 ? phv_data_156 : _GEN_3091; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3093 = 8'h9d == total_offset_14 ? phv_data_157 : _GEN_3092; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3094 = 8'h9e == total_offset_14 ? phv_data_158 : _GEN_3093; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes_3_1 = 8'h9f == total_offset_14 ? phv_data_159 : _GEN_3094; // @[executor.scala 197:66 executor.scala 197:66]
  wire  mask_3_1 = 2'h2 >= offset_3[1:0] & (2'h2 < ending_3 | ending_3 == 2'h0); // @[executor.scala 199:56]
  wire [7:0] total_offset_15 = {total_offset_hi_3,2'h3}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_3097 = 8'h1 == total_offset_15 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3098 = 8'h2 == total_offset_15 ? phv_data_2 : _GEN_3097; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3099 = 8'h3 == total_offset_15 ? phv_data_3 : _GEN_3098; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3100 = 8'h4 == total_offset_15 ? phv_data_4 : _GEN_3099; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3101 = 8'h5 == total_offset_15 ? phv_data_5 : _GEN_3100; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3102 = 8'h6 == total_offset_15 ? phv_data_6 : _GEN_3101; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3103 = 8'h7 == total_offset_15 ? phv_data_7 : _GEN_3102; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3104 = 8'h8 == total_offset_15 ? phv_data_8 : _GEN_3103; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3105 = 8'h9 == total_offset_15 ? phv_data_9 : _GEN_3104; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3106 = 8'ha == total_offset_15 ? phv_data_10 : _GEN_3105; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3107 = 8'hb == total_offset_15 ? phv_data_11 : _GEN_3106; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3108 = 8'hc == total_offset_15 ? phv_data_12 : _GEN_3107; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3109 = 8'hd == total_offset_15 ? phv_data_13 : _GEN_3108; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3110 = 8'he == total_offset_15 ? phv_data_14 : _GEN_3109; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3111 = 8'hf == total_offset_15 ? phv_data_15 : _GEN_3110; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3112 = 8'h10 == total_offset_15 ? phv_data_16 : _GEN_3111; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3113 = 8'h11 == total_offset_15 ? phv_data_17 : _GEN_3112; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3114 = 8'h12 == total_offset_15 ? phv_data_18 : _GEN_3113; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3115 = 8'h13 == total_offset_15 ? phv_data_19 : _GEN_3114; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3116 = 8'h14 == total_offset_15 ? phv_data_20 : _GEN_3115; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3117 = 8'h15 == total_offset_15 ? phv_data_21 : _GEN_3116; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3118 = 8'h16 == total_offset_15 ? phv_data_22 : _GEN_3117; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3119 = 8'h17 == total_offset_15 ? phv_data_23 : _GEN_3118; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3120 = 8'h18 == total_offset_15 ? phv_data_24 : _GEN_3119; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3121 = 8'h19 == total_offset_15 ? phv_data_25 : _GEN_3120; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3122 = 8'h1a == total_offset_15 ? phv_data_26 : _GEN_3121; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3123 = 8'h1b == total_offset_15 ? phv_data_27 : _GEN_3122; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3124 = 8'h1c == total_offset_15 ? phv_data_28 : _GEN_3123; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3125 = 8'h1d == total_offset_15 ? phv_data_29 : _GEN_3124; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3126 = 8'h1e == total_offset_15 ? phv_data_30 : _GEN_3125; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3127 = 8'h1f == total_offset_15 ? phv_data_31 : _GEN_3126; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3128 = 8'h20 == total_offset_15 ? phv_data_32 : _GEN_3127; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3129 = 8'h21 == total_offset_15 ? phv_data_33 : _GEN_3128; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3130 = 8'h22 == total_offset_15 ? phv_data_34 : _GEN_3129; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3131 = 8'h23 == total_offset_15 ? phv_data_35 : _GEN_3130; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3132 = 8'h24 == total_offset_15 ? phv_data_36 : _GEN_3131; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3133 = 8'h25 == total_offset_15 ? phv_data_37 : _GEN_3132; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3134 = 8'h26 == total_offset_15 ? phv_data_38 : _GEN_3133; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3135 = 8'h27 == total_offset_15 ? phv_data_39 : _GEN_3134; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3136 = 8'h28 == total_offset_15 ? phv_data_40 : _GEN_3135; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3137 = 8'h29 == total_offset_15 ? phv_data_41 : _GEN_3136; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3138 = 8'h2a == total_offset_15 ? phv_data_42 : _GEN_3137; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3139 = 8'h2b == total_offset_15 ? phv_data_43 : _GEN_3138; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3140 = 8'h2c == total_offset_15 ? phv_data_44 : _GEN_3139; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3141 = 8'h2d == total_offset_15 ? phv_data_45 : _GEN_3140; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3142 = 8'h2e == total_offset_15 ? phv_data_46 : _GEN_3141; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3143 = 8'h2f == total_offset_15 ? phv_data_47 : _GEN_3142; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3144 = 8'h30 == total_offset_15 ? phv_data_48 : _GEN_3143; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3145 = 8'h31 == total_offset_15 ? phv_data_49 : _GEN_3144; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3146 = 8'h32 == total_offset_15 ? phv_data_50 : _GEN_3145; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3147 = 8'h33 == total_offset_15 ? phv_data_51 : _GEN_3146; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3148 = 8'h34 == total_offset_15 ? phv_data_52 : _GEN_3147; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3149 = 8'h35 == total_offset_15 ? phv_data_53 : _GEN_3148; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3150 = 8'h36 == total_offset_15 ? phv_data_54 : _GEN_3149; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3151 = 8'h37 == total_offset_15 ? phv_data_55 : _GEN_3150; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3152 = 8'h38 == total_offset_15 ? phv_data_56 : _GEN_3151; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3153 = 8'h39 == total_offset_15 ? phv_data_57 : _GEN_3152; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3154 = 8'h3a == total_offset_15 ? phv_data_58 : _GEN_3153; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3155 = 8'h3b == total_offset_15 ? phv_data_59 : _GEN_3154; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3156 = 8'h3c == total_offset_15 ? phv_data_60 : _GEN_3155; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3157 = 8'h3d == total_offset_15 ? phv_data_61 : _GEN_3156; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3158 = 8'h3e == total_offset_15 ? phv_data_62 : _GEN_3157; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3159 = 8'h3f == total_offset_15 ? phv_data_63 : _GEN_3158; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3160 = 8'h40 == total_offset_15 ? phv_data_64 : _GEN_3159; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3161 = 8'h41 == total_offset_15 ? phv_data_65 : _GEN_3160; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3162 = 8'h42 == total_offset_15 ? phv_data_66 : _GEN_3161; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3163 = 8'h43 == total_offset_15 ? phv_data_67 : _GEN_3162; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3164 = 8'h44 == total_offset_15 ? phv_data_68 : _GEN_3163; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3165 = 8'h45 == total_offset_15 ? phv_data_69 : _GEN_3164; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3166 = 8'h46 == total_offset_15 ? phv_data_70 : _GEN_3165; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3167 = 8'h47 == total_offset_15 ? phv_data_71 : _GEN_3166; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3168 = 8'h48 == total_offset_15 ? phv_data_72 : _GEN_3167; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3169 = 8'h49 == total_offset_15 ? phv_data_73 : _GEN_3168; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3170 = 8'h4a == total_offset_15 ? phv_data_74 : _GEN_3169; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3171 = 8'h4b == total_offset_15 ? phv_data_75 : _GEN_3170; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3172 = 8'h4c == total_offset_15 ? phv_data_76 : _GEN_3171; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3173 = 8'h4d == total_offset_15 ? phv_data_77 : _GEN_3172; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3174 = 8'h4e == total_offset_15 ? phv_data_78 : _GEN_3173; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3175 = 8'h4f == total_offset_15 ? phv_data_79 : _GEN_3174; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3176 = 8'h50 == total_offset_15 ? phv_data_80 : _GEN_3175; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3177 = 8'h51 == total_offset_15 ? phv_data_81 : _GEN_3176; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3178 = 8'h52 == total_offset_15 ? phv_data_82 : _GEN_3177; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3179 = 8'h53 == total_offset_15 ? phv_data_83 : _GEN_3178; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3180 = 8'h54 == total_offset_15 ? phv_data_84 : _GEN_3179; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3181 = 8'h55 == total_offset_15 ? phv_data_85 : _GEN_3180; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3182 = 8'h56 == total_offset_15 ? phv_data_86 : _GEN_3181; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3183 = 8'h57 == total_offset_15 ? phv_data_87 : _GEN_3182; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3184 = 8'h58 == total_offset_15 ? phv_data_88 : _GEN_3183; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3185 = 8'h59 == total_offset_15 ? phv_data_89 : _GEN_3184; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3186 = 8'h5a == total_offset_15 ? phv_data_90 : _GEN_3185; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3187 = 8'h5b == total_offset_15 ? phv_data_91 : _GEN_3186; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3188 = 8'h5c == total_offset_15 ? phv_data_92 : _GEN_3187; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3189 = 8'h5d == total_offset_15 ? phv_data_93 : _GEN_3188; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3190 = 8'h5e == total_offset_15 ? phv_data_94 : _GEN_3189; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3191 = 8'h5f == total_offset_15 ? phv_data_95 : _GEN_3190; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3192 = 8'h60 == total_offset_15 ? phv_data_96 : _GEN_3191; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3193 = 8'h61 == total_offset_15 ? phv_data_97 : _GEN_3192; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3194 = 8'h62 == total_offset_15 ? phv_data_98 : _GEN_3193; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3195 = 8'h63 == total_offset_15 ? phv_data_99 : _GEN_3194; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3196 = 8'h64 == total_offset_15 ? phv_data_100 : _GEN_3195; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3197 = 8'h65 == total_offset_15 ? phv_data_101 : _GEN_3196; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3198 = 8'h66 == total_offset_15 ? phv_data_102 : _GEN_3197; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3199 = 8'h67 == total_offset_15 ? phv_data_103 : _GEN_3198; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3200 = 8'h68 == total_offset_15 ? phv_data_104 : _GEN_3199; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3201 = 8'h69 == total_offset_15 ? phv_data_105 : _GEN_3200; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3202 = 8'h6a == total_offset_15 ? phv_data_106 : _GEN_3201; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3203 = 8'h6b == total_offset_15 ? phv_data_107 : _GEN_3202; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3204 = 8'h6c == total_offset_15 ? phv_data_108 : _GEN_3203; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3205 = 8'h6d == total_offset_15 ? phv_data_109 : _GEN_3204; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3206 = 8'h6e == total_offset_15 ? phv_data_110 : _GEN_3205; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3207 = 8'h6f == total_offset_15 ? phv_data_111 : _GEN_3206; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3208 = 8'h70 == total_offset_15 ? phv_data_112 : _GEN_3207; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3209 = 8'h71 == total_offset_15 ? phv_data_113 : _GEN_3208; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3210 = 8'h72 == total_offset_15 ? phv_data_114 : _GEN_3209; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3211 = 8'h73 == total_offset_15 ? phv_data_115 : _GEN_3210; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3212 = 8'h74 == total_offset_15 ? phv_data_116 : _GEN_3211; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3213 = 8'h75 == total_offset_15 ? phv_data_117 : _GEN_3212; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3214 = 8'h76 == total_offset_15 ? phv_data_118 : _GEN_3213; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3215 = 8'h77 == total_offset_15 ? phv_data_119 : _GEN_3214; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3216 = 8'h78 == total_offset_15 ? phv_data_120 : _GEN_3215; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3217 = 8'h79 == total_offset_15 ? phv_data_121 : _GEN_3216; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3218 = 8'h7a == total_offset_15 ? phv_data_122 : _GEN_3217; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3219 = 8'h7b == total_offset_15 ? phv_data_123 : _GEN_3218; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3220 = 8'h7c == total_offset_15 ? phv_data_124 : _GEN_3219; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3221 = 8'h7d == total_offset_15 ? phv_data_125 : _GEN_3220; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3222 = 8'h7e == total_offset_15 ? phv_data_126 : _GEN_3221; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3223 = 8'h7f == total_offset_15 ? phv_data_127 : _GEN_3222; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3224 = 8'h80 == total_offset_15 ? phv_data_128 : _GEN_3223; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3225 = 8'h81 == total_offset_15 ? phv_data_129 : _GEN_3224; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3226 = 8'h82 == total_offset_15 ? phv_data_130 : _GEN_3225; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3227 = 8'h83 == total_offset_15 ? phv_data_131 : _GEN_3226; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3228 = 8'h84 == total_offset_15 ? phv_data_132 : _GEN_3227; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3229 = 8'h85 == total_offset_15 ? phv_data_133 : _GEN_3228; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3230 = 8'h86 == total_offset_15 ? phv_data_134 : _GEN_3229; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3231 = 8'h87 == total_offset_15 ? phv_data_135 : _GEN_3230; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3232 = 8'h88 == total_offset_15 ? phv_data_136 : _GEN_3231; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3233 = 8'h89 == total_offset_15 ? phv_data_137 : _GEN_3232; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3234 = 8'h8a == total_offset_15 ? phv_data_138 : _GEN_3233; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3235 = 8'h8b == total_offset_15 ? phv_data_139 : _GEN_3234; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3236 = 8'h8c == total_offset_15 ? phv_data_140 : _GEN_3235; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3237 = 8'h8d == total_offset_15 ? phv_data_141 : _GEN_3236; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3238 = 8'h8e == total_offset_15 ? phv_data_142 : _GEN_3237; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3239 = 8'h8f == total_offset_15 ? phv_data_143 : _GEN_3238; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3240 = 8'h90 == total_offset_15 ? phv_data_144 : _GEN_3239; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3241 = 8'h91 == total_offset_15 ? phv_data_145 : _GEN_3240; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3242 = 8'h92 == total_offset_15 ? phv_data_146 : _GEN_3241; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3243 = 8'h93 == total_offset_15 ? phv_data_147 : _GEN_3242; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3244 = 8'h94 == total_offset_15 ? phv_data_148 : _GEN_3243; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3245 = 8'h95 == total_offset_15 ? phv_data_149 : _GEN_3244; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3246 = 8'h96 == total_offset_15 ? phv_data_150 : _GEN_3245; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3247 = 8'h97 == total_offset_15 ? phv_data_151 : _GEN_3246; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3248 = 8'h98 == total_offset_15 ? phv_data_152 : _GEN_3247; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3249 = 8'h99 == total_offset_15 ? phv_data_153 : _GEN_3248; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3250 = 8'h9a == total_offset_15 ? phv_data_154 : _GEN_3249; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3251 = 8'h9b == total_offset_15 ? phv_data_155 : _GEN_3250; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3252 = 8'h9c == total_offset_15 ? phv_data_156 : _GEN_3251; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3253 = 8'h9d == total_offset_15 ? phv_data_157 : _GEN_3252; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3254 = 8'h9e == total_offset_15 ? phv_data_158 : _GEN_3253; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes_3_0 = 8'h9f == total_offset_15 ? phv_data_159 : _GEN_3254; // @[executor.scala 197:66 executor.scala 197:66]
  wire [31:0] _io_field_out_3_T = {bytes_3_0,bytes_3_1,bytes_3_2,bytes_3_3}; // @[Cat.scala 30:58]
  wire [3:0] _io_mask_out_3_T = {_mask_3_T_24,mask_3_1,mask_3_2,mask_3_3}; // @[Cat.scala 30:58]
  wire [17:0] io_field_out_3_hi_4 = io_field_out_3_lo[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _io_field_out_3_T_4 = {io_field_out_3_hi_4,io_field_out_3_lo}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_3481 = 4'hb == opcode_3 ? _io_field_out_3_T_4 : 32'h0; // @[executor.scala 230:56 executor.scala 231:41]
  wire [1:0] _GEN_3482 = from_header_3 ? bias_3 : 2'h0; // @[executor.scala 178:36 executor.scala 203:36 executor.scala 174:29]
  wire [31:0] _GEN_3483 = from_header_3 ? _io_field_out_3_T : _GEN_3481; // @[executor.scala 178:36 executor.scala 204:37]
  wire [3:0] _GEN_3484 = from_header_3 ? _io_mask_out_3_T : 4'h0; // @[executor.scala 178:36 executor.scala 205:37 executor.scala 173:29]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_96 = phv_data_96; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_97 = phv_data_97; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_98 = phv_data_98; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_99 = phv_data_99; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_100 = phv_data_100; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_101 = phv_data_101; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_102 = phv_data_102; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_103 = phv_data_103; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_104 = phv_data_104; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_105 = phv_data_105; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_106 = phv_data_106; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_107 = phv_data_107; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_108 = phv_data_108; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_109 = phv_data_109; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_110 = phv_data_110; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_111 = phv_data_111; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_112 = phv_data_112; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_113 = phv_data_113; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_114 = phv_data_114; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_115 = phv_data_115; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_116 = phv_data_116; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_117 = phv_data_117; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_118 = phv_data_118; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_119 = phv_data_119; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_120 = phv_data_120; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_121 = phv_data_121; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_122 = phv_data_122; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_123 = phv_data_123; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_124 = phv_data_124; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_125 = phv_data_125; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_126 = phv_data_126; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_127 = phv_data_127; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_128 = phv_data_128; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_129 = phv_data_129; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_130 = phv_data_130; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_131 = phv_data_131; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_132 = phv_data_132; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_133 = phv_data_133; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_134 = phv_data_134; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_135 = phv_data_135; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_136 = phv_data_136; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_137 = phv_data_137; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_138 = phv_data_138; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_139 = phv_data_139; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_140 = phv_data_140; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_141 = phv_data_141; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_142 = phv_data_142; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_143 = phv_data_143; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_144 = phv_data_144; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_145 = phv_data_145; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_146 = phv_data_146; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_147 = phv_data_147; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_148 = phv_data_148; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_149 = phv_data_149; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_150 = phv_data_150; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_151 = phv_data_151; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_152 = phv_data_152; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_153 = phv_data_153; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_154 = phv_data_154; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_155 = phv_data_155; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_156 = phv_data_156; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_157 = phv_data_157; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_158 = phv_data_158; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_159 = phv_data_159; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[executor.scala 153:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[executor.scala 153:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[executor.scala 153:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[executor.scala 153:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[executor.scala 153:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[executor.scala 153:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[executor.scala 153:25]
  assign io_pipe_phv_out_valid = phv_valid; // @[executor.scala 153:25]
  assign io_pipe_phv_out_last = phv_last; // @[executor.scala 153:25]
  assign io_vliw_out_0 = vliw_0; // @[executor.scala 160:21]
  assign io_vliw_out_1 = vliw_1; // @[executor.scala 160:21]
  assign io_vliw_out_2 = vliw_2; // @[executor.scala 160:21]
  assign io_vliw_out_3 = vliw_3; // @[executor.scala 160:21]
  assign io_field_out_0 = phv_is_valid_processor ? _GEN_867 : 32'h0; // @[executor.scala 176:43 executor.scala 172:29]
  assign io_field_out_1 = phv_is_valid_processor ? _GEN_1739 : 32'h0; // @[executor.scala 176:43 executor.scala 172:29]
  assign io_field_out_2 = phv_is_valid_processor ? _GEN_2611 : 32'h0; // @[executor.scala 176:43 executor.scala 172:29]
  assign io_field_out_3 = phv_is_valid_processor ? _GEN_3483 : 32'h0; // @[executor.scala 176:43 executor.scala 172:29]
  assign io_mask_out_0 = phv_is_valid_processor ? _GEN_868 : 4'h0; // @[executor.scala 176:43 executor.scala 173:29]
  assign io_mask_out_1 = phv_is_valid_processor ? _GEN_1740 : 4'h0; // @[executor.scala 176:43 executor.scala 173:29]
  assign io_mask_out_2 = phv_is_valid_processor ? _GEN_2612 : 4'h0; // @[executor.scala 176:43 executor.scala 173:29]
  assign io_mask_out_3 = phv_is_valid_processor ? _GEN_3484 : 4'h0; // @[executor.scala 176:43 executor.scala 173:29]
  assign io_bias_out_0 = phv_is_valid_processor ? _GEN_866 : 2'h0; // @[executor.scala 176:43 executor.scala 174:29]
  assign io_bias_out_1 = phv_is_valid_processor ? _GEN_1738 : 2'h0; // @[executor.scala 176:43 executor.scala 174:29]
  assign io_bias_out_2 = phv_is_valid_processor ? _GEN_2610 : 2'h0; // @[executor.scala 176:43 executor.scala 174:29]
  assign io_bias_out_3 = phv_is_valid_processor ? _GEN_3482 : 2'h0; // @[executor.scala 176:43 executor.scala 174:29]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[executor.scala 152:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[executor.scala 152:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[executor.scala 152:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[executor.scala 152:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[executor.scala 152:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[executor.scala 152:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[executor.scala 152:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[executor.scala 152:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[executor.scala 152:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[executor.scala 152:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[executor.scala 152:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[executor.scala 152:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[executor.scala 152:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[executor.scala 152:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[executor.scala 152:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[executor.scala 152:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[executor.scala 152:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[executor.scala 152:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[executor.scala 152:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[executor.scala 152:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[executor.scala 152:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[executor.scala 152:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[executor.scala 152:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[executor.scala 152:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[executor.scala 152:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[executor.scala 152:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[executor.scala 152:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[executor.scala 152:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[executor.scala 152:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[executor.scala 152:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[executor.scala 152:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[executor.scala 152:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[executor.scala 152:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[executor.scala 152:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[executor.scala 152:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[executor.scala 152:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[executor.scala 152:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[executor.scala 152:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[executor.scala 152:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[executor.scala 152:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[executor.scala 152:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[executor.scala 152:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[executor.scala 152:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[executor.scala 152:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[executor.scala 152:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[executor.scala 152:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[executor.scala 152:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[executor.scala 152:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[executor.scala 152:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[executor.scala 152:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[executor.scala 152:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[executor.scala 152:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[executor.scala 152:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[executor.scala 152:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[executor.scala 152:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[executor.scala 152:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[executor.scala 152:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[executor.scala 152:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[executor.scala 152:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[executor.scala 152:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[executor.scala 152:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[executor.scala 152:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[executor.scala 152:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[executor.scala 152:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[executor.scala 152:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[executor.scala 152:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[executor.scala 152:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[executor.scala 152:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[executor.scala 152:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[executor.scala 152:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[executor.scala 152:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[executor.scala 152:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[executor.scala 152:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[executor.scala 152:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[executor.scala 152:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[executor.scala 152:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[executor.scala 152:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[executor.scala 152:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[executor.scala 152:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[executor.scala 152:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[executor.scala 152:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[executor.scala 152:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[executor.scala 152:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[executor.scala 152:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[executor.scala 152:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[executor.scala 152:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[executor.scala 152:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[executor.scala 152:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[executor.scala 152:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[executor.scala 152:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[executor.scala 152:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[executor.scala 152:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[executor.scala 152:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[executor.scala 152:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[executor.scala 152:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[executor.scala 152:13]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[executor.scala 152:13]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[executor.scala 152:13]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[executor.scala 152:13]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[executor.scala 152:13]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[executor.scala 152:13]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[executor.scala 152:13]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[executor.scala 152:13]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[executor.scala 152:13]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[executor.scala 152:13]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[executor.scala 152:13]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[executor.scala 152:13]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[executor.scala 152:13]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[executor.scala 152:13]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[executor.scala 152:13]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[executor.scala 152:13]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[executor.scala 152:13]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[executor.scala 152:13]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[executor.scala 152:13]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[executor.scala 152:13]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[executor.scala 152:13]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[executor.scala 152:13]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[executor.scala 152:13]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[executor.scala 152:13]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[executor.scala 152:13]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[executor.scala 152:13]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[executor.scala 152:13]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[executor.scala 152:13]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[executor.scala 152:13]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[executor.scala 152:13]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[executor.scala 152:13]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[executor.scala 152:13]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[executor.scala 152:13]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[executor.scala 152:13]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[executor.scala 152:13]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[executor.scala 152:13]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[executor.scala 152:13]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[executor.scala 152:13]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[executor.scala 152:13]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[executor.scala 152:13]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[executor.scala 152:13]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[executor.scala 152:13]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[executor.scala 152:13]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[executor.scala 152:13]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[executor.scala 152:13]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[executor.scala 152:13]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[executor.scala 152:13]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[executor.scala 152:13]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[executor.scala 152:13]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[executor.scala 152:13]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[executor.scala 152:13]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[executor.scala 152:13]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[executor.scala 152:13]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[executor.scala 152:13]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[executor.scala 152:13]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[executor.scala 152:13]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[executor.scala 152:13]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[executor.scala 152:13]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[executor.scala 152:13]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[executor.scala 152:13]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[executor.scala 152:13]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[executor.scala 152:13]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[executor.scala 152:13]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[executor.scala 152:13]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[executor.scala 152:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[executor.scala 152:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[executor.scala 152:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[executor.scala 152:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[executor.scala 152:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[executor.scala 152:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[executor.scala 152:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[executor.scala 152:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[executor.scala 152:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[executor.scala 152:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[executor.scala 152:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[executor.scala 152:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[executor.scala 152:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[executor.scala 152:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[executor.scala 152:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[executor.scala 152:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[executor.scala 152:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[executor.scala 152:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[executor.scala 152:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[executor.scala 152:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[executor.scala 152:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[executor.scala 152:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[executor.scala 152:13]
    phv_valid <= io_pipe_phv_in_valid; // @[executor.scala 152:13]
    phv_last <= io_pipe_phv_in_last; // @[executor.scala 152:13]
    vliw_0 <= io_vliw_in_0; // @[executor.scala 159:14]
    vliw_1 <= io_vliw_in_1; // @[executor.scala 159:14]
    vliw_2 <= io_vliw_in_2; // @[executor.scala 159:14]
    vliw_3 <= io_vliw_in_3; // @[executor.scala 159:14]
    offset_0 <= io_offset_in_0; // @[executor.scala 164:16]
    offset_1 <= io_offset_in_1; // @[executor.scala 164:16]
    offset_2 <= io_offset_in_2; // @[executor.scala 164:16]
    offset_3 <= io_offset_in_3; // @[executor.scala 164:16]
    length_0 <= io_length_in_0; // @[executor.scala 165:16]
    length_1 <= io_length_in_1; // @[executor.scala 165:16]
    length_2 <= io_length_in_2; // @[executor.scala 165:16]
    length_3 <= io_length_in_3; // @[executor.scala 165:16]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_header_0 = _RAND_160[15:0];
  _RAND_161 = {1{`RANDOM}};
  phv_header_1 = _RAND_161[15:0];
  _RAND_162 = {1{`RANDOM}};
  phv_header_2 = _RAND_162[15:0];
  _RAND_163 = {1{`RANDOM}};
  phv_header_3 = _RAND_163[15:0];
  _RAND_164 = {1{`RANDOM}};
  phv_header_4 = _RAND_164[15:0];
  _RAND_165 = {1{`RANDOM}};
  phv_header_5 = _RAND_165[15:0];
  _RAND_166 = {1{`RANDOM}};
  phv_header_6 = _RAND_166[15:0];
  _RAND_167 = {1{`RANDOM}};
  phv_header_7 = _RAND_167[15:0];
  _RAND_168 = {1{`RANDOM}};
  phv_header_8 = _RAND_168[15:0];
  _RAND_169 = {1{`RANDOM}};
  phv_header_9 = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  phv_header_10 = _RAND_170[15:0];
  _RAND_171 = {1{`RANDOM}};
  phv_header_11 = _RAND_171[15:0];
  _RAND_172 = {1{`RANDOM}};
  phv_header_12 = _RAND_172[15:0];
  _RAND_173 = {1{`RANDOM}};
  phv_header_13 = _RAND_173[15:0];
  _RAND_174 = {1{`RANDOM}};
  phv_header_14 = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  phv_header_15 = _RAND_175[15:0];
  _RAND_176 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_178[15:0];
  _RAND_179 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_179[3:0];
  _RAND_180 = {1{`RANDOM}};
  phv_next_config_id = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  phv_valid = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  phv_last = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  vliw_0 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  vliw_1 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  vliw_2 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  vliw_3 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  offset_0 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  offset_1 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  offset_2 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  offset_3 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  length_0 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  length_1 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  length_2 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  length_3 = _RAND_195[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
