module ParseAction(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [7:0]  io_pipe_phv_in_data_160,
  input  [7:0]  io_pipe_phv_in_data_161,
  input  [7:0]  io_pipe_phv_in_data_162,
  input  [7:0]  io_pipe_phv_in_data_163,
  input  [7:0]  io_pipe_phv_in_data_164,
  input  [7:0]  io_pipe_phv_in_data_165,
  input  [7:0]  io_pipe_phv_in_data_166,
  input  [7:0]  io_pipe_phv_in_data_167,
  input  [7:0]  io_pipe_phv_in_data_168,
  input  [7:0]  io_pipe_phv_in_data_169,
  input  [7:0]  io_pipe_phv_in_data_170,
  input  [7:0]  io_pipe_phv_in_data_171,
  input  [7:0]  io_pipe_phv_in_data_172,
  input  [7:0]  io_pipe_phv_in_data_173,
  input  [7:0]  io_pipe_phv_in_data_174,
  input  [7:0]  io_pipe_phv_in_data_175,
  input  [7:0]  io_pipe_phv_in_data_176,
  input  [7:0]  io_pipe_phv_in_data_177,
  input  [7:0]  io_pipe_phv_in_data_178,
  input  [7:0]  io_pipe_phv_in_data_179,
  input  [7:0]  io_pipe_phv_in_data_180,
  input  [7:0]  io_pipe_phv_in_data_181,
  input  [7:0]  io_pipe_phv_in_data_182,
  input  [7:0]  io_pipe_phv_in_data_183,
  input  [7:0]  io_pipe_phv_in_data_184,
  input  [7:0]  io_pipe_phv_in_data_185,
  input  [7:0]  io_pipe_phv_in_data_186,
  input  [7:0]  io_pipe_phv_in_data_187,
  input  [7:0]  io_pipe_phv_in_data_188,
  input  [7:0]  io_pipe_phv_in_data_189,
  input  [7:0]  io_pipe_phv_in_data_190,
  input  [7:0]  io_pipe_phv_in_data_191,
  input  [7:0]  io_pipe_phv_in_data_192,
  input  [7:0]  io_pipe_phv_in_data_193,
  input  [7:0]  io_pipe_phv_in_data_194,
  input  [7:0]  io_pipe_phv_in_data_195,
  input  [7:0]  io_pipe_phv_in_data_196,
  input  [7:0]  io_pipe_phv_in_data_197,
  input  [7:0]  io_pipe_phv_in_data_198,
  input  [7:0]  io_pipe_phv_in_data_199,
  input  [7:0]  io_pipe_phv_in_data_200,
  input  [7:0]  io_pipe_phv_in_data_201,
  input  [7:0]  io_pipe_phv_in_data_202,
  input  [7:0]  io_pipe_phv_in_data_203,
  input  [7:0]  io_pipe_phv_in_data_204,
  input  [7:0]  io_pipe_phv_in_data_205,
  input  [7:0]  io_pipe_phv_in_data_206,
  input  [7:0]  io_pipe_phv_in_data_207,
  input  [7:0]  io_pipe_phv_in_data_208,
  input  [7:0]  io_pipe_phv_in_data_209,
  input  [7:0]  io_pipe_phv_in_data_210,
  input  [7:0]  io_pipe_phv_in_data_211,
  input  [7:0]  io_pipe_phv_in_data_212,
  input  [7:0]  io_pipe_phv_in_data_213,
  input  [7:0]  io_pipe_phv_in_data_214,
  input  [7:0]  io_pipe_phv_in_data_215,
  input  [7:0]  io_pipe_phv_in_data_216,
  input  [7:0]  io_pipe_phv_in_data_217,
  input  [7:0]  io_pipe_phv_in_data_218,
  input  [7:0]  io_pipe_phv_in_data_219,
  input  [7:0]  io_pipe_phv_in_data_220,
  input  [7:0]  io_pipe_phv_in_data_221,
  input  [7:0]  io_pipe_phv_in_data_222,
  input  [7:0]  io_pipe_phv_in_data_223,
  input  [7:0]  io_pipe_phv_in_data_224,
  input  [7:0]  io_pipe_phv_in_data_225,
  input  [7:0]  io_pipe_phv_in_data_226,
  input  [7:0]  io_pipe_phv_in_data_227,
  input  [7:0]  io_pipe_phv_in_data_228,
  input  [7:0]  io_pipe_phv_in_data_229,
  input  [7:0]  io_pipe_phv_in_data_230,
  input  [7:0]  io_pipe_phv_in_data_231,
  input  [7:0]  io_pipe_phv_in_data_232,
  input  [7:0]  io_pipe_phv_in_data_233,
  input  [7:0]  io_pipe_phv_in_data_234,
  input  [7:0]  io_pipe_phv_in_data_235,
  input  [7:0]  io_pipe_phv_in_data_236,
  input  [7:0]  io_pipe_phv_in_data_237,
  input  [7:0]  io_pipe_phv_in_data_238,
  input  [7:0]  io_pipe_phv_in_data_239,
  input  [7:0]  io_pipe_phv_in_data_240,
  input  [7:0]  io_pipe_phv_in_data_241,
  input  [7:0]  io_pipe_phv_in_data_242,
  input  [7:0]  io_pipe_phv_in_data_243,
  input  [7:0]  io_pipe_phv_in_data_244,
  input  [7:0]  io_pipe_phv_in_data_245,
  input  [7:0]  io_pipe_phv_in_data_246,
  input  [7:0]  io_pipe_phv_in_data_247,
  input  [7:0]  io_pipe_phv_in_data_248,
  input  [7:0]  io_pipe_phv_in_data_249,
  input  [7:0]  io_pipe_phv_in_data_250,
  input  [7:0]  io_pipe_phv_in_data_251,
  input  [7:0]  io_pipe_phv_in_data_252,
  input  [7:0]  io_pipe_phv_in_data_253,
  input  [7:0]  io_pipe_phv_in_data_254,
  input  [7:0]  io_pipe_phv_in_data_255,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [7:0]  io_pipe_phv_out_data_160,
  output [7:0]  io_pipe_phv_out_data_161,
  output [7:0]  io_pipe_phv_out_data_162,
  output [7:0]  io_pipe_phv_out_data_163,
  output [7:0]  io_pipe_phv_out_data_164,
  output [7:0]  io_pipe_phv_out_data_165,
  output [7:0]  io_pipe_phv_out_data_166,
  output [7:0]  io_pipe_phv_out_data_167,
  output [7:0]  io_pipe_phv_out_data_168,
  output [7:0]  io_pipe_phv_out_data_169,
  output [7:0]  io_pipe_phv_out_data_170,
  output [7:0]  io_pipe_phv_out_data_171,
  output [7:0]  io_pipe_phv_out_data_172,
  output [7:0]  io_pipe_phv_out_data_173,
  output [7:0]  io_pipe_phv_out_data_174,
  output [7:0]  io_pipe_phv_out_data_175,
  output [7:0]  io_pipe_phv_out_data_176,
  output [7:0]  io_pipe_phv_out_data_177,
  output [7:0]  io_pipe_phv_out_data_178,
  output [7:0]  io_pipe_phv_out_data_179,
  output [7:0]  io_pipe_phv_out_data_180,
  output [7:0]  io_pipe_phv_out_data_181,
  output [7:0]  io_pipe_phv_out_data_182,
  output [7:0]  io_pipe_phv_out_data_183,
  output [7:0]  io_pipe_phv_out_data_184,
  output [7:0]  io_pipe_phv_out_data_185,
  output [7:0]  io_pipe_phv_out_data_186,
  output [7:0]  io_pipe_phv_out_data_187,
  output [7:0]  io_pipe_phv_out_data_188,
  output [7:0]  io_pipe_phv_out_data_189,
  output [7:0]  io_pipe_phv_out_data_190,
  output [7:0]  io_pipe_phv_out_data_191,
  output [7:0]  io_pipe_phv_out_data_192,
  output [7:0]  io_pipe_phv_out_data_193,
  output [7:0]  io_pipe_phv_out_data_194,
  output [7:0]  io_pipe_phv_out_data_195,
  output [7:0]  io_pipe_phv_out_data_196,
  output [7:0]  io_pipe_phv_out_data_197,
  output [7:0]  io_pipe_phv_out_data_198,
  output [7:0]  io_pipe_phv_out_data_199,
  output [7:0]  io_pipe_phv_out_data_200,
  output [7:0]  io_pipe_phv_out_data_201,
  output [7:0]  io_pipe_phv_out_data_202,
  output [7:0]  io_pipe_phv_out_data_203,
  output [7:0]  io_pipe_phv_out_data_204,
  output [7:0]  io_pipe_phv_out_data_205,
  output [7:0]  io_pipe_phv_out_data_206,
  output [7:0]  io_pipe_phv_out_data_207,
  output [7:0]  io_pipe_phv_out_data_208,
  output [7:0]  io_pipe_phv_out_data_209,
  output [7:0]  io_pipe_phv_out_data_210,
  output [7:0]  io_pipe_phv_out_data_211,
  output [7:0]  io_pipe_phv_out_data_212,
  output [7:0]  io_pipe_phv_out_data_213,
  output [7:0]  io_pipe_phv_out_data_214,
  output [7:0]  io_pipe_phv_out_data_215,
  output [7:0]  io_pipe_phv_out_data_216,
  output [7:0]  io_pipe_phv_out_data_217,
  output [7:0]  io_pipe_phv_out_data_218,
  output [7:0]  io_pipe_phv_out_data_219,
  output [7:0]  io_pipe_phv_out_data_220,
  output [7:0]  io_pipe_phv_out_data_221,
  output [7:0]  io_pipe_phv_out_data_222,
  output [7:0]  io_pipe_phv_out_data_223,
  output [7:0]  io_pipe_phv_out_data_224,
  output [7:0]  io_pipe_phv_out_data_225,
  output [7:0]  io_pipe_phv_out_data_226,
  output [7:0]  io_pipe_phv_out_data_227,
  output [7:0]  io_pipe_phv_out_data_228,
  output [7:0]  io_pipe_phv_out_data_229,
  output [7:0]  io_pipe_phv_out_data_230,
  output [7:0]  io_pipe_phv_out_data_231,
  output [7:0]  io_pipe_phv_out_data_232,
  output [7:0]  io_pipe_phv_out_data_233,
  output [7:0]  io_pipe_phv_out_data_234,
  output [7:0]  io_pipe_phv_out_data_235,
  output [7:0]  io_pipe_phv_out_data_236,
  output [7:0]  io_pipe_phv_out_data_237,
  output [7:0]  io_pipe_phv_out_data_238,
  output [7:0]  io_pipe_phv_out_data_239,
  output [7:0]  io_pipe_phv_out_data_240,
  output [7:0]  io_pipe_phv_out_data_241,
  output [7:0]  io_pipe_phv_out_data_242,
  output [7:0]  io_pipe_phv_out_data_243,
  output [7:0]  io_pipe_phv_out_data_244,
  output [7:0]  io_pipe_phv_out_data_245,
  output [7:0]  io_pipe_phv_out_data_246,
  output [7:0]  io_pipe_phv_out_data_247,
  output [7:0]  io_pipe_phv_out_data_248,
  output [7:0]  io_pipe_phv_out_data_249,
  output [7:0]  io_pipe_phv_out_data_250,
  output [7:0]  io_pipe_phv_out_data_251,
  output [7:0]  io_pipe_phv_out_data_252,
  output [7:0]  io_pipe_phv_out_data_253,
  output [7:0]  io_pipe_phv_out_data_254,
  output [7:0]  io_pipe_phv_out_data_255,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input  [63:0] io_rdata,
  input         io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_1; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_2; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_3; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_4; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_5; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_6; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_7; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_8; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_9; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_10; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_11; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_12; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_13; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_14; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_15; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_16; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_17; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_18; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_19; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_20; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_21; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_22; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_23; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_24; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_25; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_26; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_27; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_28; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_29; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_30; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_31; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_32; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_33; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_34; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_35; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_36; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_37; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_38; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_39; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_40; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_41; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_42; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_43; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_44; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_45; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_46; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_47; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_48; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_49; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_50; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_51; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_52; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_53; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_54; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_55; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_56; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_57; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_58; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_59; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_60; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_61; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_62; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_63; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_64; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_65; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_66; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_67; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_68; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_69; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_70; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_71; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_72; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_73; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_74; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_75; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_76; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_77; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_78; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_79; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_80; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_81; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_82; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_83; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_84; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_85; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_86; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_87; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_88; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_89; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_90; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_91; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_92; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_93; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_94; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_95; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_96; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_97; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_98; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_99; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_100; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_101; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_102; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_103; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_104; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_105; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_106; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_107; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_108; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_109; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_110; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_111; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_112; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_113; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_114; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_115; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_116; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_117; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_118; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_119; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_120; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_121; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_122; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_123; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_124; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_125; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_126; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_127; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_128; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_129; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_130; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_131; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_132; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_133; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_134; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_135; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_136; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_137; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_138; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_139; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_140; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_141; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_142; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_143; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_144; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_145; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_146; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_147; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_148; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_149; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_150; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_151; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_152; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_153; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_154; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_155; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_156; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_157; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_158; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_159; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_160; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_161; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_162; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_163; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_164; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_165; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_166; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_167; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_168; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_169; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_170; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_171; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_172; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_173; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_174; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_175; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_176; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_177; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_178; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_179; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_180; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_181; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_182; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_183; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_184; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_185; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_186; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_187; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_188; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_189; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_190; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_191; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_192; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_193; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_194; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_195; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_196; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_197; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_198; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_199; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_200; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_201; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_202; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_203; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_204; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_205; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_206; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_207; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_208; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_209; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_210; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_211; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_212; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_213; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_214; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_215; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_216; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_217; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_218; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_219; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_220; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_221; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_222; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_223; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_224; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_225; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_226; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_227; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_228; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_229; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_230; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_231; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_232; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_233; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_234; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_235; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_236; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_237; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_238; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_239; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_240; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_241; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_242; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_243; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_244; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_245; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_246; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_247; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_248; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_249; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_250; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_251; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_252; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_253; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_254; // @[parse_module.scala 50:20]
  reg [7:0] phv_data_255; // @[parse_module.scala 50:20]
  reg [15:0] phv_header_0; // @[parse_module.scala 50:20]
  reg [15:0] phv_header_1; // @[parse_module.scala 50:20]
  reg [15:0] phv_header_2; // @[parse_module.scala 50:20]
  reg [15:0] phv_header_3; // @[parse_module.scala 50:20]
  reg [15:0] phv_header_4; // @[parse_module.scala 50:20]
  reg [15:0] phv_header_5; // @[parse_module.scala 50:20]
  reg [15:0] phv_header_6; // @[parse_module.scala 50:20]
  reg [15:0] phv_header_7; // @[parse_module.scala 50:20]
  reg [15:0] phv_header_8; // @[parse_module.scala 50:20]
  reg [15:0] phv_header_9; // @[parse_module.scala 50:20]
  reg [15:0] phv_header_10; // @[parse_module.scala 50:20]
  reg [15:0] phv_header_11; // @[parse_module.scala 50:20]
  reg [15:0] phv_header_12; // @[parse_module.scala 50:20]
  reg [15:0] phv_header_13; // @[parse_module.scala 50:20]
  reg [15:0] phv_header_14; // @[parse_module.scala 50:20]
  reg [15:0] phv_header_15; // @[parse_module.scala 50:20]
  reg [7:0] phv_parse_current_state; // @[parse_module.scala 50:20]
  reg [7:0] phv_parse_current_offset; // @[parse_module.scala 50:20]
  reg [15:0] phv_parse_transition_field; // @[parse_module.scala 50:20]
  reg  phv_next_config_id; // @[parse_module.scala 50:20]
  reg  phv_is_valid_processor; // @[parse_module.scala 50:20]
  wire  is_valid = io_valid & io_pipe_phv_in_is_valid_processor; // @[parse_module.scala 54:29]
  wire [7:0] match_val_transition_field_header_id = io_rdata[55:48]; // @[parse_module.scala 59:61]
  wire [15:0] match_val_transition_field_mask = io_rdata[47:32]; // @[parse_module.scala 60:61]
  wire [7:0] match_val_transition_field_internal_offset = io_rdata[31:24]; // @[parse_module.scala 62:67]
  wire [7:0] phv_header_lo = io_rdata[23:16]; // @[parse_module.scala 63:50]
  wire [7:0] match_val_header_id = io_rdata[15:8]; // @[parse_module.scala 64:50]
  wire [7:0] match_val_next_state = io_rdata[7:0]; // @[parse_module.scala 65:50]
  wire [7:0] _phv_parse_current_offset_T_1 = io_pipe_phv_in_parse_current_offset + phv_header_lo; // @[parse_module.scala 68:73]
  wire [15:0] _GEN_1 = 4'h1 == match_val_transition_field_header_id[3:0] ? io_pipe_phv_in_header_1 :
    io_pipe_phv_in_header_0; // @[const.scala 34:43 const.scala 34:43]
  wire [15:0] _GEN_2 = 4'h2 == match_val_transition_field_header_id[3:0] ? io_pipe_phv_in_header_2 : _GEN_1; // @[const.scala 34:43 const.scala 34:43]
  wire [15:0] _GEN_3 = 4'h3 == match_val_transition_field_header_id[3:0] ? io_pipe_phv_in_header_3 : _GEN_2; // @[const.scala 34:43 const.scala 34:43]
  wire [15:0] _GEN_4 = 4'h4 == match_val_transition_field_header_id[3:0] ? io_pipe_phv_in_header_4 : _GEN_3; // @[const.scala 34:43 const.scala 34:43]
  wire [15:0] _GEN_5 = 4'h5 == match_val_transition_field_header_id[3:0] ? io_pipe_phv_in_header_5 : _GEN_4; // @[const.scala 34:43 const.scala 34:43]
  wire [15:0] _GEN_6 = 4'h6 == match_val_transition_field_header_id[3:0] ? io_pipe_phv_in_header_6 : _GEN_5; // @[const.scala 34:43 const.scala 34:43]
  wire [15:0] _GEN_7 = 4'h7 == match_val_transition_field_header_id[3:0] ? io_pipe_phv_in_header_7 : _GEN_6; // @[const.scala 34:43 const.scala 34:43]
  wire [15:0] _GEN_8 = 4'h8 == match_val_transition_field_header_id[3:0] ? io_pipe_phv_in_header_8 : _GEN_7; // @[const.scala 34:43 const.scala 34:43]
  wire [15:0] _GEN_9 = 4'h9 == match_val_transition_field_header_id[3:0] ? io_pipe_phv_in_header_9 : _GEN_8; // @[const.scala 34:43 const.scala 34:43]
  wire [15:0] _GEN_10 = 4'ha == match_val_transition_field_header_id[3:0] ? io_pipe_phv_in_header_10 : _GEN_9; // @[const.scala 34:43 const.scala 34:43]
  wire [15:0] _GEN_11 = 4'hb == match_val_transition_field_header_id[3:0] ? io_pipe_phv_in_header_11 : _GEN_10; // @[const.scala 34:43 const.scala 34:43]
  wire [15:0] _GEN_12 = 4'hc == match_val_transition_field_header_id[3:0] ? io_pipe_phv_in_header_12 : _GEN_11; // @[const.scala 34:43 const.scala 34:43]
  wire [15:0] _GEN_13 = 4'hd == match_val_transition_field_header_id[3:0] ? io_pipe_phv_in_header_13 : _GEN_12; // @[const.scala 34:43 const.scala 34:43]
  wire [15:0] _GEN_14 = 4'he == match_val_transition_field_header_id[3:0] ? io_pipe_phv_in_header_14 : _GEN_13; // @[const.scala 34:43 const.scala 34:43]
  wire [15:0] _GEN_15 = 4'hf == match_val_transition_field_header_id[3:0] ? io_pipe_phv_in_header_15 : _GEN_14; // @[const.scala 34:43 const.scala 34:43]
  wire [7:0] transition_field_header_offset = _GEN_15[15:8]; // @[const.scala 34:43]
  wire [7:0] transition_field_offset = transition_field_header_offset + match_val_transition_field_internal_offset; // @[parse_module.scala 71:70]
  wire [7:0] _transition_field_raw_data_T_1 = transition_field_offset + 8'h1; // @[parse_module.scala 73:57]
  wire [7:0] _GEN_17 = 8'h1 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_1 : io_pipe_phv_in_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_18 = 8'h2 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_2 : _GEN_17; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_19 = 8'h3 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_3 : _GEN_18; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_20 = 8'h4 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_4 : _GEN_19; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_21 = 8'h5 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_5 : _GEN_20; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_22 = 8'h6 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_6 : _GEN_21; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_23 = 8'h7 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_7 : _GEN_22; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_24 = 8'h8 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_8 : _GEN_23; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_25 = 8'h9 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_9 : _GEN_24; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_26 = 8'ha == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_10 : _GEN_25; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_27 = 8'hb == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_11 : _GEN_26; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_28 = 8'hc == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_12 : _GEN_27; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_29 = 8'hd == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_13 : _GEN_28; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_30 = 8'he == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_14 : _GEN_29; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_31 = 8'hf == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_15 : _GEN_30; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_32 = 8'h10 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_16 : _GEN_31; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_33 = 8'h11 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_17 : _GEN_32; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_34 = 8'h12 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_18 : _GEN_33; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_35 = 8'h13 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_19 : _GEN_34; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_36 = 8'h14 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_20 : _GEN_35; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_37 = 8'h15 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_21 : _GEN_36; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_38 = 8'h16 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_22 : _GEN_37; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_39 = 8'h17 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_23 : _GEN_38; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_40 = 8'h18 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_24 : _GEN_39; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_41 = 8'h19 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_25 : _GEN_40; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_42 = 8'h1a == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_26 : _GEN_41; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_43 = 8'h1b == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_27 : _GEN_42; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_44 = 8'h1c == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_28 : _GEN_43; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_45 = 8'h1d == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_29 : _GEN_44; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_46 = 8'h1e == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_30 : _GEN_45; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_47 = 8'h1f == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_31 : _GEN_46; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_48 = 8'h20 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_32 : _GEN_47; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_49 = 8'h21 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_33 : _GEN_48; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_50 = 8'h22 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_34 : _GEN_49; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_51 = 8'h23 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_35 : _GEN_50; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_52 = 8'h24 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_36 : _GEN_51; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_53 = 8'h25 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_37 : _GEN_52; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_54 = 8'h26 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_38 : _GEN_53; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_55 = 8'h27 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_39 : _GEN_54; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_56 = 8'h28 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_40 : _GEN_55; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_57 = 8'h29 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_41 : _GEN_56; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_58 = 8'h2a == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_42 : _GEN_57; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_59 = 8'h2b == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_43 : _GEN_58; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_60 = 8'h2c == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_44 : _GEN_59; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_61 = 8'h2d == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_45 : _GEN_60; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_62 = 8'h2e == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_46 : _GEN_61; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_63 = 8'h2f == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_47 : _GEN_62; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_64 = 8'h30 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_48 : _GEN_63; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_65 = 8'h31 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_49 : _GEN_64; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_66 = 8'h32 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_50 : _GEN_65; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_67 = 8'h33 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_51 : _GEN_66; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_68 = 8'h34 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_52 : _GEN_67; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_69 = 8'h35 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_53 : _GEN_68; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_70 = 8'h36 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_54 : _GEN_69; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_71 = 8'h37 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_55 : _GEN_70; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_72 = 8'h38 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_56 : _GEN_71; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_73 = 8'h39 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_57 : _GEN_72; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_74 = 8'h3a == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_58 : _GEN_73; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_75 = 8'h3b == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_59 : _GEN_74; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_76 = 8'h3c == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_60 : _GEN_75; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_77 = 8'h3d == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_61 : _GEN_76; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_78 = 8'h3e == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_62 : _GEN_77; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_79 = 8'h3f == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_63 : _GEN_78; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_80 = 8'h40 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_64 : _GEN_79; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_81 = 8'h41 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_65 : _GEN_80; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_82 = 8'h42 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_66 : _GEN_81; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_83 = 8'h43 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_67 : _GEN_82; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_84 = 8'h44 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_68 : _GEN_83; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_85 = 8'h45 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_69 : _GEN_84; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_86 = 8'h46 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_70 : _GEN_85; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_87 = 8'h47 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_71 : _GEN_86; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_88 = 8'h48 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_72 : _GEN_87; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_89 = 8'h49 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_73 : _GEN_88; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_90 = 8'h4a == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_74 : _GEN_89; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_91 = 8'h4b == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_75 : _GEN_90; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_92 = 8'h4c == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_76 : _GEN_91; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_93 = 8'h4d == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_77 : _GEN_92; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_94 = 8'h4e == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_78 : _GEN_93; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_95 = 8'h4f == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_79 : _GEN_94; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_96 = 8'h50 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_80 : _GEN_95; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_97 = 8'h51 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_81 : _GEN_96; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_98 = 8'h52 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_82 : _GEN_97; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_99 = 8'h53 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_83 : _GEN_98; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_100 = 8'h54 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_84 : _GEN_99; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_101 = 8'h55 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_85 : _GEN_100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_102 = 8'h56 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_86 : _GEN_101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_103 = 8'h57 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_87 : _GEN_102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_104 = 8'h58 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_88 : _GEN_103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_105 = 8'h59 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_89 : _GEN_104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_106 = 8'h5a == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_90 : _GEN_105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_107 = 8'h5b == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_91 : _GEN_106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_108 = 8'h5c == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_92 : _GEN_107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_109 = 8'h5d == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_93 : _GEN_108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_110 = 8'h5e == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_94 : _GEN_109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_111 = 8'h5f == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_95 : _GEN_110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_112 = 8'h60 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_96 : _GEN_111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_113 = 8'h61 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_97 : _GEN_112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_114 = 8'h62 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_98 : _GEN_113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_115 = 8'h63 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_99 : _GEN_114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_116 = 8'h64 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_100 : _GEN_115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_117 = 8'h65 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_101 : _GEN_116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_118 = 8'h66 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_102 : _GEN_117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_119 = 8'h67 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_103 : _GEN_118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_120 = 8'h68 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_104 : _GEN_119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_121 = 8'h69 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_105 : _GEN_120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_122 = 8'h6a == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_106 : _GEN_121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_123 = 8'h6b == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_107 : _GEN_122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_124 = 8'h6c == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_108 : _GEN_123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_125 = 8'h6d == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_109 : _GEN_124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_126 = 8'h6e == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_110 : _GEN_125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_127 = 8'h6f == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_111 : _GEN_126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_128 = 8'h70 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_112 : _GEN_127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_129 = 8'h71 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_113 : _GEN_128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_130 = 8'h72 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_114 : _GEN_129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_131 = 8'h73 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_115 : _GEN_130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_132 = 8'h74 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_116 : _GEN_131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_133 = 8'h75 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_117 : _GEN_132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_134 = 8'h76 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_118 : _GEN_133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_135 = 8'h77 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_119 : _GEN_134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_136 = 8'h78 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_120 : _GEN_135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_137 = 8'h79 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_121 : _GEN_136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_138 = 8'h7a == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_122 : _GEN_137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_139 = 8'h7b == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_123 : _GEN_138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_140 = 8'h7c == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_124 : _GEN_139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_141 = 8'h7d == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_125 : _GEN_140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_142 = 8'h7e == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_126 : _GEN_141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_143 = 8'h7f == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_127 : _GEN_142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_144 = 8'h80 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_128 : _GEN_143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_145 = 8'h81 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_129 : _GEN_144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_146 = 8'h82 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_130 : _GEN_145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_147 = 8'h83 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_131 : _GEN_146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_148 = 8'h84 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_132 : _GEN_147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_149 = 8'h85 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_133 : _GEN_148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_150 = 8'h86 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_134 : _GEN_149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_151 = 8'h87 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_135 : _GEN_150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_152 = 8'h88 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_136 : _GEN_151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_153 = 8'h89 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_137 : _GEN_152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_154 = 8'h8a == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_138 : _GEN_153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_155 = 8'h8b == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_139 : _GEN_154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_156 = 8'h8c == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_140 : _GEN_155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_157 = 8'h8d == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_141 : _GEN_156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_158 = 8'h8e == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_142 : _GEN_157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_159 = 8'h8f == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_143 : _GEN_158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_160 = 8'h90 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_144 : _GEN_159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_161 = 8'h91 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_145 : _GEN_160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_162 = 8'h92 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_146 : _GEN_161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_163 = 8'h93 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_147 : _GEN_162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_164 = 8'h94 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_148 : _GEN_163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_165 = 8'h95 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_149 : _GEN_164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_166 = 8'h96 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_150 : _GEN_165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_167 = 8'h97 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_151 : _GEN_166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_168 = 8'h98 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_152 : _GEN_167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_169 = 8'h99 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_153 : _GEN_168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_170 = 8'h9a == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_154 : _GEN_169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_171 = 8'h9b == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_155 : _GEN_170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_172 = 8'h9c == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_156 : _GEN_171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_173 = 8'h9d == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_157 : _GEN_172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_174 = 8'h9e == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_158 : _GEN_173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_175 = 8'h9f == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_159 : _GEN_174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_176 = 8'ha0 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_160 : _GEN_175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_177 = 8'ha1 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_161 : _GEN_176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_178 = 8'ha2 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_162 : _GEN_177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_179 = 8'ha3 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_163 : _GEN_178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_180 = 8'ha4 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_164 : _GEN_179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_181 = 8'ha5 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_165 : _GEN_180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_182 = 8'ha6 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_166 : _GEN_181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_183 = 8'ha7 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_167 : _GEN_182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_184 = 8'ha8 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_168 : _GEN_183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_185 = 8'ha9 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_169 : _GEN_184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_186 = 8'haa == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_170 : _GEN_185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_187 = 8'hab == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_171 : _GEN_186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_188 = 8'hac == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_172 : _GEN_187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_189 = 8'had == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_173 : _GEN_188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_190 = 8'hae == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_174 : _GEN_189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_191 = 8'haf == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_175 : _GEN_190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_192 = 8'hb0 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_176 : _GEN_191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_193 = 8'hb1 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_177 : _GEN_192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_194 = 8'hb2 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_178 : _GEN_193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_195 = 8'hb3 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_179 : _GEN_194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_196 = 8'hb4 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_180 : _GEN_195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_197 = 8'hb5 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_181 : _GEN_196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_198 = 8'hb6 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_182 : _GEN_197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_199 = 8'hb7 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_183 : _GEN_198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_200 = 8'hb8 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_184 : _GEN_199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_201 = 8'hb9 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_185 : _GEN_200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_202 = 8'hba == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_186 : _GEN_201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_203 = 8'hbb == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_187 : _GEN_202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_204 = 8'hbc == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_188 : _GEN_203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_205 = 8'hbd == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_189 : _GEN_204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_206 = 8'hbe == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_190 : _GEN_205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_207 = 8'hbf == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_191 : _GEN_206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_208 = 8'hc0 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_192 : _GEN_207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_209 = 8'hc1 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_193 : _GEN_208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_210 = 8'hc2 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_194 : _GEN_209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_211 = 8'hc3 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_195 : _GEN_210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_212 = 8'hc4 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_196 : _GEN_211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_213 = 8'hc5 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_197 : _GEN_212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_214 = 8'hc6 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_198 : _GEN_213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_215 = 8'hc7 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_199 : _GEN_214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_216 = 8'hc8 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_200 : _GEN_215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_217 = 8'hc9 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_201 : _GEN_216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_218 = 8'hca == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_202 : _GEN_217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_219 = 8'hcb == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_203 : _GEN_218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_220 = 8'hcc == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_204 : _GEN_219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_221 = 8'hcd == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_205 : _GEN_220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_222 = 8'hce == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_206 : _GEN_221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_223 = 8'hcf == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_207 : _GEN_222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_224 = 8'hd0 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_208 : _GEN_223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_225 = 8'hd1 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_209 : _GEN_224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_226 = 8'hd2 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_210 : _GEN_225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_227 = 8'hd3 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_211 : _GEN_226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_228 = 8'hd4 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_212 : _GEN_227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_229 = 8'hd5 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_213 : _GEN_228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_230 = 8'hd6 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_214 : _GEN_229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_231 = 8'hd7 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_215 : _GEN_230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_232 = 8'hd8 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_216 : _GEN_231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_233 = 8'hd9 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_217 : _GEN_232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_234 = 8'hda == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_218 : _GEN_233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_235 = 8'hdb == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_219 : _GEN_234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_236 = 8'hdc == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_220 : _GEN_235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_237 = 8'hdd == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_221 : _GEN_236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_238 = 8'hde == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_222 : _GEN_237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_239 = 8'hdf == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_223 : _GEN_238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_240 = 8'he0 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_224 : _GEN_239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_241 = 8'he1 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_225 : _GEN_240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_242 = 8'he2 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_226 : _GEN_241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_243 = 8'he3 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_227 : _GEN_242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_244 = 8'he4 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_228 : _GEN_243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_245 = 8'he5 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_229 : _GEN_244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_246 = 8'he6 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_230 : _GEN_245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_247 = 8'he7 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_231 : _GEN_246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_248 = 8'he8 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_232 : _GEN_247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_249 = 8'he9 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_233 : _GEN_248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_250 = 8'hea == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_234 : _GEN_249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_251 = 8'heb == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_235 : _GEN_250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_252 = 8'hec == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_236 : _GEN_251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_253 = 8'hed == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_237 : _GEN_252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_254 = 8'hee == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_238 : _GEN_253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_255 = 8'hef == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_239 : _GEN_254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_256 = 8'hf0 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_240 : _GEN_255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_257 = 8'hf1 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_241 : _GEN_256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_258 = 8'hf2 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_242 : _GEN_257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_259 = 8'hf3 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_243 : _GEN_258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_260 = 8'hf4 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_244 : _GEN_259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_261 = 8'hf5 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_245 : _GEN_260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_262 = 8'hf6 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_246 : _GEN_261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_263 = 8'hf7 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_247 : _GEN_262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_264 = 8'hf8 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_248 : _GEN_263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_265 = 8'hf9 == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_249 : _GEN_264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_266 = 8'hfa == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_250 : _GEN_265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_267 = 8'hfb == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_251 : _GEN_266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_268 = 8'hfc == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_252 : _GEN_267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_269 = 8'hfd == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_253 : _GEN_268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_270 = 8'hfe == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_254 : _GEN_269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_271 = 8'hff == _transition_field_raw_data_T_1 ? io_pipe_phv_in_data_255 : _GEN_270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_273 = 8'h1 == transition_field_offset ? io_pipe_phv_in_data_1 : io_pipe_phv_in_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_274 = 8'h2 == transition_field_offset ? io_pipe_phv_in_data_2 : _GEN_273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_275 = 8'h3 == transition_field_offset ? io_pipe_phv_in_data_3 : _GEN_274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_276 = 8'h4 == transition_field_offset ? io_pipe_phv_in_data_4 : _GEN_275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_277 = 8'h5 == transition_field_offset ? io_pipe_phv_in_data_5 : _GEN_276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_278 = 8'h6 == transition_field_offset ? io_pipe_phv_in_data_6 : _GEN_277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_279 = 8'h7 == transition_field_offset ? io_pipe_phv_in_data_7 : _GEN_278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_280 = 8'h8 == transition_field_offset ? io_pipe_phv_in_data_8 : _GEN_279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_281 = 8'h9 == transition_field_offset ? io_pipe_phv_in_data_9 : _GEN_280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_282 = 8'ha == transition_field_offset ? io_pipe_phv_in_data_10 : _GEN_281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_283 = 8'hb == transition_field_offset ? io_pipe_phv_in_data_11 : _GEN_282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_284 = 8'hc == transition_field_offset ? io_pipe_phv_in_data_12 : _GEN_283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_285 = 8'hd == transition_field_offset ? io_pipe_phv_in_data_13 : _GEN_284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_286 = 8'he == transition_field_offset ? io_pipe_phv_in_data_14 : _GEN_285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_287 = 8'hf == transition_field_offset ? io_pipe_phv_in_data_15 : _GEN_286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_288 = 8'h10 == transition_field_offset ? io_pipe_phv_in_data_16 : _GEN_287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_289 = 8'h11 == transition_field_offset ? io_pipe_phv_in_data_17 : _GEN_288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_290 = 8'h12 == transition_field_offset ? io_pipe_phv_in_data_18 : _GEN_289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_291 = 8'h13 == transition_field_offset ? io_pipe_phv_in_data_19 : _GEN_290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_292 = 8'h14 == transition_field_offset ? io_pipe_phv_in_data_20 : _GEN_291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_293 = 8'h15 == transition_field_offset ? io_pipe_phv_in_data_21 : _GEN_292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_294 = 8'h16 == transition_field_offset ? io_pipe_phv_in_data_22 : _GEN_293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_295 = 8'h17 == transition_field_offset ? io_pipe_phv_in_data_23 : _GEN_294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_296 = 8'h18 == transition_field_offset ? io_pipe_phv_in_data_24 : _GEN_295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_297 = 8'h19 == transition_field_offset ? io_pipe_phv_in_data_25 : _GEN_296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_298 = 8'h1a == transition_field_offset ? io_pipe_phv_in_data_26 : _GEN_297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_299 = 8'h1b == transition_field_offset ? io_pipe_phv_in_data_27 : _GEN_298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_300 = 8'h1c == transition_field_offset ? io_pipe_phv_in_data_28 : _GEN_299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_301 = 8'h1d == transition_field_offset ? io_pipe_phv_in_data_29 : _GEN_300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_302 = 8'h1e == transition_field_offset ? io_pipe_phv_in_data_30 : _GEN_301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_303 = 8'h1f == transition_field_offset ? io_pipe_phv_in_data_31 : _GEN_302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_304 = 8'h20 == transition_field_offset ? io_pipe_phv_in_data_32 : _GEN_303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_305 = 8'h21 == transition_field_offset ? io_pipe_phv_in_data_33 : _GEN_304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_306 = 8'h22 == transition_field_offset ? io_pipe_phv_in_data_34 : _GEN_305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_307 = 8'h23 == transition_field_offset ? io_pipe_phv_in_data_35 : _GEN_306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_308 = 8'h24 == transition_field_offset ? io_pipe_phv_in_data_36 : _GEN_307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_309 = 8'h25 == transition_field_offset ? io_pipe_phv_in_data_37 : _GEN_308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_310 = 8'h26 == transition_field_offset ? io_pipe_phv_in_data_38 : _GEN_309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_311 = 8'h27 == transition_field_offset ? io_pipe_phv_in_data_39 : _GEN_310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_312 = 8'h28 == transition_field_offset ? io_pipe_phv_in_data_40 : _GEN_311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_313 = 8'h29 == transition_field_offset ? io_pipe_phv_in_data_41 : _GEN_312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_314 = 8'h2a == transition_field_offset ? io_pipe_phv_in_data_42 : _GEN_313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_315 = 8'h2b == transition_field_offset ? io_pipe_phv_in_data_43 : _GEN_314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_316 = 8'h2c == transition_field_offset ? io_pipe_phv_in_data_44 : _GEN_315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_317 = 8'h2d == transition_field_offset ? io_pipe_phv_in_data_45 : _GEN_316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_318 = 8'h2e == transition_field_offset ? io_pipe_phv_in_data_46 : _GEN_317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_319 = 8'h2f == transition_field_offset ? io_pipe_phv_in_data_47 : _GEN_318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_320 = 8'h30 == transition_field_offset ? io_pipe_phv_in_data_48 : _GEN_319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_321 = 8'h31 == transition_field_offset ? io_pipe_phv_in_data_49 : _GEN_320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_322 = 8'h32 == transition_field_offset ? io_pipe_phv_in_data_50 : _GEN_321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_323 = 8'h33 == transition_field_offset ? io_pipe_phv_in_data_51 : _GEN_322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_324 = 8'h34 == transition_field_offset ? io_pipe_phv_in_data_52 : _GEN_323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_325 = 8'h35 == transition_field_offset ? io_pipe_phv_in_data_53 : _GEN_324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_326 = 8'h36 == transition_field_offset ? io_pipe_phv_in_data_54 : _GEN_325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_327 = 8'h37 == transition_field_offset ? io_pipe_phv_in_data_55 : _GEN_326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_328 = 8'h38 == transition_field_offset ? io_pipe_phv_in_data_56 : _GEN_327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_329 = 8'h39 == transition_field_offset ? io_pipe_phv_in_data_57 : _GEN_328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_330 = 8'h3a == transition_field_offset ? io_pipe_phv_in_data_58 : _GEN_329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_331 = 8'h3b == transition_field_offset ? io_pipe_phv_in_data_59 : _GEN_330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_332 = 8'h3c == transition_field_offset ? io_pipe_phv_in_data_60 : _GEN_331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_333 = 8'h3d == transition_field_offset ? io_pipe_phv_in_data_61 : _GEN_332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_334 = 8'h3e == transition_field_offset ? io_pipe_phv_in_data_62 : _GEN_333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_335 = 8'h3f == transition_field_offset ? io_pipe_phv_in_data_63 : _GEN_334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_336 = 8'h40 == transition_field_offset ? io_pipe_phv_in_data_64 : _GEN_335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_337 = 8'h41 == transition_field_offset ? io_pipe_phv_in_data_65 : _GEN_336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_338 = 8'h42 == transition_field_offset ? io_pipe_phv_in_data_66 : _GEN_337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_339 = 8'h43 == transition_field_offset ? io_pipe_phv_in_data_67 : _GEN_338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_340 = 8'h44 == transition_field_offset ? io_pipe_phv_in_data_68 : _GEN_339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_341 = 8'h45 == transition_field_offset ? io_pipe_phv_in_data_69 : _GEN_340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_342 = 8'h46 == transition_field_offset ? io_pipe_phv_in_data_70 : _GEN_341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_343 = 8'h47 == transition_field_offset ? io_pipe_phv_in_data_71 : _GEN_342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_344 = 8'h48 == transition_field_offset ? io_pipe_phv_in_data_72 : _GEN_343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_345 = 8'h49 == transition_field_offset ? io_pipe_phv_in_data_73 : _GEN_344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_346 = 8'h4a == transition_field_offset ? io_pipe_phv_in_data_74 : _GEN_345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_347 = 8'h4b == transition_field_offset ? io_pipe_phv_in_data_75 : _GEN_346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_348 = 8'h4c == transition_field_offset ? io_pipe_phv_in_data_76 : _GEN_347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_349 = 8'h4d == transition_field_offset ? io_pipe_phv_in_data_77 : _GEN_348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_350 = 8'h4e == transition_field_offset ? io_pipe_phv_in_data_78 : _GEN_349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_351 = 8'h4f == transition_field_offset ? io_pipe_phv_in_data_79 : _GEN_350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_352 = 8'h50 == transition_field_offset ? io_pipe_phv_in_data_80 : _GEN_351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_353 = 8'h51 == transition_field_offset ? io_pipe_phv_in_data_81 : _GEN_352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_354 = 8'h52 == transition_field_offset ? io_pipe_phv_in_data_82 : _GEN_353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_355 = 8'h53 == transition_field_offset ? io_pipe_phv_in_data_83 : _GEN_354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_356 = 8'h54 == transition_field_offset ? io_pipe_phv_in_data_84 : _GEN_355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_357 = 8'h55 == transition_field_offset ? io_pipe_phv_in_data_85 : _GEN_356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_358 = 8'h56 == transition_field_offset ? io_pipe_phv_in_data_86 : _GEN_357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_359 = 8'h57 == transition_field_offset ? io_pipe_phv_in_data_87 : _GEN_358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_360 = 8'h58 == transition_field_offset ? io_pipe_phv_in_data_88 : _GEN_359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_361 = 8'h59 == transition_field_offset ? io_pipe_phv_in_data_89 : _GEN_360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_362 = 8'h5a == transition_field_offset ? io_pipe_phv_in_data_90 : _GEN_361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_363 = 8'h5b == transition_field_offset ? io_pipe_phv_in_data_91 : _GEN_362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_364 = 8'h5c == transition_field_offset ? io_pipe_phv_in_data_92 : _GEN_363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_365 = 8'h5d == transition_field_offset ? io_pipe_phv_in_data_93 : _GEN_364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_366 = 8'h5e == transition_field_offset ? io_pipe_phv_in_data_94 : _GEN_365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_367 = 8'h5f == transition_field_offset ? io_pipe_phv_in_data_95 : _GEN_366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_368 = 8'h60 == transition_field_offset ? io_pipe_phv_in_data_96 : _GEN_367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_369 = 8'h61 == transition_field_offset ? io_pipe_phv_in_data_97 : _GEN_368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_370 = 8'h62 == transition_field_offset ? io_pipe_phv_in_data_98 : _GEN_369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_371 = 8'h63 == transition_field_offset ? io_pipe_phv_in_data_99 : _GEN_370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_372 = 8'h64 == transition_field_offset ? io_pipe_phv_in_data_100 : _GEN_371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_373 = 8'h65 == transition_field_offset ? io_pipe_phv_in_data_101 : _GEN_372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_374 = 8'h66 == transition_field_offset ? io_pipe_phv_in_data_102 : _GEN_373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_375 = 8'h67 == transition_field_offset ? io_pipe_phv_in_data_103 : _GEN_374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_376 = 8'h68 == transition_field_offset ? io_pipe_phv_in_data_104 : _GEN_375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_377 = 8'h69 == transition_field_offset ? io_pipe_phv_in_data_105 : _GEN_376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_378 = 8'h6a == transition_field_offset ? io_pipe_phv_in_data_106 : _GEN_377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_379 = 8'h6b == transition_field_offset ? io_pipe_phv_in_data_107 : _GEN_378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_380 = 8'h6c == transition_field_offset ? io_pipe_phv_in_data_108 : _GEN_379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_381 = 8'h6d == transition_field_offset ? io_pipe_phv_in_data_109 : _GEN_380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_382 = 8'h6e == transition_field_offset ? io_pipe_phv_in_data_110 : _GEN_381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_383 = 8'h6f == transition_field_offset ? io_pipe_phv_in_data_111 : _GEN_382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_384 = 8'h70 == transition_field_offset ? io_pipe_phv_in_data_112 : _GEN_383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_385 = 8'h71 == transition_field_offset ? io_pipe_phv_in_data_113 : _GEN_384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_386 = 8'h72 == transition_field_offset ? io_pipe_phv_in_data_114 : _GEN_385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_387 = 8'h73 == transition_field_offset ? io_pipe_phv_in_data_115 : _GEN_386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_388 = 8'h74 == transition_field_offset ? io_pipe_phv_in_data_116 : _GEN_387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_389 = 8'h75 == transition_field_offset ? io_pipe_phv_in_data_117 : _GEN_388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_390 = 8'h76 == transition_field_offset ? io_pipe_phv_in_data_118 : _GEN_389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_391 = 8'h77 == transition_field_offset ? io_pipe_phv_in_data_119 : _GEN_390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_392 = 8'h78 == transition_field_offset ? io_pipe_phv_in_data_120 : _GEN_391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_393 = 8'h79 == transition_field_offset ? io_pipe_phv_in_data_121 : _GEN_392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_394 = 8'h7a == transition_field_offset ? io_pipe_phv_in_data_122 : _GEN_393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_395 = 8'h7b == transition_field_offset ? io_pipe_phv_in_data_123 : _GEN_394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_396 = 8'h7c == transition_field_offset ? io_pipe_phv_in_data_124 : _GEN_395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_397 = 8'h7d == transition_field_offset ? io_pipe_phv_in_data_125 : _GEN_396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_398 = 8'h7e == transition_field_offset ? io_pipe_phv_in_data_126 : _GEN_397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_399 = 8'h7f == transition_field_offset ? io_pipe_phv_in_data_127 : _GEN_398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_400 = 8'h80 == transition_field_offset ? io_pipe_phv_in_data_128 : _GEN_399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_401 = 8'h81 == transition_field_offset ? io_pipe_phv_in_data_129 : _GEN_400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_402 = 8'h82 == transition_field_offset ? io_pipe_phv_in_data_130 : _GEN_401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_403 = 8'h83 == transition_field_offset ? io_pipe_phv_in_data_131 : _GEN_402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_404 = 8'h84 == transition_field_offset ? io_pipe_phv_in_data_132 : _GEN_403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_405 = 8'h85 == transition_field_offset ? io_pipe_phv_in_data_133 : _GEN_404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_406 = 8'h86 == transition_field_offset ? io_pipe_phv_in_data_134 : _GEN_405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_407 = 8'h87 == transition_field_offset ? io_pipe_phv_in_data_135 : _GEN_406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_408 = 8'h88 == transition_field_offset ? io_pipe_phv_in_data_136 : _GEN_407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_409 = 8'h89 == transition_field_offset ? io_pipe_phv_in_data_137 : _GEN_408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_410 = 8'h8a == transition_field_offset ? io_pipe_phv_in_data_138 : _GEN_409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_411 = 8'h8b == transition_field_offset ? io_pipe_phv_in_data_139 : _GEN_410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_412 = 8'h8c == transition_field_offset ? io_pipe_phv_in_data_140 : _GEN_411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_413 = 8'h8d == transition_field_offset ? io_pipe_phv_in_data_141 : _GEN_412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_414 = 8'h8e == transition_field_offset ? io_pipe_phv_in_data_142 : _GEN_413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_415 = 8'h8f == transition_field_offset ? io_pipe_phv_in_data_143 : _GEN_414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_416 = 8'h90 == transition_field_offset ? io_pipe_phv_in_data_144 : _GEN_415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_417 = 8'h91 == transition_field_offset ? io_pipe_phv_in_data_145 : _GEN_416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_418 = 8'h92 == transition_field_offset ? io_pipe_phv_in_data_146 : _GEN_417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_419 = 8'h93 == transition_field_offset ? io_pipe_phv_in_data_147 : _GEN_418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_420 = 8'h94 == transition_field_offset ? io_pipe_phv_in_data_148 : _GEN_419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_421 = 8'h95 == transition_field_offset ? io_pipe_phv_in_data_149 : _GEN_420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_422 = 8'h96 == transition_field_offset ? io_pipe_phv_in_data_150 : _GEN_421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_423 = 8'h97 == transition_field_offset ? io_pipe_phv_in_data_151 : _GEN_422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_424 = 8'h98 == transition_field_offset ? io_pipe_phv_in_data_152 : _GEN_423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_425 = 8'h99 == transition_field_offset ? io_pipe_phv_in_data_153 : _GEN_424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_426 = 8'h9a == transition_field_offset ? io_pipe_phv_in_data_154 : _GEN_425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_427 = 8'h9b == transition_field_offset ? io_pipe_phv_in_data_155 : _GEN_426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_428 = 8'h9c == transition_field_offset ? io_pipe_phv_in_data_156 : _GEN_427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_429 = 8'h9d == transition_field_offset ? io_pipe_phv_in_data_157 : _GEN_428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_430 = 8'h9e == transition_field_offset ? io_pipe_phv_in_data_158 : _GEN_429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_431 = 8'h9f == transition_field_offset ? io_pipe_phv_in_data_159 : _GEN_430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_432 = 8'ha0 == transition_field_offset ? io_pipe_phv_in_data_160 : _GEN_431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_433 = 8'ha1 == transition_field_offset ? io_pipe_phv_in_data_161 : _GEN_432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_434 = 8'ha2 == transition_field_offset ? io_pipe_phv_in_data_162 : _GEN_433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_435 = 8'ha3 == transition_field_offset ? io_pipe_phv_in_data_163 : _GEN_434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_436 = 8'ha4 == transition_field_offset ? io_pipe_phv_in_data_164 : _GEN_435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_437 = 8'ha5 == transition_field_offset ? io_pipe_phv_in_data_165 : _GEN_436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_438 = 8'ha6 == transition_field_offset ? io_pipe_phv_in_data_166 : _GEN_437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_439 = 8'ha7 == transition_field_offset ? io_pipe_phv_in_data_167 : _GEN_438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_440 = 8'ha8 == transition_field_offset ? io_pipe_phv_in_data_168 : _GEN_439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_441 = 8'ha9 == transition_field_offset ? io_pipe_phv_in_data_169 : _GEN_440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_442 = 8'haa == transition_field_offset ? io_pipe_phv_in_data_170 : _GEN_441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_443 = 8'hab == transition_field_offset ? io_pipe_phv_in_data_171 : _GEN_442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_444 = 8'hac == transition_field_offset ? io_pipe_phv_in_data_172 : _GEN_443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_445 = 8'had == transition_field_offset ? io_pipe_phv_in_data_173 : _GEN_444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_446 = 8'hae == transition_field_offset ? io_pipe_phv_in_data_174 : _GEN_445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_447 = 8'haf == transition_field_offset ? io_pipe_phv_in_data_175 : _GEN_446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_448 = 8'hb0 == transition_field_offset ? io_pipe_phv_in_data_176 : _GEN_447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_449 = 8'hb1 == transition_field_offset ? io_pipe_phv_in_data_177 : _GEN_448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_450 = 8'hb2 == transition_field_offset ? io_pipe_phv_in_data_178 : _GEN_449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_451 = 8'hb3 == transition_field_offset ? io_pipe_phv_in_data_179 : _GEN_450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_452 = 8'hb4 == transition_field_offset ? io_pipe_phv_in_data_180 : _GEN_451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_453 = 8'hb5 == transition_field_offset ? io_pipe_phv_in_data_181 : _GEN_452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_454 = 8'hb6 == transition_field_offset ? io_pipe_phv_in_data_182 : _GEN_453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_455 = 8'hb7 == transition_field_offset ? io_pipe_phv_in_data_183 : _GEN_454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_456 = 8'hb8 == transition_field_offset ? io_pipe_phv_in_data_184 : _GEN_455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_457 = 8'hb9 == transition_field_offset ? io_pipe_phv_in_data_185 : _GEN_456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_458 = 8'hba == transition_field_offset ? io_pipe_phv_in_data_186 : _GEN_457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_459 = 8'hbb == transition_field_offset ? io_pipe_phv_in_data_187 : _GEN_458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_460 = 8'hbc == transition_field_offset ? io_pipe_phv_in_data_188 : _GEN_459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_461 = 8'hbd == transition_field_offset ? io_pipe_phv_in_data_189 : _GEN_460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_462 = 8'hbe == transition_field_offset ? io_pipe_phv_in_data_190 : _GEN_461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_463 = 8'hbf == transition_field_offset ? io_pipe_phv_in_data_191 : _GEN_462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_464 = 8'hc0 == transition_field_offset ? io_pipe_phv_in_data_192 : _GEN_463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_465 = 8'hc1 == transition_field_offset ? io_pipe_phv_in_data_193 : _GEN_464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_466 = 8'hc2 == transition_field_offset ? io_pipe_phv_in_data_194 : _GEN_465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_467 = 8'hc3 == transition_field_offset ? io_pipe_phv_in_data_195 : _GEN_466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_468 = 8'hc4 == transition_field_offset ? io_pipe_phv_in_data_196 : _GEN_467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_469 = 8'hc5 == transition_field_offset ? io_pipe_phv_in_data_197 : _GEN_468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_470 = 8'hc6 == transition_field_offset ? io_pipe_phv_in_data_198 : _GEN_469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_471 = 8'hc7 == transition_field_offset ? io_pipe_phv_in_data_199 : _GEN_470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_472 = 8'hc8 == transition_field_offset ? io_pipe_phv_in_data_200 : _GEN_471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_473 = 8'hc9 == transition_field_offset ? io_pipe_phv_in_data_201 : _GEN_472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_474 = 8'hca == transition_field_offset ? io_pipe_phv_in_data_202 : _GEN_473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_475 = 8'hcb == transition_field_offset ? io_pipe_phv_in_data_203 : _GEN_474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_476 = 8'hcc == transition_field_offset ? io_pipe_phv_in_data_204 : _GEN_475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_477 = 8'hcd == transition_field_offset ? io_pipe_phv_in_data_205 : _GEN_476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_478 = 8'hce == transition_field_offset ? io_pipe_phv_in_data_206 : _GEN_477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_479 = 8'hcf == transition_field_offset ? io_pipe_phv_in_data_207 : _GEN_478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_480 = 8'hd0 == transition_field_offset ? io_pipe_phv_in_data_208 : _GEN_479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_481 = 8'hd1 == transition_field_offset ? io_pipe_phv_in_data_209 : _GEN_480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_482 = 8'hd2 == transition_field_offset ? io_pipe_phv_in_data_210 : _GEN_481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_483 = 8'hd3 == transition_field_offset ? io_pipe_phv_in_data_211 : _GEN_482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_484 = 8'hd4 == transition_field_offset ? io_pipe_phv_in_data_212 : _GEN_483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_485 = 8'hd5 == transition_field_offset ? io_pipe_phv_in_data_213 : _GEN_484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_486 = 8'hd6 == transition_field_offset ? io_pipe_phv_in_data_214 : _GEN_485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_487 = 8'hd7 == transition_field_offset ? io_pipe_phv_in_data_215 : _GEN_486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_488 = 8'hd8 == transition_field_offset ? io_pipe_phv_in_data_216 : _GEN_487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_489 = 8'hd9 == transition_field_offset ? io_pipe_phv_in_data_217 : _GEN_488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_490 = 8'hda == transition_field_offset ? io_pipe_phv_in_data_218 : _GEN_489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_491 = 8'hdb == transition_field_offset ? io_pipe_phv_in_data_219 : _GEN_490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_492 = 8'hdc == transition_field_offset ? io_pipe_phv_in_data_220 : _GEN_491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_493 = 8'hdd == transition_field_offset ? io_pipe_phv_in_data_221 : _GEN_492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_494 = 8'hde == transition_field_offset ? io_pipe_phv_in_data_222 : _GEN_493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_495 = 8'hdf == transition_field_offset ? io_pipe_phv_in_data_223 : _GEN_494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_496 = 8'he0 == transition_field_offset ? io_pipe_phv_in_data_224 : _GEN_495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_497 = 8'he1 == transition_field_offset ? io_pipe_phv_in_data_225 : _GEN_496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_498 = 8'he2 == transition_field_offset ? io_pipe_phv_in_data_226 : _GEN_497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_499 = 8'he3 == transition_field_offset ? io_pipe_phv_in_data_227 : _GEN_498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_500 = 8'he4 == transition_field_offset ? io_pipe_phv_in_data_228 : _GEN_499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_501 = 8'he5 == transition_field_offset ? io_pipe_phv_in_data_229 : _GEN_500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_502 = 8'he6 == transition_field_offset ? io_pipe_phv_in_data_230 : _GEN_501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_503 = 8'he7 == transition_field_offset ? io_pipe_phv_in_data_231 : _GEN_502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_504 = 8'he8 == transition_field_offset ? io_pipe_phv_in_data_232 : _GEN_503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_505 = 8'he9 == transition_field_offset ? io_pipe_phv_in_data_233 : _GEN_504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_506 = 8'hea == transition_field_offset ? io_pipe_phv_in_data_234 : _GEN_505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_507 = 8'heb == transition_field_offset ? io_pipe_phv_in_data_235 : _GEN_506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_508 = 8'hec == transition_field_offset ? io_pipe_phv_in_data_236 : _GEN_507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_509 = 8'hed == transition_field_offset ? io_pipe_phv_in_data_237 : _GEN_508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_510 = 8'hee == transition_field_offset ? io_pipe_phv_in_data_238 : _GEN_509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_511 = 8'hef == transition_field_offset ? io_pipe_phv_in_data_239 : _GEN_510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_512 = 8'hf0 == transition_field_offset ? io_pipe_phv_in_data_240 : _GEN_511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_513 = 8'hf1 == transition_field_offset ? io_pipe_phv_in_data_241 : _GEN_512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_514 = 8'hf2 == transition_field_offset ? io_pipe_phv_in_data_242 : _GEN_513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_515 = 8'hf3 == transition_field_offset ? io_pipe_phv_in_data_243 : _GEN_514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_516 = 8'hf4 == transition_field_offset ? io_pipe_phv_in_data_244 : _GEN_515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_517 = 8'hf5 == transition_field_offset ? io_pipe_phv_in_data_245 : _GEN_516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_518 = 8'hf6 == transition_field_offset ? io_pipe_phv_in_data_246 : _GEN_517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_519 = 8'hf7 == transition_field_offset ? io_pipe_phv_in_data_247 : _GEN_518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_520 = 8'hf8 == transition_field_offset ? io_pipe_phv_in_data_248 : _GEN_519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_521 = 8'hf9 == transition_field_offset ? io_pipe_phv_in_data_249 : _GEN_520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_522 = 8'hfa == transition_field_offset ? io_pipe_phv_in_data_250 : _GEN_521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_523 = 8'hfb == transition_field_offset ? io_pipe_phv_in_data_251 : _GEN_522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_524 = 8'hfc == transition_field_offset ? io_pipe_phv_in_data_252 : _GEN_523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_525 = 8'hfd == transition_field_offset ? io_pipe_phv_in_data_253 : _GEN_524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_526 = 8'hfe == transition_field_offset ? io_pipe_phv_in_data_254 : _GEN_525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_527 = 8'hff == transition_field_offset ? io_pipe_phv_in_data_255 : _GEN_526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [15:0] transition_field_raw_data = {_GEN_271,_GEN_527}; // @[Cat.scala 30:58]
  wire [15:0] transition_field = transition_field_raw_data ^ match_val_transition_field_mask; // @[parse_module.scala 76:58]
  wire [15:0] _phv_header_T = {io_pipe_phv_in_parse_current_offset,phv_header_lo}; // @[Cat.scala 30:58]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_96 = phv_data_96; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_97 = phv_data_97; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_98 = phv_data_98; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_99 = phv_data_99; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_100 = phv_data_100; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_101 = phv_data_101; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_102 = phv_data_102; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_103 = phv_data_103; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_104 = phv_data_104; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_105 = phv_data_105; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_106 = phv_data_106; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_107 = phv_data_107; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_108 = phv_data_108; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_109 = phv_data_109; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_110 = phv_data_110; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_111 = phv_data_111; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_112 = phv_data_112; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_113 = phv_data_113; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_114 = phv_data_114; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_115 = phv_data_115; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_116 = phv_data_116; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_117 = phv_data_117; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_118 = phv_data_118; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_119 = phv_data_119; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_120 = phv_data_120; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_121 = phv_data_121; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_122 = phv_data_122; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_123 = phv_data_123; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_124 = phv_data_124; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_125 = phv_data_125; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_126 = phv_data_126; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_127 = phv_data_127; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_128 = phv_data_128; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_129 = phv_data_129; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_130 = phv_data_130; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_131 = phv_data_131; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_132 = phv_data_132; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_133 = phv_data_133; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_134 = phv_data_134; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_135 = phv_data_135; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_136 = phv_data_136; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_137 = phv_data_137; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_138 = phv_data_138; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_139 = phv_data_139; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_140 = phv_data_140; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_141 = phv_data_141; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_142 = phv_data_142; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_143 = phv_data_143; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_144 = phv_data_144; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_145 = phv_data_145; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_146 = phv_data_146; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_147 = phv_data_147; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_148 = phv_data_148; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_149 = phv_data_149; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_150 = phv_data_150; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_151 = phv_data_151; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_152 = phv_data_152; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_153 = phv_data_153; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_154 = phv_data_154; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_155 = phv_data_155; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_156 = phv_data_156; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_157 = phv_data_157; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_158 = phv_data_158; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_159 = phv_data_159; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_160 = phv_data_160; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_161 = phv_data_161; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_162 = phv_data_162; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_163 = phv_data_163; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_164 = phv_data_164; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_165 = phv_data_165; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_166 = phv_data_166; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_167 = phv_data_167; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_168 = phv_data_168; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_169 = phv_data_169; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_170 = phv_data_170; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_171 = phv_data_171; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_172 = phv_data_172; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_173 = phv_data_173; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_174 = phv_data_174; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_175 = phv_data_175; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_176 = phv_data_176; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_177 = phv_data_177; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_178 = phv_data_178; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_179 = phv_data_179; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_180 = phv_data_180; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_181 = phv_data_181; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_182 = phv_data_182; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_183 = phv_data_183; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_184 = phv_data_184; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_185 = phv_data_185; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_186 = phv_data_186; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_187 = phv_data_187; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_188 = phv_data_188; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_189 = phv_data_189; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_190 = phv_data_190; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_191 = phv_data_191; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_192 = phv_data_192; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_193 = phv_data_193; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_194 = phv_data_194; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_195 = phv_data_195; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_196 = phv_data_196; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_197 = phv_data_197; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_198 = phv_data_198; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_199 = phv_data_199; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_200 = phv_data_200; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_201 = phv_data_201; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_202 = phv_data_202; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_203 = phv_data_203; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_204 = phv_data_204; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_205 = phv_data_205; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_206 = phv_data_206; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_207 = phv_data_207; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_208 = phv_data_208; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_209 = phv_data_209; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_210 = phv_data_210; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_211 = phv_data_211; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_212 = phv_data_212; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_213 = phv_data_213; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_214 = phv_data_214; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_215 = phv_data_215; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_216 = phv_data_216; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_217 = phv_data_217; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_218 = phv_data_218; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_219 = phv_data_219; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_220 = phv_data_220; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_221 = phv_data_221; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_222 = phv_data_222; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_223 = phv_data_223; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_224 = phv_data_224; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_225 = phv_data_225; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_226 = phv_data_226; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_227 = phv_data_227; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_228 = phv_data_228; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_229 = phv_data_229; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_230 = phv_data_230; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_231 = phv_data_231; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_232 = phv_data_232; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_233 = phv_data_233; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_234 = phv_data_234; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_235 = phv_data_235; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_236 = phv_data_236; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_237 = phv_data_237; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_238 = phv_data_238; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_239 = phv_data_239; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_240 = phv_data_240; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_241 = phv_data_241; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_242 = phv_data_242; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_243 = phv_data_243; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_244 = phv_data_244; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_245 = phv_data_245; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_246 = phv_data_246; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_247 = phv_data_247; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_248 = phv_data_248; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_249 = phv_data_249; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_250 = phv_data_250; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_251 = phv_data_251; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_252 = phv_data_252; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_253 = phv_data_253; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_254 = phv_data_254; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_data_255 = phv_data_255; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[parse_module.scala 52:21]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[parse_module.scala 52:21]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[parse_module.scala 51:9]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[parse_module.scala 51:9]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[parse_module.scala 51:9]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[parse_module.scala 51:9]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[parse_module.scala 51:9]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[parse_module.scala 51:9]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[parse_module.scala 51:9]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[parse_module.scala 51:9]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[parse_module.scala 51:9]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[parse_module.scala 51:9]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[parse_module.scala 51:9]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[parse_module.scala 51:9]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[parse_module.scala 51:9]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[parse_module.scala 51:9]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[parse_module.scala 51:9]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[parse_module.scala 51:9]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[parse_module.scala 51:9]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[parse_module.scala 51:9]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[parse_module.scala 51:9]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[parse_module.scala 51:9]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[parse_module.scala 51:9]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[parse_module.scala 51:9]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[parse_module.scala 51:9]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[parse_module.scala 51:9]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[parse_module.scala 51:9]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[parse_module.scala 51:9]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[parse_module.scala 51:9]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[parse_module.scala 51:9]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[parse_module.scala 51:9]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[parse_module.scala 51:9]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[parse_module.scala 51:9]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[parse_module.scala 51:9]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[parse_module.scala 51:9]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[parse_module.scala 51:9]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[parse_module.scala 51:9]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[parse_module.scala 51:9]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[parse_module.scala 51:9]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[parse_module.scala 51:9]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[parse_module.scala 51:9]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[parse_module.scala 51:9]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[parse_module.scala 51:9]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[parse_module.scala 51:9]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[parse_module.scala 51:9]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[parse_module.scala 51:9]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[parse_module.scala 51:9]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[parse_module.scala 51:9]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[parse_module.scala 51:9]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[parse_module.scala 51:9]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[parse_module.scala 51:9]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[parse_module.scala 51:9]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[parse_module.scala 51:9]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[parse_module.scala 51:9]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[parse_module.scala 51:9]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[parse_module.scala 51:9]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[parse_module.scala 51:9]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[parse_module.scala 51:9]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[parse_module.scala 51:9]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[parse_module.scala 51:9]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[parse_module.scala 51:9]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[parse_module.scala 51:9]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[parse_module.scala 51:9]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[parse_module.scala 51:9]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[parse_module.scala 51:9]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[parse_module.scala 51:9]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[parse_module.scala 51:9]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[parse_module.scala 51:9]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[parse_module.scala 51:9]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[parse_module.scala 51:9]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[parse_module.scala 51:9]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[parse_module.scala 51:9]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[parse_module.scala 51:9]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[parse_module.scala 51:9]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[parse_module.scala 51:9]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[parse_module.scala 51:9]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[parse_module.scala 51:9]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[parse_module.scala 51:9]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[parse_module.scala 51:9]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[parse_module.scala 51:9]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[parse_module.scala 51:9]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[parse_module.scala 51:9]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[parse_module.scala 51:9]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[parse_module.scala 51:9]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[parse_module.scala 51:9]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[parse_module.scala 51:9]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[parse_module.scala 51:9]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[parse_module.scala 51:9]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[parse_module.scala 51:9]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[parse_module.scala 51:9]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[parse_module.scala 51:9]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[parse_module.scala 51:9]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[parse_module.scala 51:9]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[parse_module.scala 51:9]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[parse_module.scala 51:9]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[parse_module.scala 51:9]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[parse_module.scala 51:9]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[parse_module.scala 51:9]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[parse_module.scala 51:9]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[parse_module.scala 51:9]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[parse_module.scala 51:9]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[parse_module.scala 51:9]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[parse_module.scala 51:9]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[parse_module.scala 51:9]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[parse_module.scala 51:9]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[parse_module.scala 51:9]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[parse_module.scala 51:9]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[parse_module.scala 51:9]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[parse_module.scala 51:9]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[parse_module.scala 51:9]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[parse_module.scala 51:9]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[parse_module.scala 51:9]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[parse_module.scala 51:9]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[parse_module.scala 51:9]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[parse_module.scala 51:9]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[parse_module.scala 51:9]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[parse_module.scala 51:9]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[parse_module.scala 51:9]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[parse_module.scala 51:9]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[parse_module.scala 51:9]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[parse_module.scala 51:9]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[parse_module.scala 51:9]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[parse_module.scala 51:9]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[parse_module.scala 51:9]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[parse_module.scala 51:9]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[parse_module.scala 51:9]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[parse_module.scala 51:9]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[parse_module.scala 51:9]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[parse_module.scala 51:9]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[parse_module.scala 51:9]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[parse_module.scala 51:9]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[parse_module.scala 51:9]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[parse_module.scala 51:9]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[parse_module.scala 51:9]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[parse_module.scala 51:9]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[parse_module.scala 51:9]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[parse_module.scala 51:9]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[parse_module.scala 51:9]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[parse_module.scala 51:9]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[parse_module.scala 51:9]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[parse_module.scala 51:9]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[parse_module.scala 51:9]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[parse_module.scala 51:9]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[parse_module.scala 51:9]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[parse_module.scala 51:9]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[parse_module.scala 51:9]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[parse_module.scala 51:9]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[parse_module.scala 51:9]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[parse_module.scala 51:9]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[parse_module.scala 51:9]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[parse_module.scala 51:9]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[parse_module.scala 51:9]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[parse_module.scala 51:9]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[parse_module.scala 51:9]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[parse_module.scala 51:9]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[parse_module.scala 51:9]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[parse_module.scala 51:9]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[parse_module.scala 51:9]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[parse_module.scala 51:9]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[parse_module.scala 51:9]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[parse_module.scala 51:9]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[parse_module.scala 51:9]
    phv_data_160 <= io_pipe_phv_in_data_160; // @[parse_module.scala 51:9]
    phv_data_161 <= io_pipe_phv_in_data_161; // @[parse_module.scala 51:9]
    phv_data_162 <= io_pipe_phv_in_data_162; // @[parse_module.scala 51:9]
    phv_data_163 <= io_pipe_phv_in_data_163; // @[parse_module.scala 51:9]
    phv_data_164 <= io_pipe_phv_in_data_164; // @[parse_module.scala 51:9]
    phv_data_165 <= io_pipe_phv_in_data_165; // @[parse_module.scala 51:9]
    phv_data_166 <= io_pipe_phv_in_data_166; // @[parse_module.scala 51:9]
    phv_data_167 <= io_pipe_phv_in_data_167; // @[parse_module.scala 51:9]
    phv_data_168 <= io_pipe_phv_in_data_168; // @[parse_module.scala 51:9]
    phv_data_169 <= io_pipe_phv_in_data_169; // @[parse_module.scala 51:9]
    phv_data_170 <= io_pipe_phv_in_data_170; // @[parse_module.scala 51:9]
    phv_data_171 <= io_pipe_phv_in_data_171; // @[parse_module.scala 51:9]
    phv_data_172 <= io_pipe_phv_in_data_172; // @[parse_module.scala 51:9]
    phv_data_173 <= io_pipe_phv_in_data_173; // @[parse_module.scala 51:9]
    phv_data_174 <= io_pipe_phv_in_data_174; // @[parse_module.scala 51:9]
    phv_data_175 <= io_pipe_phv_in_data_175; // @[parse_module.scala 51:9]
    phv_data_176 <= io_pipe_phv_in_data_176; // @[parse_module.scala 51:9]
    phv_data_177 <= io_pipe_phv_in_data_177; // @[parse_module.scala 51:9]
    phv_data_178 <= io_pipe_phv_in_data_178; // @[parse_module.scala 51:9]
    phv_data_179 <= io_pipe_phv_in_data_179; // @[parse_module.scala 51:9]
    phv_data_180 <= io_pipe_phv_in_data_180; // @[parse_module.scala 51:9]
    phv_data_181 <= io_pipe_phv_in_data_181; // @[parse_module.scala 51:9]
    phv_data_182 <= io_pipe_phv_in_data_182; // @[parse_module.scala 51:9]
    phv_data_183 <= io_pipe_phv_in_data_183; // @[parse_module.scala 51:9]
    phv_data_184 <= io_pipe_phv_in_data_184; // @[parse_module.scala 51:9]
    phv_data_185 <= io_pipe_phv_in_data_185; // @[parse_module.scala 51:9]
    phv_data_186 <= io_pipe_phv_in_data_186; // @[parse_module.scala 51:9]
    phv_data_187 <= io_pipe_phv_in_data_187; // @[parse_module.scala 51:9]
    phv_data_188 <= io_pipe_phv_in_data_188; // @[parse_module.scala 51:9]
    phv_data_189 <= io_pipe_phv_in_data_189; // @[parse_module.scala 51:9]
    phv_data_190 <= io_pipe_phv_in_data_190; // @[parse_module.scala 51:9]
    phv_data_191 <= io_pipe_phv_in_data_191; // @[parse_module.scala 51:9]
    phv_data_192 <= io_pipe_phv_in_data_192; // @[parse_module.scala 51:9]
    phv_data_193 <= io_pipe_phv_in_data_193; // @[parse_module.scala 51:9]
    phv_data_194 <= io_pipe_phv_in_data_194; // @[parse_module.scala 51:9]
    phv_data_195 <= io_pipe_phv_in_data_195; // @[parse_module.scala 51:9]
    phv_data_196 <= io_pipe_phv_in_data_196; // @[parse_module.scala 51:9]
    phv_data_197 <= io_pipe_phv_in_data_197; // @[parse_module.scala 51:9]
    phv_data_198 <= io_pipe_phv_in_data_198; // @[parse_module.scala 51:9]
    phv_data_199 <= io_pipe_phv_in_data_199; // @[parse_module.scala 51:9]
    phv_data_200 <= io_pipe_phv_in_data_200; // @[parse_module.scala 51:9]
    phv_data_201 <= io_pipe_phv_in_data_201; // @[parse_module.scala 51:9]
    phv_data_202 <= io_pipe_phv_in_data_202; // @[parse_module.scala 51:9]
    phv_data_203 <= io_pipe_phv_in_data_203; // @[parse_module.scala 51:9]
    phv_data_204 <= io_pipe_phv_in_data_204; // @[parse_module.scala 51:9]
    phv_data_205 <= io_pipe_phv_in_data_205; // @[parse_module.scala 51:9]
    phv_data_206 <= io_pipe_phv_in_data_206; // @[parse_module.scala 51:9]
    phv_data_207 <= io_pipe_phv_in_data_207; // @[parse_module.scala 51:9]
    phv_data_208 <= io_pipe_phv_in_data_208; // @[parse_module.scala 51:9]
    phv_data_209 <= io_pipe_phv_in_data_209; // @[parse_module.scala 51:9]
    phv_data_210 <= io_pipe_phv_in_data_210; // @[parse_module.scala 51:9]
    phv_data_211 <= io_pipe_phv_in_data_211; // @[parse_module.scala 51:9]
    phv_data_212 <= io_pipe_phv_in_data_212; // @[parse_module.scala 51:9]
    phv_data_213 <= io_pipe_phv_in_data_213; // @[parse_module.scala 51:9]
    phv_data_214 <= io_pipe_phv_in_data_214; // @[parse_module.scala 51:9]
    phv_data_215 <= io_pipe_phv_in_data_215; // @[parse_module.scala 51:9]
    phv_data_216 <= io_pipe_phv_in_data_216; // @[parse_module.scala 51:9]
    phv_data_217 <= io_pipe_phv_in_data_217; // @[parse_module.scala 51:9]
    phv_data_218 <= io_pipe_phv_in_data_218; // @[parse_module.scala 51:9]
    phv_data_219 <= io_pipe_phv_in_data_219; // @[parse_module.scala 51:9]
    phv_data_220 <= io_pipe_phv_in_data_220; // @[parse_module.scala 51:9]
    phv_data_221 <= io_pipe_phv_in_data_221; // @[parse_module.scala 51:9]
    phv_data_222 <= io_pipe_phv_in_data_222; // @[parse_module.scala 51:9]
    phv_data_223 <= io_pipe_phv_in_data_223; // @[parse_module.scala 51:9]
    phv_data_224 <= io_pipe_phv_in_data_224; // @[parse_module.scala 51:9]
    phv_data_225 <= io_pipe_phv_in_data_225; // @[parse_module.scala 51:9]
    phv_data_226 <= io_pipe_phv_in_data_226; // @[parse_module.scala 51:9]
    phv_data_227 <= io_pipe_phv_in_data_227; // @[parse_module.scala 51:9]
    phv_data_228 <= io_pipe_phv_in_data_228; // @[parse_module.scala 51:9]
    phv_data_229 <= io_pipe_phv_in_data_229; // @[parse_module.scala 51:9]
    phv_data_230 <= io_pipe_phv_in_data_230; // @[parse_module.scala 51:9]
    phv_data_231 <= io_pipe_phv_in_data_231; // @[parse_module.scala 51:9]
    phv_data_232 <= io_pipe_phv_in_data_232; // @[parse_module.scala 51:9]
    phv_data_233 <= io_pipe_phv_in_data_233; // @[parse_module.scala 51:9]
    phv_data_234 <= io_pipe_phv_in_data_234; // @[parse_module.scala 51:9]
    phv_data_235 <= io_pipe_phv_in_data_235; // @[parse_module.scala 51:9]
    phv_data_236 <= io_pipe_phv_in_data_236; // @[parse_module.scala 51:9]
    phv_data_237 <= io_pipe_phv_in_data_237; // @[parse_module.scala 51:9]
    phv_data_238 <= io_pipe_phv_in_data_238; // @[parse_module.scala 51:9]
    phv_data_239 <= io_pipe_phv_in_data_239; // @[parse_module.scala 51:9]
    phv_data_240 <= io_pipe_phv_in_data_240; // @[parse_module.scala 51:9]
    phv_data_241 <= io_pipe_phv_in_data_241; // @[parse_module.scala 51:9]
    phv_data_242 <= io_pipe_phv_in_data_242; // @[parse_module.scala 51:9]
    phv_data_243 <= io_pipe_phv_in_data_243; // @[parse_module.scala 51:9]
    phv_data_244 <= io_pipe_phv_in_data_244; // @[parse_module.scala 51:9]
    phv_data_245 <= io_pipe_phv_in_data_245; // @[parse_module.scala 51:9]
    phv_data_246 <= io_pipe_phv_in_data_246; // @[parse_module.scala 51:9]
    phv_data_247 <= io_pipe_phv_in_data_247; // @[parse_module.scala 51:9]
    phv_data_248 <= io_pipe_phv_in_data_248; // @[parse_module.scala 51:9]
    phv_data_249 <= io_pipe_phv_in_data_249; // @[parse_module.scala 51:9]
    phv_data_250 <= io_pipe_phv_in_data_250; // @[parse_module.scala 51:9]
    phv_data_251 <= io_pipe_phv_in_data_251; // @[parse_module.scala 51:9]
    phv_data_252 <= io_pipe_phv_in_data_252; // @[parse_module.scala 51:9]
    phv_data_253 <= io_pipe_phv_in_data_253; // @[parse_module.scala 51:9]
    phv_data_254 <= io_pipe_phv_in_data_254; // @[parse_module.scala 51:9]
    phv_data_255 <= io_pipe_phv_in_data_255; // @[parse_module.scala 51:9]
    if (is_valid) begin // @[parse_module.scala 56:21]
      if (4'h0 == match_val_header_id[3:0]) begin // @[parse_module.scala 79:41]
        phv_header_0 <= _phv_header_T; // @[parse_module.scala 79:41]
      end else begin
        phv_header_0 <= io_pipe_phv_in_header_0; // @[parse_module.scala 51:9]
      end
    end else begin
      phv_header_0 <= io_pipe_phv_in_header_0; // @[parse_module.scala 51:9]
    end
    if (is_valid) begin // @[parse_module.scala 56:21]
      if (4'h1 == match_val_header_id[3:0]) begin // @[parse_module.scala 79:41]
        phv_header_1 <= _phv_header_T; // @[parse_module.scala 79:41]
      end else begin
        phv_header_1 <= io_pipe_phv_in_header_1; // @[parse_module.scala 51:9]
      end
    end else begin
      phv_header_1 <= io_pipe_phv_in_header_1; // @[parse_module.scala 51:9]
    end
    if (is_valid) begin // @[parse_module.scala 56:21]
      if (4'h2 == match_val_header_id[3:0]) begin // @[parse_module.scala 79:41]
        phv_header_2 <= _phv_header_T; // @[parse_module.scala 79:41]
      end else begin
        phv_header_2 <= io_pipe_phv_in_header_2; // @[parse_module.scala 51:9]
      end
    end else begin
      phv_header_2 <= io_pipe_phv_in_header_2; // @[parse_module.scala 51:9]
    end
    if (is_valid) begin // @[parse_module.scala 56:21]
      if (4'h3 == match_val_header_id[3:0]) begin // @[parse_module.scala 79:41]
        phv_header_3 <= _phv_header_T; // @[parse_module.scala 79:41]
      end else begin
        phv_header_3 <= io_pipe_phv_in_header_3; // @[parse_module.scala 51:9]
      end
    end else begin
      phv_header_3 <= io_pipe_phv_in_header_3; // @[parse_module.scala 51:9]
    end
    if (is_valid) begin // @[parse_module.scala 56:21]
      if (4'h4 == match_val_header_id[3:0]) begin // @[parse_module.scala 79:41]
        phv_header_4 <= _phv_header_T; // @[parse_module.scala 79:41]
      end else begin
        phv_header_4 <= io_pipe_phv_in_header_4; // @[parse_module.scala 51:9]
      end
    end else begin
      phv_header_4 <= io_pipe_phv_in_header_4; // @[parse_module.scala 51:9]
    end
    if (is_valid) begin // @[parse_module.scala 56:21]
      if (4'h5 == match_val_header_id[3:0]) begin // @[parse_module.scala 79:41]
        phv_header_5 <= _phv_header_T; // @[parse_module.scala 79:41]
      end else begin
        phv_header_5 <= io_pipe_phv_in_header_5; // @[parse_module.scala 51:9]
      end
    end else begin
      phv_header_5 <= io_pipe_phv_in_header_5; // @[parse_module.scala 51:9]
    end
    if (is_valid) begin // @[parse_module.scala 56:21]
      if (4'h6 == match_val_header_id[3:0]) begin // @[parse_module.scala 79:41]
        phv_header_6 <= _phv_header_T; // @[parse_module.scala 79:41]
      end else begin
        phv_header_6 <= io_pipe_phv_in_header_6; // @[parse_module.scala 51:9]
      end
    end else begin
      phv_header_6 <= io_pipe_phv_in_header_6; // @[parse_module.scala 51:9]
    end
    if (is_valid) begin // @[parse_module.scala 56:21]
      if (4'h7 == match_val_header_id[3:0]) begin // @[parse_module.scala 79:41]
        phv_header_7 <= _phv_header_T; // @[parse_module.scala 79:41]
      end else begin
        phv_header_7 <= io_pipe_phv_in_header_7; // @[parse_module.scala 51:9]
      end
    end else begin
      phv_header_7 <= io_pipe_phv_in_header_7; // @[parse_module.scala 51:9]
    end
    if (is_valid) begin // @[parse_module.scala 56:21]
      if (4'h8 == match_val_header_id[3:0]) begin // @[parse_module.scala 79:41]
        phv_header_8 <= _phv_header_T; // @[parse_module.scala 79:41]
      end else begin
        phv_header_8 <= io_pipe_phv_in_header_8; // @[parse_module.scala 51:9]
      end
    end else begin
      phv_header_8 <= io_pipe_phv_in_header_8; // @[parse_module.scala 51:9]
    end
    if (is_valid) begin // @[parse_module.scala 56:21]
      if (4'h9 == match_val_header_id[3:0]) begin // @[parse_module.scala 79:41]
        phv_header_9 <= _phv_header_T; // @[parse_module.scala 79:41]
      end else begin
        phv_header_9 <= io_pipe_phv_in_header_9; // @[parse_module.scala 51:9]
      end
    end else begin
      phv_header_9 <= io_pipe_phv_in_header_9; // @[parse_module.scala 51:9]
    end
    if (is_valid) begin // @[parse_module.scala 56:21]
      if (4'ha == match_val_header_id[3:0]) begin // @[parse_module.scala 79:41]
        phv_header_10 <= _phv_header_T; // @[parse_module.scala 79:41]
      end else begin
        phv_header_10 <= io_pipe_phv_in_header_10; // @[parse_module.scala 51:9]
      end
    end else begin
      phv_header_10 <= io_pipe_phv_in_header_10; // @[parse_module.scala 51:9]
    end
    if (is_valid) begin // @[parse_module.scala 56:21]
      if (4'hb == match_val_header_id[3:0]) begin // @[parse_module.scala 79:41]
        phv_header_11 <= _phv_header_T; // @[parse_module.scala 79:41]
      end else begin
        phv_header_11 <= io_pipe_phv_in_header_11; // @[parse_module.scala 51:9]
      end
    end else begin
      phv_header_11 <= io_pipe_phv_in_header_11; // @[parse_module.scala 51:9]
    end
    if (is_valid) begin // @[parse_module.scala 56:21]
      if (4'hc == match_val_header_id[3:0]) begin // @[parse_module.scala 79:41]
        phv_header_12 <= _phv_header_T; // @[parse_module.scala 79:41]
      end else begin
        phv_header_12 <= io_pipe_phv_in_header_12; // @[parse_module.scala 51:9]
      end
    end else begin
      phv_header_12 <= io_pipe_phv_in_header_12; // @[parse_module.scala 51:9]
    end
    if (is_valid) begin // @[parse_module.scala 56:21]
      if (4'hd == match_val_header_id[3:0]) begin // @[parse_module.scala 79:41]
        phv_header_13 <= _phv_header_T; // @[parse_module.scala 79:41]
      end else begin
        phv_header_13 <= io_pipe_phv_in_header_13; // @[parse_module.scala 51:9]
      end
    end else begin
      phv_header_13 <= io_pipe_phv_in_header_13; // @[parse_module.scala 51:9]
    end
    if (is_valid) begin // @[parse_module.scala 56:21]
      if (4'he == match_val_header_id[3:0]) begin // @[parse_module.scala 79:41]
        phv_header_14 <= _phv_header_T; // @[parse_module.scala 79:41]
      end else begin
        phv_header_14 <= io_pipe_phv_in_header_14; // @[parse_module.scala 51:9]
      end
    end else begin
      phv_header_14 <= io_pipe_phv_in_header_14; // @[parse_module.scala 51:9]
    end
    if (is_valid) begin // @[parse_module.scala 56:21]
      if (4'hf == match_val_header_id[3:0]) begin // @[parse_module.scala 79:41]
        phv_header_15 <= _phv_header_T; // @[parse_module.scala 79:41]
      end else begin
        phv_header_15 <= io_pipe_phv_in_header_15; // @[parse_module.scala 51:9]
      end
    end else begin
      phv_header_15 <= io_pipe_phv_in_header_15; // @[parse_module.scala 51:9]
    end
    if (is_valid) begin // @[parse_module.scala 56:21]
      phv_parse_current_state <= match_val_next_state; // @[parse_module.scala 67:34]
    end else begin
      phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[parse_module.scala 51:9]
    end
    if (is_valid) begin // @[parse_module.scala 56:21]
      phv_parse_current_offset <= _phv_parse_current_offset_T_1; // @[parse_module.scala 68:34]
    end else begin
      phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[parse_module.scala 51:9]
    end
    if (is_valid) begin // @[parse_module.scala 56:21]
      phv_parse_transition_field <= transition_field; // @[parse_module.scala 77:36]
    end else begin
      phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[parse_module.scala 51:9]
    end
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[parse_module.scala 51:9]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[parse_module.scala 51:9]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_data_160 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  phv_data_161 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  phv_data_162 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  phv_data_163 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  phv_data_164 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  phv_data_165 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  phv_data_166 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  phv_data_167 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  phv_data_168 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  phv_data_169 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  phv_data_170 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  phv_data_171 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  phv_data_172 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  phv_data_173 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  phv_data_174 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  phv_data_175 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  phv_data_176 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_data_177 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_data_178 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  phv_data_179 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  phv_data_180 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  phv_data_181 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  phv_data_182 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  phv_data_183 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  phv_data_184 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  phv_data_185 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  phv_data_186 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  phv_data_187 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  phv_data_188 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  phv_data_189 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  phv_data_190 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  phv_data_191 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  phv_data_192 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  phv_data_193 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  phv_data_194 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  phv_data_195 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  phv_data_196 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  phv_data_197 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  phv_data_198 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  phv_data_199 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  phv_data_200 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  phv_data_201 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  phv_data_202 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  phv_data_203 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  phv_data_204 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  phv_data_205 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  phv_data_206 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  phv_data_207 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  phv_data_208 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  phv_data_209 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  phv_data_210 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  phv_data_211 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  phv_data_212 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  phv_data_213 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  phv_data_214 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  phv_data_215 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  phv_data_216 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  phv_data_217 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  phv_data_218 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  phv_data_219 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  phv_data_220 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  phv_data_221 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  phv_data_222 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  phv_data_223 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  phv_data_224 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  phv_data_225 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  phv_data_226 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  phv_data_227 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  phv_data_228 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  phv_data_229 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  phv_data_230 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  phv_data_231 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  phv_data_232 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  phv_data_233 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  phv_data_234 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  phv_data_235 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  phv_data_236 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  phv_data_237 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  phv_data_238 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  phv_data_239 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  phv_data_240 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  phv_data_241 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  phv_data_242 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  phv_data_243 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  phv_data_244 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  phv_data_245 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  phv_data_246 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  phv_data_247 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  phv_data_248 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  phv_data_249 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  phv_data_250 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  phv_data_251 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  phv_data_252 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  phv_data_253 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  phv_data_254 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  phv_data_255 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  phv_header_0 = _RAND_256[15:0];
  _RAND_257 = {1{`RANDOM}};
  phv_header_1 = _RAND_257[15:0];
  _RAND_258 = {1{`RANDOM}};
  phv_header_2 = _RAND_258[15:0];
  _RAND_259 = {1{`RANDOM}};
  phv_header_3 = _RAND_259[15:0];
  _RAND_260 = {1{`RANDOM}};
  phv_header_4 = _RAND_260[15:0];
  _RAND_261 = {1{`RANDOM}};
  phv_header_5 = _RAND_261[15:0];
  _RAND_262 = {1{`RANDOM}};
  phv_header_6 = _RAND_262[15:0];
  _RAND_263 = {1{`RANDOM}};
  phv_header_7 = _RAND_263[15:0];
  _RAND_264 = {1{`RANDOM}};
  phv_header_8 = _RAND_264[15:0];
  _RAND_265 = {1{`RANDOM}};
  phv_header_9 = _RAND_265[15:0];
  _RAND_266 = {1{`RANDOM}};
  phv_header_10 = _RAND_266[15:0];
  _RAND_267 = {1{`RANDOM}};
  phv_header_11 = _RAND_267[15:0];
  _RAND_268 = {1{`RANDOM}};
  phv_header_12 = _RAND_268[15:0];
  _RAND_269 = {1{`RANDOM}};
  phv_header_13 = _RAND_269[15:0];
  _RAND_270 = {1{`RANDOM}};
  phv_header_14 = _RAND_270[15:0];
  _RAND_271 = {1{`RANDOM}};
  phv_header_15 = _RAND_271[15:0];
  _RAND_272 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_272[7:0];
  _RAND_273 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_273[7:0];
  _RAND_274 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_274[15:0];
  _RAND_275 = {1{`RANDOM}};
  phv_next_config_id = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_276[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
