module IPSASP(
  input         clock,
  input         reset,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [7:0]  io_pipe_phv_in_data_160,
  input  [7:0]  io_pipe_phv_in_data_161,
  input  [7:0]  io_pipe_phv_in_data_162,
  input  [7:0]  io_pipe_phv_in_data_163,
  input  [7:0]  io_pipe_phv_in_data_164,
  input  [7:0]  io_pipe_phv_in_data_165,
  input  [7:0]  io_pipe_phv_in_data_166,
  input  [7:0]  io_pipe_phv_in_data_167,
  input  [7:0]  io_pipe_phv_in_data_168,
  input  [7:0]  io_pipe_phv_in_data_169,
  input  [7:0]  io_pipe_phv_in_data_170,
  input  [7:0]  io_pipe_phv_in_data_171,
  input  [7:0]  io_pipe_phv_in_data_172,
  input  [7:0]  io_pipe_phv_in_data_173,
  input  [7:0]  io_pipe_phv_in_data_174,
  input  [7:0]  io_pipe_phv_in_data_175,
  input  [7:0]  io_pipe_phv_in_data_176,
  input  [7:0]  io_pipe_phv_in_data_177,
  input  [7:0]  io_pipe_phv_in_data_178,
  input  [7:0]  io_pipe_phv_in_data_179,
  input  [7:0]  io_pipe_phv_in_data_180,
  input  [7:0]  io_pipe_phv_in_data_181,
  input  [7:0]  io_pipe_phv_in_data_182,
  input  [7:0]  io_pipe_phv_in_data_183,
  input  [7:0]  io_pipe_phv_in_data_184,
  input  [7:0]  io_pipe_phv_in_data_185,
  input  [7:0]  io_pipe_phv_in_data_186,
  input  [7:0]  io_pipe_phv_in_data_187,
  input  [7:0]  io_pipe_phv_in_data_188,
  input  [7:0]  io_pipe_phv_in_data_189,
  input  [7:0]  io_pipe_phv_in_data_190,
  input  [7:0]  io_pipe_phv_in_data_191,
  input  [7:0]  io_pipe_phv_in_data_192,
  input  [7:0]  io_pipe_phv_in_data_193,
  input  [7:0]  io_pipe_phv_in_data_194,
  input  [7:0]  io_pipe_phv_in_data_195,
  input  [7:0]  io_pipe_phv_in_data_196,
  input  [7:0]  io_pipe_phv_in_data_197,
  input  [7:0]  io_pipe_phv_in_data_198,
  input  [7:0]  io_pipe_phv_in_data_199,
  input  [7:0]  io_pipe_phv_in_data_200,
  input  [7:0]  io_pipe_phv_in_data_201,
  input  [7:0]  io_pipe_phv_in_data_202,
  input  [7:0]  io_pipe_phv_in_data_203,
  input  [7:0]  io_pipe_phv_in_data_204,
  input  [7:0]  io_pipe_phv_in_data_205,
  input  [7:0]  io_pipe_phv_in_data_206,
  input  [7:0]  io_pipe_phv_in_data_207,
  input  [7:0]  io_pipe_phv_in_data_208,
  input  [7:0]  io_pipe_phv_in_data_209,
  input  [7:0]  io_pipe_phv_in_data_210,
  input  [7:0]  io_pipe_phv_in_data_211,
  input  [7:0]  io_pipe_phv_in_data_212,
  input  [7:0]  io_pipe_phv_in_data_213,
  input  [7:0]  io_pipe_phv_in_data_214,
  input  [7:0]  io_pipe_phv_in_data_215,
  input  [7:0]  io_pipe_phv_in_data_216,
  input  [7:0]  io_pipe_phv_in_data_217,
  input  [7:0]  io_pipe_phv_in_data_218,
  input  [7:0]  io_pipe_phv_in_data_219,
  input  [7:0]  io_pipe_phv_in_data_220,
  input  [7:0]  io_pipe_phv_in_data_221,
  input  [7:0]  io_pipe_phv_in_data_222,
  input  [7:0]  io_pipe_phv_in_data_223,
  input  [7:0]  io_pipe_phv_in_data_224,
  input  [7:0]  io_pipe_phv_in_data_225,
  input  [7:0]  io_pipe_phv_in_data_226,
  input  [7:0]  io_pipe_phv_in_data_227,
  input  [7:0]  io_pipe_phv_in_data_228,
  input  [7:0]  io_pipe_phv_in_data_229,
  input  [7:0]  io_pipe_phv_in_data_230,
  input  [7:0]  io_pipe_phv_in_data_231,
  input  [7:0]  io_pipe_phv_in_data_232,
  input  [7:0]  io_pipe_phv_in_data_233,
  input  [7:0]  io_pipe_phv_in_data_234,
  input  [7:0]  io_pipe_phv_in_data_235,
  input  [7:0]  io_pipe_phv_in_data_236,
  input  [7:0]  io_pipe_phv_in_data_237,
  input  [7:0]  io_pipe_phv_in_data_238,
  input  [7:0]  io_pipe_phv_in_data_239,
  input  [7:0]  io_pipe_phv_in_data_240,
  input  [7:0]  io_pipe_phv_in_data_241,
  input  [7:0]  io_pipe_phv_in_data_242,
  input  [7:0]  io_pipe_phv_in_data_243,
  input  [7:0]  io_pipe_phv_in_data_244,
  input  [7:0]  io_pipe_phv_in_data_245,
  input  [7:0]  io_pipe_phv_in_data_246,
  input  [7:0]  io_pipe_phv_in_data_247,
  input  [7:0]  io_pipe_phv_in_data_248,
  input  [7:0]  io_pipe_phv_in_data_249,
  input  [7:0]  io_pipe_phv_in_data_250,
  input  [7:0]  io_pipe_phv_in_data_251,
  input  [7:0]  io_pipe_phv_in_data_252,
  input  [7:0]  io_pipe_phv_in_data_253,
  input  [7:0]  io_pipe_phv_in_data_254,
  input  [7:0]  io_pipe_phv_in_data_255,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [3:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [7:0]  io_pipe_phv_out_data_160,
  output [7:0]  io_pipe_phv_out_data_161,
  output [7:0]  io_pipe_phv_out_data_162,
  output [7:0]  io_pipe_phv_out_data_163,
  output [7:0]  io_pipe_phv_out_data_164,
  output [7:0]  io_pipe_phv_out_data_165,
  output [7:0]  io_pipe_phv_out_data_166,
  output [7:0]  io_pipe_phv_out_data_167,
  output [7:0]  io_pipe_phv_out_data_168,
  output [7:0]  io_pipe_phv_out_data_169,
  output [7:0]  io_pipe_phv_out_data_170,
  output [7:0]  io_pipe_phv_out_data_171,
  output [7:0]  io_pipe_phv_out_data_172,
  output [7:0]  io_pipe_phv_out_data_173,
  output [7:0]  io_pipe_phv_out_data_174,
  output [7:0]  io_pipe_phv_out_data_175,
  output [7:0]  io_pipe_phv_out_data_176,
  output [7:0]  io_pipe_phv_out_data_177,
  output [7:0]  io_pipe_phv_out_data_178,
  output [7:0]  io_pipe_phv_out_data_179,
  output [7:0]  io_pipe_phv_out_data_180,
  output [7:0]  io_pipe_phv_out_data_181,
  output [7:0]  io_pipe_phv_out_data_182,
  output [7:0]  io_pipe_phv_out_data_183,
  output [7:0]  io_pipe_phv_out_data_184,
  output [7:0]  io_pipe_phv_out_data_185,
  output [7:0]  io_pipe_phv_out_data_186,
  output [7:0]  io_pipe_phv_out_data_187,
  output [7:0]  io_pipe_phv_out_data_188,
  output [7:0]  io_pipe_phv_out_data_189,
  output [7:0]  io_pipe_phv_out_data_190,
  output [7:0]  io_pipe_phv_out_data_191,
  output [7:0]  io_pipe_phv_out_data_192,
  output [7:0]  io_pipe_phv_out_data_193,
  output [7:0]  io_pipe_phv_out_data_194,
  output [7:0]  io_pipe_phv_out_data_195,
  output [7:0]  io_pipe_phv_out_data_196,
  output [7:0]  io_pipe_phv_out_data_197,
  output [7:0]  io_pipe_phv_out_data_198,
  output [7:0]  io_pipe_phv_out_data_199,
  output [7:0]  io_pipe_phv_out_data_200,
  output [7:0]  io_pipe_phv_out_data_201,
  output [7:0]  io_pipe_phv_out_data_202,
  output [7:0]  io_pipe_phv_out_data_203,
  output [7:0]  io_pipe_phv_out_data_204,
  output [7:0]  io_pipe_phv_out_data_205,
  output [7:0]  io_pipe_phv_out_data_206,
  output [7:0]  io_pipe_phv_out_data_207,
  output [7:0]  io_pipe_phv_out_data_208,
  output [7:0]  io_pipe_phv_out_data_209,
  output [7:0]  io_pipe_phv_out_data_210,
  output [7:0]  io_pipe_phv_out_data_211,
  output [7:0]  io_pipe_phv_out_data_212,
  output [7:0]  io_pipe_phv_out_data_213,
  output [7:0]  io_pipe_phv_out_data_214,
  output [7:0]  io_pipe_phv_out_data_215,
  output [7:0]  io_pipe_phv_out_data_216,
  output [7:0]  io_pipe_phv_out_data_217,
  output [7:0]  io_pipe_phv_out_data_218,
  output [7:0]  io_pipe_phv_out_data_219,
  output [7:0]  io_pipe_phv_out_data_220,
  output [7:0]  io_pipe_phv_out_data_221,
  output [7:0]  io_pipe_phv_out_data_222,
  output [7:0]  io_pipe_phv_out_data_223,
  output [7:0]  io_pipe_phv_out_data_224,
  output [7:0]  io_pipe_phv_out_data_225,
  output [7:0]  io_pipe_phv_out_data_226,
  output [7:0]  io_pipe_phv_out_data_227,
  output [7:0]  io_pipe_phv_out_data_228,
  output [7:0]  io_pipe_phv_out_data_229,
  output [7:0]  io_pipe_phv_out_data_230,
  output [7:0]  io_pipe_phv_out_data_231,
  output [7:0]  io_pipe_phv_out_data_232,
  output [7:0]  io_pipe_phv_out_data_233,
  output [7:0]  io_pipe_phv_out_data_234,
  output [7:0]  io_pipe_phv_out_data_235,
  output [7:0]  io_pipe_phv_out_data_236,
  output [7:0]  io_pipe_phv_out_data_237,
  output [7:0]  io_pipe_phv_out_data_238,
  output [7:0]  io_pipe_phv_out_data_239,
  output [7:0]  io_pipe_phv_out_data_240,
  output [7:0]  io_pipe_phv_out_data_241,
  output [7:0]  io_pipe_phv_out_data_242,
  output [7:0]  io_pipe_phv_out_data_243,
  output [7:0]  io_pipe_phv_out_data_244,
  output [7:0]  io_pipe_phv_out_data_245,
  output [7:0]  io_pipe_phv_out_data_246,
  output [7:0]  io_pipe_phv_out_data_247,
  output [7:0]  io_pipe_phv_out_data_248,
  output [7:0]  io_pipe_phv_out_data_249,
  output [7:0]  io_pipe_phv_out_data_250,
  output [7:0]  io_pipe_phv_out_data_251,
  output [7:0]  io_pipe_phv_out_data_252,
  output [7:0]  io_pipe_phv_out_data_253,
  output [7:0]  io_pipe_phv_out_data_254,
  output [7:0]  io_pipe_phv_out_data_255,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [3:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input         io_mod_par_mod_en,
  input         io_mod_par_mod_last_mau_id_mod,
  input  [1:0]  io_mod_par_mod_last_mau_id,
  input  [1:0]  io_mod_par_mod_cs,
  input         io_mod_par_mod_module_mod_state_id_mod,
  input  [7:0]  io_mod_par_mod_module_mod_state_id,
  input         io_mod_par_mod_module_mod_sram_w_cs,
  input         io_mod_par_mod_module_mod_sram_w_en,
  input  [7:0]  io_mod_par_mod_module_mod_sram_w_addr,
  input  [63:0] io_mod_par_mod_module_mod_sram_w_data,
  input         io_mod_mat_mod_en,
  input         io_mod_mat_mod_config_id,
  input  [7:0]  io_mod_mat_mod_key_mod_header_id,
  input  [7:0]  io_mod_mat_mod_key_mod_internal_offset,
  input  [7:0]  io_mod_mat_mod_key_mod_key_length,
  input  [3:0]  io_mod_mat_mod_key_mod_val_length,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_0,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_1,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_2,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_3,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_4,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_5,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_6,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_7,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_8,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_9,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_10,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_11,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_12,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_13,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_14,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_15,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_16,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_17,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_18,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_19,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_20,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_21,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_22,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_23,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_24,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_25,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_26,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_27,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_28,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_29,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_30,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_31,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_32,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_33,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_34,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_35,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_36,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_37,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_38,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_39,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_40,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_41,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_42,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_43,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_44,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_45,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_46,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_47,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_48,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_49,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_50,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_51,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_52,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_53,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_54,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_55,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_56,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_57,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_58,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_59,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_60,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_61,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_62,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_63,
  input  [6:0]  io_mod_mat_mod_table_mod_table_width,
  input  [6:0]  io_mod_mat_mod_table_mod_table_depth,
  input         io_mod_act_mod_en_0,
  input         io_mod_act_mod_en_1,
  input  [7:0]  io_mod_act_mod_addr,
  input  [63:0] io_mod_act_mod_data_0,
  input  [63:0] io_mod_act_mod_data_1,
  input  [5:0]  io_w_wcs,
  input         io_w_w_en,
  input  [7:0]  io_w_w_addr,
  input  [63:0] io_w_w_data
);
  wire  proc_clock; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_0; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_1; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_2; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_3; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_4; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_5; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_6; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_7; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_8; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_9; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_10; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_11; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_12; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_13; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_14; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_15; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_16; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_17; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_18; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_19; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_20; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_21; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_22; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_23; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_24; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_25; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_26; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_27; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_28; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_29; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_30; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_31; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_32; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_33; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_34; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_35; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_36; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_37; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_38; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_39; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_40; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_41; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_42; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_43; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_44; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_45; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_46; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_47; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_48; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_49; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_50; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_51; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_52; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_53; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_54; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_55; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_56; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_57; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_58; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_59; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_60; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_61; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_62; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_63; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_64; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_65; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_66; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_67; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_68; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_69; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_70; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_71; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_72; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_73; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_74; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_75; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_76; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_77; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_78; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_79; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_80; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_81; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_82; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_83; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_84; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_85; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_86; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_87; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_88; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_89; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_90; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_91; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_92; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_93; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_94; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_95; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_96; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_97; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_98; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_99; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_100; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_101; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_102; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_103; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_104; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_105; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_106; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_107; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_108; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_109; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_110; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_111; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_112; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_113; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_114; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_115; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_116; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_117; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_118; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_119; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_120; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_121; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_122; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_123; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_124; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_125; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_126; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_127; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_128; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_129; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_130; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_131; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_132; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_133; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_134; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_135; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_136; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_137; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_138; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_139; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_140; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_141; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_142; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_143; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_144; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_145; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_146; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_147; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_148; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_149; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_150; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_151; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_152; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_153; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_154; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_155; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_156; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_157; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_158; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_159; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_160; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_161; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_162; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_163; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_164; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_165; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_166; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_167; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_168; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_169; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_170; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_171; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_172; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_173; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_174; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_175; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_176; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_177; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_178; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_179; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_180; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_181; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_182; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_183; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_184; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_185; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_186; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_187; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_188; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_189; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_190; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_191; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_192; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_193; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_194; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_195; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_196; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_197; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_198; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_199; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_200; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_201; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_202; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_203; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_204; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_205; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_206; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_207; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_208; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_209; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_210; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_211; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_212; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_213; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_214; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_215; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_216; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_217; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_218; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_219; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_220; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_221; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_222; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_223; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_224; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_225; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_226; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_227; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_228; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_229; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_230; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_231; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_232; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_233; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_234; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_235; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_236; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_237; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_238; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_239; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_240; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_241; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_242; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_243; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_244; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_245; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_246; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_247; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_248; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_249; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_250; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_251; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_252; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_253; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_254; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_data_255; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_in_header_0; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_in_header_1; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_in_header_2; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_in_header_3; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_in_header_4; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_in_header_5; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_in_header_6; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_in_header_7; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_in_header_8; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_in_header_9; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_in_header_10; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_in_header_11; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_in_header_12; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_in_header_13; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_in_header_14; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_in_header_15; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_parse_current_state; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_in_parse_current_offset; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_in_parse_transition_field; // @[ipsa_single_processor.scala 14:22]
  wire [3:0] proc_io_pipe_phv_in_next_processor_id; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_pipe_phv_in_next_config_id; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_pipe_phv_in_is_valid_processor; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_0; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_1; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_2; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_3; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_4; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_5; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_6; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_7; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_8; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_9; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_10; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_11; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_12; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_13; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_14; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_15; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_16; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_17; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_18; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_19; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_20; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_21; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_22; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_23; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_24; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_25; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_26; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_27; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_28; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_29; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_30; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_31; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_32; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_33; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_34; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_35; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_36; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_37; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_38; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_39; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_40; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_41; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_42; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_43; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_44; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_45; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_46; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_47; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_48; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_49; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_50; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_51; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_52; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_53; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_54; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_55; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_56; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_57; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_58; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_59; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_60; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_61; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_62; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_63; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_64; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_65; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_66; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_67; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_68; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_69; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_70; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_71; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_72; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_73; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_74; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_75; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_76; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_77; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_78; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_79; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_80; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_81; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_82; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_83; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_84; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_85; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_86; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_87; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_88; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_89; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_90; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_91; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_92; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_93; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_94; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_95; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_96; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_97; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_98; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_99; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_100; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_101; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_102; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_103; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_104; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_105; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_106; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_107; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_108; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_109; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_110; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_111; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_112; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_113; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_114; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_115; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_116; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_117; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_118; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_119; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_120; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_121; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_122; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_123; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_124; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_125; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_126; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_127; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_128; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_129; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_130; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_131; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_132; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_133; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_134; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_135; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_136; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_137; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_138; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_139; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_140; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_141; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_142; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_143; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_144; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_145; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_146; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_147; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_148; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_149; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_150; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_151; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_152; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_153; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_154; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_155; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_156; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_157; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_158; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_159; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_160; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_161; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_162; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_163; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_164; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_165; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_166; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_167; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_168; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_169; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_170; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_171; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_172; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_173; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_174; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_175; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_176; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_177; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_178; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_179; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_180; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_181; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_182; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_183; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_184; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_185; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_186; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_187; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_188; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_189; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_190; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_191; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_192; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_193; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_194; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_195; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_196; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_197; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_198; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_199; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_200; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_201; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_202; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_203; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_204; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_205; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_206; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_207; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_208; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_209; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_210; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_211; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_212; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_213; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_214; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_215; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_216; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_217; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_218; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_219; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_220; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_221; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_222; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_223; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_224; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_225; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_226; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_227; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_228; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_229; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_230; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_231; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_232; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_233; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_234; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_235; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_236; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_237; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_238; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_239; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_240; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_241; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_242; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_243; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_244; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_245; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_246; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_247; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_248; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_249; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_250; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_251; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_252; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_253; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_254; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_data_255; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_out_header_0; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_out_header_1; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_out_header_2; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_out_header_3; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_out_header_4; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_out_header_5; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_out_header_6; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_out_header_7; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_out_header_8; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_out_header_9; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_out_header_10; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_out_header_11; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_out_header_12; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_out_header_13; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_out_header_14; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_out_header_15; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_parse_current_state; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_pipe_phv_out_parse_current_offset; // @[ipsa_single_processor.scala 14:22]
  wire [15:0] proc_io_pipe_phv_out_parse_transition_field; // @[ipsa_single_processor.scala 14:22]
  wire [3:0] proc_io_pipe_phv_out_next_processor_id; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_pipe_phv_out_next_config_id; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_pipe_phv_out_is_valid_processor; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mod_par_mod_en; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mod_par_mod_last_mau_id_mod; // @[ipsa_single_processor.scala 14:22]
  wire [1:0] proc_io_mod_par_mod_last_mau_id; // @[ipsa_single_processor.scala 14:22]
  wire [1:0] proc_io_mod_par_mod_cs; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mod_par_mod_module_mod_state_id_mod; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mod_par_mod_module_mod_state_id; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mod_par_mod_module_mod_sram_w_cs; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mod_par_mod_module_mod_sram_w_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mod_par_mod_module_mod_sram_w_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mod_par_mod_module_mod_sram_w_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mod_mat_mod_en; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mod_mat_mod_config_id; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mod_mat_mod_key_mod_header_id; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mod_mat_mod_key_mod_internal_offset; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mod_mat_mod_key_mod_key_length; // @[ipsa_single_processor.scala 14:22]
  wire [6:0] proc_io_mod_mat_mod_table_mod_table_width; // @[ipsa_single_processor.scala 14:22]
  wire [6:0] proc_io_mod_mat_mod_table_mod_table_depth; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mod_act_mod_en_0; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mod_act_mod_en_1; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mod_act_mod_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mod_act_mod_data_0; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mod_act_mod_data_1; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_0_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_0_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_0_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_1_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_1_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_1_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_2_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_2_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_2_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_3_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_3_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_3_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_4_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_4_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_4_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_5_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_5_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_5_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_6_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_6_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_6_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_7_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_7_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_7_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_8_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_8_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_8_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_9_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_9_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_9_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_10_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_10_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_10_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_11_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_11_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_11_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_12_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_12_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_12_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_13_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_13_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_13_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_14_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_14_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_14_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_15_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_15_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_15_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_16_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_16_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_16_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_17_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_17_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_17_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_18_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_18_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_18_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_19_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_19_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_19_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_20_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_20_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_20_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_21_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_21_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_21_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_22_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_22_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_22_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_23_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_23_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_23_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_24_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_24_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_24_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_25_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_25_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_25_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_26_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_26_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_26_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_27_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_27_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_27_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_28_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_28_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_28_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_29_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_29_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_29_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_30_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_30_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_30_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_31_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_31_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_31_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_32_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_32_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_32_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_33_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_33_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_33_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_34_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_34_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_34_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_35_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_35_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_35_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_36_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_36_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_36_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_37_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_37_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_37_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_38_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_38_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_38_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_39_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_39_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_39_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_40_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_40_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_40_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_41_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_41_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_41_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_42_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_42_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_42_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_43_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_43_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_43_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_44_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_44_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_44_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_45_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_45_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_45_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_46_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_46_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_46_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_47_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_47_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_47_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_48_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_48_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_48_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_49_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_49_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_49_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_50_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_50_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_50_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_51_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_51_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_51_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_52_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_52_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_52_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_53_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_53_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_53_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_54_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_54_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_54_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_55_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_55_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_55_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_56_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_56_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_56_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_57_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_57_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_57_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_58_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_58_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_58_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_59_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_59_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_59_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_60_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_60_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_60_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_61_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_61_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_61_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_62_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_62_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_62_data; // @[ipsa_single_processor.scala 14:22]
  wire  proc_io_mem_cluster_63_en; // @[ipsa_single_processor.scala 14:22]
  wire [7:0] proc_io_mem_cluster_63_addr; // @[ipsa_single_processor.scala 14:22]
  wire [63:0] proc_io_mem_cluster_63_data; // @[ipsa_single_processor.scala 14:22]
  wire  sram_cluster_clock; // @[ipsa_single_processor.scala 19:30]
  wire [5:0] sram_cluster_io_w_wcs; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_w_w_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_w_w_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_w_w_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_0_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_0_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_0_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_1_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_1_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_1_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_2_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_2_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_2_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_3_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_3_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_3_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_4_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_4_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_4_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_5_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_5_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_5_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_6_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_6_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_6_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_7_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_7_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_7_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_8_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_8_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_8_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_9_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_9_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_9_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_10_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_10_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_10_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_11_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_11_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_11_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_12_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_12_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_12_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_13_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_13_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_13_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_14_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_14_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_14_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_15_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_15_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_15_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_16_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_16_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_16_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_17_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_17_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_17_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_18_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_18_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_18_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_19_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_19_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_19_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_20_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_20_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_20_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_21_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_21_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_21_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_22_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_22_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_22_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_23_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_23_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_23_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_24_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_24_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_24_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_25_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_25_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_25_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_26_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_26_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_26_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_27_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_27_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_27_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_28_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_28_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_28_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_29_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_29_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_29_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_30_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_30_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_30_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_31_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_31_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_31_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_32_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_32_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_32_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_33_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_33_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_33_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_34_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_34_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_34_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_35_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_35_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_35_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_36_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_36_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_36_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_37_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_37_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_37_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_38_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_38_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_38_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_39_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_39_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_39_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_40_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_40_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_40_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_41_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_41_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_41_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_42_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_42_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_42_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_43_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_43_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_43_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_44_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_44_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_44_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_45_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_45_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_45_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_46_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_46_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_46_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_47_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_47_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_47_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_48_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_48_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_48_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_49_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_49_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_49_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_50_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_50_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_50_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_51_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_51_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_51_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_52_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_52_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_52_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_53_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_53_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_53_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_54_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_54_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_54_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_55_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_55_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_55_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_56_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_56_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_56_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_57_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_57_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_57_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_58_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_58_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_58_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_59_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_59_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_59_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_60_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_60_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_60_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_61_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_61_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_61_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_62_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_62_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_62_data; // @[ipsa_single_processor.scala 19:30]
  wire  sram_cluster_io_r_0_cluster_63_en; // @[ipsa_single_processor.scala 19:30]
  wire [7:0] sram_cluster_io_r_0_cluster_63_addr; // @[ipsa_single_processor.scala 19:30]
  wire [63:0] sram_cluster_io_r_0_cluster_63_data; // @[ipsa_single_processor.scala 19:30]
  Processor proc ( // @[ipsa_single_processor.scala 14:22]
    .clock(proc_clock),
    .io_pipe_phv_in_data_0(proc_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(proc_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(proc_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(proc_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(proc_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(proc_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(proc_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(proc_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(proc_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(proc_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(proc_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(proc_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(proc_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(proc_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(proc_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(proc_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(proc_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(proc_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(proc_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(proc_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(proc_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(proc_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(proc_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(proc_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(proc_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(proc_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(proc_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(proc_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(proc_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(proc_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(proc_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(proc_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(proc_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(proc_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(proc_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(proc_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(proc_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(proc_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(proc_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(proc_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(proc_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(proc_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(proc_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(proc_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(proc_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(proc_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(proc_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(proc_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(proc_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(proc_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(proc_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(proc_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(proc_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(proc_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(proc_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(proc_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(proc_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(proc_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(proc_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(proc_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(proc_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(proc_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(proc_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(proc_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(proc_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(proc_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(proc_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(proc_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(proc_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(proc_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(proc_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(proc_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(proc_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(proc_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(proc_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(proc_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(proc_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(proc_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(proc_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(proc_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(proc_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(proc_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(proc_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(proc_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(proc_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(proc_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(proc_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(proc_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(proc_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(proc_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(proc_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(proc_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(proc_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(proc_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(proc_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(proc_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(proc_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(proc_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(proc_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(proc_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(proc_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(proc_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(proc_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(proc_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(proc_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(proc_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(proc_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(proc_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(proc_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(proc_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(proc_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(proc_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(proc_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(proc_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(proc_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(proc_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(proc_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(proc_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(proc_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(proc_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(proc_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(proc_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(proc_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(proc_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(proc_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(proc_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(proc_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(proc_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(proc_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(proc_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(proc_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(proc_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(proc_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(proc_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(proc_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(proc_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(proc_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(proc_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(proc_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(proc_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(proc_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(proc_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(proc_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(proc_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(proc_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(proc_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(proc_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(proc_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(proc_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(proc_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(proc_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(proc_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(proc_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(proc_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(proc_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(proc_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(proc_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(proc_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(proc_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(proc_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(proc_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(proc_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(proc_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(proc_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(proc_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(proc_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(proc_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(proc_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(proc_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(proc_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(proc_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(proc_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(proc_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(proc_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(proc_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(proc_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(proc_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(proc_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(proc_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(proc_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(proc_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(proc_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(proc_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(proc_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(proc_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(proc_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(proc_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(proc_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(proc_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(proc_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(proc_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(proc_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(proc_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(proc_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(proc_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(proc_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(proc_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(proc_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(proc_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(proc_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(proc_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(proc_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(proc_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(proc_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(proc_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(proc_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(proc_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(proc_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(proc_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(proc_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(proc_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(proc_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(proc_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(proc_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(proc_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(proc_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(proc_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(proc_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(proc_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(proc_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(proc_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(proc_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(proc_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(proc_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(proc_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(proc_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(proc_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(proc_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(proc_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(proc_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(proc_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(proc_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(proc_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(proc_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(proc_io_pipe_phv_out_is_valid_processor),
    .io_mod_par_mod_en(proc_io_mod_par_mod_en),
    .io_mod_par_mod_last_mau_id_mod(proc_io_mod_par_mod_last_mau_id_mod),
    .io_mod_par_mod_last_mau_id(proc_io_mod_par_mod_last_mau_id),
    .io_mod_par_mod_cs(proc_io_mod_par_mod_cs),
    .io_mod_par_mod_module_mod_state_id_mod(proc_io_mod_par_mod_module_mod_state_id_mod),
    .io_mod_par_mod_module_mod_state_id(proc_io_mod_par_mod_module_mod_state_id),
    .io_mod_par_mod_module_mod_sram_w_cs(proc_io_mod_par_mod_module_mod_sram_w_cs),
    .io_mod_par_mod_module_mod_sram_w_en(proc_io_mod_par_mod_module_mod_sram_w_en),
    .io_mod_par_mod_module_mod_sram_w_addr(proc_io_mod_par_mod_module_mod_sram_w_addr),
    .io_mod_par_mod_module_mod_sram_w_data(proc_io_mod_par_mod_module_mod_sram_w_data),
    .io_mod_mat_mod_en(proc_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_header_id(proc_io_mod_mat_mod_key_mod_header_id),
    .io_mod_mat_mod_key_mod_internal_offset(proc_io_mod_mat_mod_key_mod_internal_offset),
    .io_mod_mat_mod_key_mod_key_length(proc_io_mod_mat_mod_key_mod_key_length),
    .io_mod_mat_mod_table_mod_table_width(proc_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_table_mod_table_depth(proc_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_act_mod_en_0(proc_io_mod_act_mod_en_0),
    .io_mod_act_mod_en_1(proc_io_mod_act_mod_en_1),
    .io_mod_act_mod_addr(proc_io_mod_act_mod_addr),
    .io_mod_act_mod_data_0(proc_io_mod_act_mod_data_0),
    .io_mod_act_mod_data_1(proc_io_mod_act_mod_data_1),
    .io_mem_cluster_0_en(proc_io_mem_cluster_0_en),
    .io_mem_cluster_0_addr(proc_io_mem_cluster_0_addr),
    .io_mem_cluster_0_data(proc_io_mem_cluster_0_data),
    .io_mem_cluster_1_en(proc_io_mem_cluster_1_en),
    .io_mem_cluster_1_addr(proc_io_mem_cluster_1_addr),
    .io_mem_cluster_1_data(proc_io_mem_cluster_1_data),
    .io_mem_cluster_2_en(proc_io_mem_cluster_2_en),
    .io_mem_cluster_2_addr(proc_io_mem_cluster_2_addr),
    .io_mem_cluster_2_data(proc_io_mem_cluster_2_data),
    .io_mem_cluster_3_en(proc_io_mem_cluster_3_en),
    .io_mem_cluster_3_addr(proc_io_mem_cluster_3_addr),
    .io_mem_cluster_3_data(proc_io_mem_cluster_3_data),
    .io_mem_cluster_4_en(proc_io_mem_cluster_4_en),
    .io_mem_cluster_4_addr(proc_io_mem_cluster_4_addr),
    .io_mem_cluster_4_data(proc_io_mem_cluster_4_data),
    .io_mem_cluster_5_en(proc_io_mem_cluster_5_en),
    .io_mem_cluster_5_addr(proc_io_mem_cluster_5_addr),
    .io_mem_cluster_5_data(proc_io_mem_cluster_5_data),
    .io_mem_cluster_6_en(proc_io_mem_cluster_6_en),
    .io_mem_cluster_6_addr(proc_io_mem_cluster_6_addr),
    .io_mem_cluster_6_data(proc_io_mem_cluster_6_data),
    .io_mem_cluster_7_en(proc_io_mem_cluster_7_en),
    .io_mem_cluster_7_addr(proc_io_mem_cluster_7_addr),
    .io_mem_cluster_7_data(proc_io_mem_cluster_7_data),
    .io_mem_cluster_8_en(proc_io_mem_cluster_8_en),
    .io_mem_cluster_8_addr(proc_io_mem_cluster_8_addr),
    .io_mem_cluster_8_data(proc_io_mem_cluster_8_data),
    .io_mem_cluster_9_en(proc_io_mem_cluster_9_en),
    .io_mem_cluster_9_addr(proc_io_mem_cluster_9_addr),
    .io_mem_cluster_9_data(proc_io_mem_cluster_9_data),
    .io_mem_cluster_10_en(proc_io_mem_cluster_10_en),
    .io_mem_cluster_10_addr(proc_io_mem_cluster_10_addr),
    .io_mem_cluster_10_data(proc_io_mem_cluster_10_data),
    .io_mem_cluster_11_en(proc_io_mem_cluster_11_en),
    .io_mem_cluster_11_addr(proc_io_mem_cluster_11_addr),
    .io_mem_cluster_11_data(proc_io_mem_cluster_11_data),
    .io_mem_cluster_12_en(proc_io_mem_cluster_12_en),
    .io_mem_cluster_12_addr(proc_io_mem_cluster_12_addr),
    .io_mem_cluster_12_data(proc_io_mem_cluster_12_data),
    .io_mem_cluster_13_en(proc_io_mem_cluster_13_en),
    .io_mem_cluster_13_addr(proc_io_mem_cluster_13_addr),
    .io_mem_cluster_13_data(proc_io_mem_cluster_13_data),
    .io_mem_cluster_14_en(proc_io_mem_cluster_14_en),
    .io_mem_cluster_14_addr(proc_io_mem_cluster_14_addr),
    .io_mem_cluster_14_data(proc_io_mem_cluster_14_data),
    .io_mem_cluster_15_en(proc_io_mem_cluster_15_en),
    .io_mem_cluster_15_addr(proc_io_mem_cluster_15_addr),
    .io_mem_cluster_15_data(proc_io_mem_cluster_15_data),
    .io_mem_cluster_16_en(proc_io_mem_cluster_16_en),
    .io_mem_cluster_16_addr(proc_io_mem_cluster_16_addr),
    .io_mem_cluster_16_data(proc_io_mem_cluster_16_data),
    .io_mem_cluster_17_en(proc_io_mem_cluster_17_en),
    .io_mem_cluster_17_addr(proc_io_mem_cluster_17_addr),
    .io_mem_cluster_17_data(proc_io_mem_cluster_17_data),
    .io_mem_cluster_18_en(proc_io_mem_cluster_18_en),
    .io_mem_cluster_18_addr(proc_io_mem_cluster_18_addr),
    .io_mem_cluster_18_data(proc_io_mem_cluster_18_data),
    .io_mem_cluster_19_en(proc_io_mem_cluster_19_en),
    .io_mem_cluster_19_addr(proc_io_mem_cluster_19_addr),
    .io_mem_cluster_19_data(proc_io_mem_cluster_19_data),
    .io_mem_cluster_20_en(proc_io_mem_cluster_20_en),
    .io_mem_cluster_20_addr(proc_io_mem_cluster_20_addr),
    .io_mem_cluster_20_data(proc_io_mem_cluster_20_data),
    .io_mem_cluster_21_en(proc_io_mem_cluster_21_en),
    .io_mem_cluster_21_addr(proc_io_mem_cluster_21_addr),
    .io_mem_cluster_21_data(proc_io_mem_cluster_21_data),
    .io_mem_cluster_22_en(proc_io_mem_cluster_22_en),
    .io_mem_cluster_22_addr(proc_io_mem_cluster_22_addr),
    .io_mem_cluster_22_data(proc_io_mem_cluster_22_data),
    .io_mem_cluster_23_en(proc_io_mem_cluster_23_en),
    .io_mem_cluster_23_addr(proc_io_mem_cluster_23_addr),
    .io_mem_cluster_23_data(proc_io_mem_cluster_23_data),
    .io_mem_cluster_24_en(proc_io_mem_cluster_24_en),
    .io_mem_cluster_24_addr(proc_io_mem_cluster_24_addr),
    .io_mem_cluster_24_data(proc_io_mem_cluster_24_data),
    .io_mem_cluster_25_en(proc_io_mem_cluster_25_en),
    .io_mem_cluster_25_addr(proc_io_mem_cluster_25_addr),
    .io_mem_cluster_25_data(proc_io_mem_cluster_25_data),
    .io_mem_cluster_26_en(proc_io_mem_cluster_26_en),
    .io_mem_cluster_26_addr(proc_io_mem_cluster_26_addr),
    .io_mem_cluster_26_data(proc_io_mem_cluster_26_data),
    .io_mem_cluster_27_en(proc_io_mem_cluster_27_en),
    .io_mem_cluster_27_addr(proc_io_mem_cluster_27_addr),
    .io_mem_cluster_27_data(proc_io_mem_cluster_27_data),
    .io_mem_cluster_28_en(proc_io_mem_cluster_28_en),
    .io_mem_cluster_28_addr(proc_io_mem_cluster_28_addr),
    .io_mem_cluster_28_data(proc_io_mem_cluster_28_data),
    .io_mem_cluster_29_en(proc_io_mem_cluster_29_en),
    .io_mem_cluster_29_addr(proc_io_mem_cluster_29_addr),
    .io_mem_cluster_29_data(proc_io_mem_cluster_29_data),
    .io_mem_cluster_30_en(proc_io_mem_cluster_30_en),
    .io_mem_cluster_30_addr(proc_io_mem_cluster_30_addr),
    .io_mem_cluster_30_data(proc_io_mem_cluster_30_data),
    .io_mem_cluster_31_en(proc_io_mem_cluster_31_en),
    .io_mem_cluster_31_addr(proc_io_mem_cluster_31_addr),
    .io_mem_cluster_31_data(proc_io_mem_cluster_31_data),
    .io_mem_cluster_32_en(proc_io_mem_cluster_32_en),
    .io_mem_cluster_32_addr(proc_io_mem_cluster_32_addr),
    .io_mem_cluster_32_data(proc_io_mem_cluster_32_data),
    .io_mem_cluster_33_en(proc_io_mem_cluster_33_en),
    .io_mem_cluster_33_addr(proc_io_mem_cluster_33_addr),
    .io_mem_cluster_33_data(proc_io_mem_cluster_33_data),
    .io_mem_cluster_34_en(proc_io_mem_cluster_34_en),
    .io_mem_cluster_34_addr(proc_io_mem_cluster_34_addr),
    .io_mem_cluster_34_data(proc_io_mem_cluster_34_data),
    .io_mem_cluster_35_en(proc_io_mem_cluster_35_en),
    .io_mem_cluster_35_addr(proc_io_mem_cluster_35_addr),
    .io_mem_cluster_35_data(proc_io_mem_cluster_35_data),
    .io_mem_cluster_36_en(proc_io_mem_cluster_36_en),
    .io_mem_cluster_36_addr(proc_io_mem_cluster_36_addr),
    .io_mem_cluster_36_data(proc_io_mem_cluster_36_data),
    .io_mem_cluster_37_en(proc_io_mem_cluster_37_en),
    .io_mem_cluster_37_addr(proc_io_mem_cluster_37_addr),
    .io_mem_cluster_37_data(proc_io_mem_cluster_37_data),
    .io_mem_cluster_38_en(proc_io_mem_cluster_38_en),
    .io_mem_cluster_38_addr(proc_io_mem_cluster_38_addr),
    .io_mem_cluster_38_data(proc_io_mem_cluster_38_data),
    .io_mem_cluster_39_en(proc_io_mem_cluster_39_en),
    .io_mem_cluster_39_addr(proc_io_mem_cluster_39_addr),
    .io_mem_cluster_39_data(proc_io_mem_cluster_39_data),
    .io_mem_cluster_40_en(proc_io_mem_cluster_40_en),
    .io_mem_cluster_40_addr(proc_io_mem_cluster_40_addr),
    .io_mem_cluster_40_data(proc_io_mem_cluster_40_data),
    .io_mem_cluster_41_en(proc_io_mem_cluster_41_en),
    .io_mem_cluster_41_addr(proc_io_mem_cluster_41_addr),
    .io_mem_cluster_41_data(proc_io_mem_cluster_41_data),
    .io_mem_cluster_42_en(proc_io_mem_cluster_42_en),
    .io_mem_cluster_42_addr(proc_io_mem_cluster_42_addr),
    .io_mem_cluster_42_data(proc_io_mem_cluster_42_data),
    .io_mem_cluster_43_en(proc_io_mem_cluster_43_en),
    .io_mem_cluster_43_addr(proc_io_mem_cluster_43_addr),
    .io_mem_cluster_43_data(proc_io_mem_cluster_43_data),
    .io_mem_cluster_44_en(proc_io_mem_cluster_44_en),
    .io_mem_cluster_44_addr(proc_io_mem_cluster_44_addr),
    .io_mem_cluster_44_data(proc_io_mem_cluster_44_data),
    .io_mem_cluster_45_en(proc_io_mem_cluster_45_en),
    .io_mem_cluster_45_addr(proc_io_mem_cluster_45_addr),
    .io_mem_cluster_45_data(proc_io_mem_cluster_45_data),
    .io_mem_cluster_46_en(proc_io_mem_cluster_46_en),
    .io_mem_cluster_46_addr(proc_io_mem_cluster_46_addr),
    .io_mem_cluster_46_data(proc_io_mem_cluster_46_data),
    .io_mem_cluster_47_en(proc_io_mem_cluster_47_en),
    .io_mem_cluster_47_addr(proc_io_mem_cluster_47_addr),
    .io_mem_cluster_47_data(proc_io_mem_cluster_47_data),
    .io_mem_cluster_48_en(proc_io_mem_cluster_48_en),
    .io_mem_cluster_48_addr(proc_io_mem_cluster_48_addr),
    .io_mem_cluster_48_data(proc_io_mem_cluster_48_data),
    .io_mem_cluster_49_en(proc_io_mem_cluster_49_en),
    .io_mem_cluster_49_addr(proc_io_mem_cluster_49_addr),
    .io_mem_cluster_49_data(proc_io_mem_cluster_49_data),
    .io_mem_cluster_50_en(proc_io_mem_cluster_50_en),
    .io_mem_cluster_50_addr(proc_io_mem_cluster_50_addr),
    .io_mem_cluster_50_data(proc_io_mem_cluster_50_data),
    .io_mem_cluster_51_en(proc_io_mem_cluster_51_en),
    .io_mem_cluster_51_addr(proc_io_mem_cluster_51_addr),
    .io_mem_cluster_51_data(proc_io_mem_cluster_51_data),
    .io_mem_cluster_52_en(proc_io_mem_cluster_52_en),
    .io_mem_cluster_52_addr(proc_io_mem_cluster_52_addr),
    .io_mem_cluster_52_data(proc_io_mem_cluster_52_data),
    .io_mem_cluster_53_en(proc_io_mem_cluster_53_en),
    .io_mem_cluster_53_addr(proc_io_mem_cluster_53_addr),
    .io_mem_cluster_53_data(proc_io_mem_cluster_53_data),
    .io_mem_cluster_54_en(proc_io_mem_cluster_54_en),
    .io_mem_cluster_54_addr(proc_io_mem_cluster_54_addr),
    .io_mem_cluster_54_data(proc_io_mem_cluster_54_data),
    .io_mem_cluster_55_en(proc_io_mem_cluster_55_en),
    .io_mem_cluster_55_addr(proc_io_mem_cluster_55_addr),
    .io_mem_cluster_55_data(proc_io_mem_cluster_55_data),
    .io_mem_cluster_56_en(proc_io_mem_cluster_56_en),
    .io_mem_cluster_56_addr(proc_io_mem_cluster_56_addr),
    .io_mem_cluster_56_data(proc_io_mem_cluster_56_data),
    .io_mem_cluster_57_en(proc_io_mem_cluster_57_en),
    .io_mem_cluster_57_addr(proc_io_mem_cluster_57_addr),
    .io_mem_cluster_57_data(proc_io_mem_cluster_57_data),
    .io_mem_cluster_58_en(proc_io_mem_cluster_58_en),
    .io_mem_cluster_58_addr(proc_io_mem_cluster_58_addr),
    .io_mem_cluster_58_data(proc_io_mem_cluster_58_data),
    .io_mem_cluster_59_en(proc_io_mem_cluster_59_en),
    .io_mem_cluster_59_addr(proc_io_mem_cluster_59_addr),
    .io_mem_cluster_59_data(proc_io_mem_cluster_59_data),
    .io_mem_cluster_60_en(proc_io_mem_cluster_60_en),
    .io_mem_cluster_60_addr(proc_io_mem_cluster_60_addr),
    .io_mem_cluster_60_data(proc_io_mem_cluster_60_data),
    .io_mem_cluster_61_en(proc_io_mem_cluster_61_en),
    .io_mem_cluster_61_addr(proc_io_mem_cluster_61_addr),
    .io_mem_cluster_61_data(proc_io_mem_cluster_61_data),
    .io_mem_cluster_62_en(proc_io_mem_cluster_62_en),
    .io_mem_cluster_62_addr(proc_io_mem_cluster_62_addr),
    .io_mem_cluster_62_data(proc_io_mem_cluster_62_data),
    .io_mem_cluster_63_en(proc_io_mem_cluster_63_en),
    .io_mem_cluster_63_addr(proc_io_mem_cluster_63_addr),
    .io_mem_cluster_63_data(proc_io_mem_cluster_63_data)
  );
  SRAMCluster sram_cluster ( // @[ipsa_single_processor.scala 19:30]
    .clock(sram_cluster_clock),
    .io_w_wcs(sram_cluster_io_w_wcs),
    .io_w_w_en(sram_cluster_io_w_w_en),
    .io_w_w_addr(sram_cluster_io_w_w_addr),
    .io_w_w_data(sram_cluster_io_w_w_data),
    .io_r_0_cluster_0_en(sram_cluster_io_r_0_cluster_0_en),
    .io_r_0_cluster_0_addr(sram_cluster_io_r_0_cluster_0_addr),
    .io_r_0_cluster_0_data(sram_cluster_io_r_0_cluster_0_data),
    .io_r_0_cluster_1_en(sram_cluster_io_r_0_cluster_1_en),
    .io_r_0_cluster_1_addr(sram_cluster_io_r_0_cluster_1_addr),
    .io_r_0_cluster_1_data(sram_cluster_io_r_0_cluster_1_data),
    .io_r_0_cluster_2_en(sram_cluster_io_r_0_cluster_2_en),
    .io_r_0_cluster_2_addr(sram_cluster_io_r_0_cluster_2_addr),
    .io_r_0_cluster_2_data(sram_cluster_io_r_0_cluster_2_data),
    .io_r_0_cluster_3_en(sram_cluster_io_r_0_cluster_3_en),
    .io_r_0_cluster_3_addr(sram_cluster_io_r_0_cluster_3_addr),
    .io_r_0_cluster_3_data(sram_cluster_io_r_0_cluster_3_data),
    .io_r_0_cluster_4_en(sram_cluster_io_r_0_cluster_4_en),
    .io_r_0_cluster_4_addr(sram_cluster_io_r_0_cluster_4_addr),
    .io_r_0_cluster_4_data(sram_cluster_io_r_0_cluster_4_data),
    .io_r_0_cluster_5_en(sram_cluster_io_r_0_cluster_5_en),
    .io_r_0_cluster_5_addr(sram_cluster_io_r_0_cluster_5_addr),
    .io_r_0_cluster_5_data(sram_cluster_io_r_0_cluster_5_data),
    .io_r_0_cluster_6_en(sram_cluster_io_r_0_cluster_6_en),
    .io_r_0_cluster_6_addr(sram_cluster_io_r_0_cluster_6_addr),
    .io_r_0_cluster_6_data(sram_cluster_io_r_0_cluster_6_data),
    .io_r_0_cluster_7_en(sram_cluster_io_r_0_cluster_7_en),
    .io_r_0_cluster_7_addr(sram_cluster_io_r_0_cluster_7_addr),
    .io_r_0_cluster_7_data(sram_cluster_io_r_0_cluster_7_data),
    .io_r_0_cluster_8_en(sram_cluster_io_r_0_cluster_8_en),
    .io_r_0_cluster_8_addr(sram_cluster_io_r_0_cluster_8_addr),
    .io_r_0_cluster_8_data(sram_cluster_io_r_0_cluster_8_data),
    .io_r_0_cluster_9_en(sram_cluster_io_r_0_cluster_9_en),
    .io_r_0_cluster_9_addr(sram_cluster_io_r_0_cluster_9_addr),
    .io_r_0_cluster_9_data(sram_cluster_io_r_0_cluster_9_data),
    .io_r_0_cluster_10_en(sram_cluster_io_r_0_cluster_10_en),
    .io_r_0_cluster_10_addr(sram_cluster_io_r_0_cluster_10_addr),
    .io_r_0_cluster_10_data(sram_cluster_io_r_0_cluster_10_data),
    .io_r_0_cluster_11_en(sram_cluster_io_r_0_cluster_11_en),
    .io_r_0_cluster_11_addr(sram_cluster_io_r_0_cluster_11_addr),
    .io_r_0_cluster_11_data(sram_cluster_io_r_0_cluster_11_data),
    .io_r_0_cluster_12_en(sram_cluster_io_r_0_cluster_12_en),
    .io_r_0_cluster_12_addr(sram_cluster_io_r_0_cluster_12_addr),
    .io_r_0_cluster_12_data(sram_cluster_io_r_0_cluster_12_data),
    .io_r_0_cluster_13_en(sram_cluster_io_r_0_cluster_13_en),
    .io_r_0_cluster_13_addr(sram_cluster_io_r_0_cluster_13_addr),
    .io_r_0_cluster_13_data(sram_cluster_io_r_0_cluster_13_data),
    .io_r_0_cluster_14_en(sram_cluster_io_r_0_cluster_14_en),
    .io_r_0_cluster_14_addr(sram_cluster_io_r_0_cluster_14_addr),
    .io_r_0_cluster_14_data(sram_cluster_io_r_0_cluster_14_data),
    .io_r_0_cluster_15_en(sram_cluster_io_r_0_cluster_15_en),
    .io_r_0_cluster_15_addr(sram_cluster_io_r_0_cluster_15_addr),
    .io_r_0_cluster_15_data(sram_cluster_io_r_0_cluster_15_data),
    .io_r_0_cluster_16_en(sram_cluster_io_r_0_cluster_16_en),
    .io_r_0_cluster_16_addr(sram_cluster_io_r_0_cluster_16_addr),
    .io_r_0_cluster_16_data(sram_cluster_io_r_0_cluster_16_data),
    .io_r_0_cluster_17_en(sram_cluster_io_r_0_cluster_17_en),
    .io_r_0_cluster_17_addr(sram_cluster_io_r_0_cluster_17_addr),
    .io_r_0_cluster_17_data(sram_cluster_io_r_0_cluster_17_data),
    .io_r_0_cluster_18_en(sram_cluster_io_r_0_cluster_18_en),
    .io_r_0_cluster_18_addr(sram_cluster_io_r_0_cluster_18_addr),
    .io_r_0_cluster_18_data(sram_cluster_io_r_0_cluster_18_data),
    .io_r_0_cluster_19_en(sram_cluster_io_r_0_cluster_19_en),
    .io_r_0_cluster_19_addr(sram_cluster_io_r_0_cluster_19_addr),
    .io_r_0_cluster_19_data(sram_cluster_io_r_0_cluster_19_data),
    .io_r_0_cluster_20_en(sram_cluster_io_r_0_cluster_20_en),
    .io_r_0_cluster_20_addr(sram_cluster_io_r_0_cluster_20_addr),
    .io_r_0_cluster_20_data(sram_cluster_io_r_0_cluster_20_data),
    .io_r_0_cluster_21_en(sram_cluster_io_r_0_cluster_21_en),
    .io_r_0_cluster_21_addr(sram_cluster_io_r_0_cluster_21_addr),
    .io_r_0_cluster_21_data(sram_cluster_io_r_0_cluster_21_data),
    .io_r_0_cluster_22_en(sram_cluster_io_r_0_cluster_22_en),
    .io_r_0_cluster_22_addr(sram_cluster_io_r_0_cluster_22_addr),
    .io_r_0_cluster_22_data(sram_cluster_io_r_0_cluster_22_data),
    .io_r_0_cluster_23_en(sram_cluster_io_r_0_cluster_23_en),
    .io_r_0_cluster_23_addr(sram_cluster_io_r_0_cluster_23_addr),
    .io_r_0_cluster_23_data(sram_cluster_io_r_0_cluster_23_data),
    .io_r_0_cluster_24_en(sram_cluster_io_r_0_cluster_24_en),
    .io_r_0_cluster_24_addr(sram_cluster_io_r_0_cluster_24_addr),
    .io_r_0_cluster_24_data(sram_cluster_io_r_0_cluster_24_data),
    .io_r_0_cluster_25_en(sram_cluster_io_r_0_cluster_25_en),
    .io_r_0_cluster_25_addr(sram_cluster_io_r_0_cluster_25_addr),
    .io_r_0_cluster_25_data(sram_cluster_io_r_0_cluster_25_data),
    .io_r_0_cluster_26_en(sram_cluster_io_r_0_cluster_26_en),
    .io_r_0_cluster_26_addr(sram_cluster_io_r_0_cluster_26_addr),
    .io_r_0_cluster_26_data(sram_cluster_io_r_0_cluster_26_data),
    .io_r_0_cluster_27_en(sram_cluster_io_r_0_cluster_27_en),
    .io_r_0_cluster_27_addr(sram_cluster_io_r_0_cluster_27_addr),
    .io_r_0_cluster_27_data(sram_cluster_io_r_0_cluster_27_data),
    .io_r_0_cluster_28_en(sram_cluster_io_r_0_cluster_28_en),
    .io_r_0_cluster_28_addr(sram_cluster_io_r_0_cluster_28_addr),
    .io_r_0_cluster_28_data(sram_cluster_io_r_0_cluster_28_data),
    .io_r_0_cluster_29_en(sram_cluster_io_r_0_cluster_29_en),
    .io_r_0_cluster_29_addr(sram_cluster_io_r_0_cluster_29_addr),
    .io_r_0_cluster_29_data(sram_cluster_io_r_0_cluster_29_data),
    .io_r_0_cluster_30_en(sram_cluster_io_r_0_cluster_30_en),
    .io_r_0_cluster_30_addr(sram_cluster_io_r_0_cluster_30_addr),
    .io_r_0_cluster_30_data(sram_cluster_io_r_0_cluster_30_data),
    .io_r_0_cluster_31_en(sram_cluster_io_r_0_cluster_31_en),
    .io_r_0_cluster_31_addr(sram_cluster_io_r_0_cluster_31_addr),
    .io_r_0_cluster_31_data(sram_cluster_io_r_0_cluster_31_data),
    .io_r_0_cluster_32_en(sram_cluster_io_r_0_cluster_32_en),
    .io_r_0_cluster_32_addr(sram_cluster_io_r_0_cluster_32_addr),
    .io_r_0_cluster_32_data(sram_cluster_io_r_0_cluster_32_data),
    .io_r_0_cluster_33_en(sram_cluster_io_r_0_cluster_33_en),
    .io_r_0_cluster_33_addr(sram_cluster_io_r_0_cluster_33_addr),
    .io_r_0_cluster_33_data(sram_cluster_io_r_0_cluster_33_data),
    .io_r_0_cluster_34_en(sram_cluster_io_r_0_cluster_34_en),
    .io_r_0_cluster_34_addr(sram_cluster_io_r_0_cluster_34_addr),
    .io_r_0_cluster_34_data(sram_cluster_io_r_0_cluster_34_data),
    .io_r_0_cluster_35_en(sram_cluster_io_r_0_cluster_35_en),
    .io_r_0_cluster_35_addr(sram_cluster_io_r_0_cluster_35_addr),
    .io_r_0_cluster_35_data(sram_cluster_io_r_0_cluster_35_data),
    .io_r_0_cluster_36_en(sram_cluster_io_r_0_cluster_36_en),
    .io_r_0_cluster_36_addr(sram_cluster_io_r_0_cluster_36_addr),
    .io_r_0_cluster_36_data(sram_cluster_io_r_0_cluster_36_data),
    .io_r_0_cluster_37_en(sram_cluster_io_r_0_cluster_37_en),
    .io_r_0_cluster_37_addr(sram_cluster_io_r_0_cluster_37_addr),
    .io_r_0_cluster_37_data(sram_cluster_io_r_0_cluster_37_data),
    .io_r_0_cluster_38_en(sram_cluster_io_r_0_cluster_38_en),
    .io_r_0_cluster_38_addr(sram_cluster_io_r_0_cluster_38_addr),
    .io_r_0_cluster_38_data(sram_cluster_io_r_0_cluster_38_data),
    .io_r_0_cluster_39_en(sram_cluster_io_r_0_cluster_39_en),
    .io_r_0_cluster_39_addr(sram_cluster_io_r_0_cluster_39_addr),
    .io_r_0_cluster_39_data(sram_cluster_io_r_0_cluster_39_data),
    .io_r_0_cluster_40_en(sram_cluster_io_r_0_cluster_40_en),
    .io_r_0_cluster_40_addr(sram_cluster_io_r_0_cluster_40_addr),
    .io_r_0_cluster_40_data(sram_cluster_io_r_0_cluster_40_data),
    .io_r_0_cluster_41_en(sram_cluster_io_r_0_cluster_41_en),
    .io_r_0_cluster_41_addr(sram_cluster_io_r_0_cluster_41_addr),
    .io_r_0_cluster_41_data(sram_cluster_io_r_0_cluster_41_data),
    .io_r_0_cluster_42_en(sram_cluster_io_r_0_cluster_42_en),
    .io_r_0_cluster_42_addr(sram_cluster_io_r_0_cluster_42_addr),
    .io_r_0_cluster_42_data(sram_cluster_io_r_0_cluster_42_data),
    .io_r_0_cluster_43_en(sram_cluster_io_r_0_cluster_43_en),
    .io_r_0_cluster_43_addr(sram_cluster_io_r_0_cluster_43_addr),
    .io_r_0_cluster_43_data(sram_cluster_io_r_0_cluster_43_data),
    .io_r_0_cluster_44_en(sram_cluster_io_r_0_cluster_44_en),
    .io_r_0_cluster_44_addr(sram_cluster_io_r_0_cluster_44_addr),
    .io_r_0_cluster_44_data(sram_cluster_io_r_0_cluster_44_data),
    .io_r_0_cluster_45_en(sram_cluster_io_r_0_cluster_45_en),
    .io_r_0_cluster_45_addr(sram_cluster_io_r_0_cluster_45_addr),
    .io_r_0_cluster_45_data(sram_cluster_io_r_0_cluster_45_data),
    .io_r_0_cluster_46_en(sram_cluster_io_r_0_cluster_46_en),
    .io_r_0_cluster_46_addr(sram_cluster_io_r_0_cluster_46_addr),
    .io_r_0_cluster_46_data(sram_cluster_io_r_0_cluster_46_data),
    .io_r_0_cluster_47_en(sram_cluster_io_r_0_cluster_47_en),
    .io_r_0_cluster_47_addr(sram_cluster_io_r_0_cluster_47_addr),
    .io_r_0_cluster_47_data(sram_cluster_io_r_0_cluster_47_data),
    .io_r_0_cluster_48_en(sram_cluster_io_r_0_cluster_48_en),
    .io_r_0_cluster_48_addr(sram_cluster_io_r_0_cluster_48_addr),
    .io_r_0_cluster_48_data(sram_cluster_io_r_0_cluster_48_data),
    .io_r_0_cluster_49_en(sram_cluster_io_r_0_cluster_49_en),
    .io_r_0_cluster_49_addr(sram_cluster_io_r_0_cluster_49_addr),
    .io_r_0_cluster_49_data(sram_cluster_io_r_0_cluster_49_data),
    .io_r_0_cluster_50_en(sram_cluster_io_r_0_cluster_50_en),
    .io_r_0_cluster_50_addr(sram_cluster_io_r_0_cluster_50_addr),
    .io_r_0_cluster_50_data(sram_cluster_io_r_0_cluster_50_data),
    .io_r_0_cluster_51_en(sram_cluster_io_r_0_cluster_51_en),
    .io_r_0_cluster_51_addr(sram_cluster_io_r_0_cluster_51_addr),
    .io_r_0_cluster_51_data(sram_cluster_io_r_0_cluster_51_data),
    .io_r_0_cluster_52_en(sram_cluster_io_r_0_cluster_52_en),
    .io_r_0_cluster_52_addr(sram_cluster_io_r_0_cluster_52_addr),
    .io_r_0_cluster_52_data(sram_cluster_io_r_0_cluster_52_data),
    .io_r_0_cluster_53_en(sram_cluster_io_r_0_cluster_53_en),
    .io_r_0_cluster_53_addr(sram_cluster_io_r_0_cluster_53_addr),
    .io_r_0_cluster_53_data(sram_cluster_io_r_0_cluster_53_data),
    .io_r_0_cluster_54_en(sram_cluster_io_r_0_cluster_54_en),
    .io_r_0_cluster_54_addr(sram_cluster_io_r_0_cluster_54_addr),
    .io_r_0_cluster_54_data(sram_cluster_io_r_0_cluster_54_data),
    .io_r_0_cluster_55_en(sram_cluster_io_r_0_cluster_55_en),
    .io_r_0_cluster_55_addr(sram_cluster_io_r_0_cluster_55_addr),
    .io_r_0_cluster_55_data(sram_cluster_io_r_0_cluster_55_data),
    .io_r_0_cluster_56_en(sram_cluster_io_r_0_cluster_56_en),
    .io_r_0_cluster_56_addr(sram_cluster_io_r_0_cluster_56_addr),
    .io_r_0_cluster_56_data(sram_cluster_io_r_0_cluster_56_data),
    .io_r_0_cluster_57_en(sram_cluster_io_r_0_cluster_57_en),
    .io_r_0_cluster_57_addr(sram_cluster_io_r_0_cluster_57_addr),
    .io_r_0_cluster_57_data(sram_cluster_io_r_0_cluster_57_data),
    .io_r_0_cluster_58_en(sram_cluster_io_r_0_cluster_58_en),
    .io_r_0_cluster_58_addr(sram_cluster_io_r_0_cluster_58_addr),
    .io_r_0_cluster_58_data(sram_cluster_io_r_0_cluster_58_data),
    .io_r_0_cluster_59_en(sram_cluster_io_r_0_cluster_59_en),
    .io_r_0_cluster_59_addr(sram_cluster_io_r_0_cluster_59_addr),
    .io_r_0_cluster_59_data(sram_cluster_io_r_0_cluster_59_data),
    .io_r_0_cluster_60_en(sram_cluster_io_r_0_cluster_60_en),
    .io_r_0_cluster_60_addr(sram_cluster_io_r_0_cluster_60_addr),
    .io_r_0_cluster_60_data(sram_cluster_io_r_0_cluster_60_data),
    .io_r_0_cluster_61_en(sram_cluster_io_r_0_cluster_61_en),
    .io_r_0_cluster_61_addr(sram_cluster_io_r_0_cluster_61_addr),
    .io_r_0_cluster_61_data(sram_cluster_io_r_0_cluster_61_data),
    .io_r_0_cluster_62_en(sram_cluster_io_r_0_cluster_62_en),
    .io_r_0_cluster_62_addr(sram_cluster_io_r_0_cluster_62_addr),
    .io_r_0_cluster_62_data(sram_cluster_io_r_0_cluster_62_data),
    .io_r_0_cluster_63_en(sram_cluster_io_r_0_cluster_63_en),
    .io_r_0_cluster_63_addr(sram_cluster_io_r_0_cluster_63_addr),
    .io_r_0_cluster_63_data(sram_cluster_io_r_0_cluster_63_data)
  );
  assign io_pipe_phv_out_data_0 = proc_io_pipe_phv_out_data_0; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_1 = proc_io_pipe_phv_out_data_1; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_2 = proc_io_pipe_phv_out_data_2; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_3 = proc_io_pipe_phv_out_data_3; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_4 = proc_io_pipe_phv_out_data_4; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_5 = proc_io_pipe_phv_out_data_5; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_6 = proc_io_pipe_phv_out_data_6; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_7 = proc_io_pipe_phv_out_data_7; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_8 = proc_io_pipe_phv_out_data_8; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_9 = proc_io_pipe_phv_out_data_9; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_10 = proc_io_pipe_phv_out_data_10; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_11 = proc_io_pipe_phv_out_data_11; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_12 = proc_io_pipe_phv_out_data_12; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_13 = proc_io_pipe_phv_out_data_13; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_14 = proc_io_pipe_phv_out_data_14; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_15 = proc_io_pipe_phv_out_data_15; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_16 = proc_io_pipe_phv_out_data_16; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_17 = proc_io_pipe_phv_out_data_17; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_18 = proc_io_pipe_phv_out_data_18; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_19 = proc_io_pipe_phv_out_data_19; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_20 = proc_io_pipe_phv_out_data_20; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_21 = proc_io_pipe_phv_out_data_21; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_22 = proc_io_pipe_phv_out_data_22; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_23 = proc_io_pipe_phv_out_data_23; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_24 = proc_io_pipe_phv_out_data_24; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_25 = proc_io_pipe_phv_out_data_25; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_26 = proc_io_pipe_phv_out_data_26; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_27 = proc_io_pipe_phv_out_data_27; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_28 = proc_io_pipe_phv_out_data_28; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_29 = proc_io_pipe_phv_out_data_29; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_30 = proc_io_pipe_phv_out_data_30; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_31 = proc_io_pipe_phv_out_data_31; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_32 = proc_io_pipe_phv_out_data_32; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_33 = proc_io_pipe_phv_out_data_33; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_34 = proc_io_pipe_phv_out_data_34; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_35 = proc_io_pipe_phv_out_data_35; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_36 = proc_io_pipe_phv_out_data_36; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_37 = proc_io_pipe_phv_out_data_37; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_38 = proc_io_pipe_phv_out_data_38; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_39 = proc_io_pipe_phv_out_data_39; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_40 = proc_io_pipe_phv_out_data_40; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_41 = proc_io_pipe_phv_out_data_41; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_42 = proc_io_pipe_phv_out_data_42; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_43 = proc_io_pipe_phv_out_data_43; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_44 = proc_io_pipe_phv_out_data_44; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_45 = proc_io_pipe_phv_out_data_45; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_46 = proc_io_pipe_phv_out_data_46; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_47 = proc_io_pipe_phv_out_data_47; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_48 = proc_io_pipe_phv_out_data_48; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_49 = proc_io_pipe_phv_out_data_49; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_50 = proc_io_pipe_phv_out_data_50; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_51 = proc_io_pipe_phv_out_data_51; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_52 = proc_io_pipe_phv_out_data_52; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_53 = proc_io_pipe_phv_out_data_53; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_54 = proc_io_pipe_phv_out_data_54; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_55 = proc_io_pipe_phv_out_data_55; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_56 = proc_io_pipe_phv_out_data_56; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_57 = proc_io_pipe_phv_out_data_57; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_58 = proc_io_pipe_phv_out_data_58; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_59 = proc_io_pipe_phv_out_data_59; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_60 = proc_io_pipe_phv_out_data_60; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_61 = proc_io_pipe_phv_out_data_61; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_62 = proc_io_pipe_phv_out_data_62; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_63 = proc_io_pipe_phv_out_data_63; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_64 = proc_io_pipe_phv_out_data_64; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_65 = proc_io_pipe_phv_out_data_65; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_66 = proc_io_pipe_phv_out_data_66; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_67 = proc_io_pipe_phv_out_data_67; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_68 = proc_io_pipe_phv_out_data_68; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_69 = proc_io_pipe_phv_out_data_69; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_70 = proc_io_pipe_phv_out_data_70; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_71 = proc_io_pipe_phv_out_data_71; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_72 = proc_io_pipe_phv_out_data_72; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_73 = proc_io_pipe_phv_out_data_73; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_74 = proc_io_pipe_phv_out_data_74; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_75 = proc_io_pipe_phv_out_data_75; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_76 = proc_io_pipe_phv_out_data_76; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_77 = proc_io_pipe_phv_out_data_77; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_78 = proc_io_pipe_phv_out_data_78; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_79 = proc_io_pipe_phv_out_data_79; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_80 = proc_io_pipe_phv_out_data_80; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_81 = proc_io_pipe_phv_out_data_81; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_82 = proc_io_pipe_phv_out_data_82; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_83 = proc_io_pipe_phv_out_data_83; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_84 = proc_io_pipe_phv_out_data_84; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_85 = proc_io_pipe_phv_out_data_85; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_86 = proc_io_pipe_phv_out_data_86; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_87 = proc_io_pipe_phv_out_data_87; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_88 = proc_io_pipe_phv_out_data_88; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_89 = proc_io_pipe_phv_out_data_89; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_90 = proc_io_pipe_phv_out_data_90; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_91 = proc_io_pipe_phv_out_data_91; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_92 = proc_io_pipe_phv_out_data_92; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_93 = proc_io_pipe_phv_out_data_93; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_94 = proc_io_pipe_phv_out_data_94; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_95 = proc_io_pipe_phv_out_data_95; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_96 = proc_io_pipe_phv_out_data_96; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_97 = proc_io_pipe_phv_out_data_97; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_98 = proc_io_pipe_phv_out_data_98; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_99 = proc_io_pipe_phv_out_data_99; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_100 = proc_io_pipe_phv_out_data_100; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_101 = proc_io_pipe_phv_out_data_101; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_102 = proc_io_pipe_phv_out_data_102; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_103 = proc_io_pipe_phv_out_data_103; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_104 = proc_io_pipe_phv_out_data_104; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_105 = proc_io_pipe_phv_out_data_105; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_106 = proc_io_pipe_phv_out_data_106; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_107 = proc_io_pipe_phv_out_data_107; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_108 = proc_io_pipe_phv_out_data_108; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_109 = proc_io_pipe_phv_out_data_109; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_110 = proc_io_pipe_phv_out_data_110; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_111 = proc_io_pipe_phv_out_data_111; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_112 = proc_io_pipe_phv_out_data_112; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_113 = proc_io_pipe_phv_out_data_113; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_114 = proc_io_pipe_phv_out_data_114; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_115 = proc_io_pipe_phv_out_data_115; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_116 = proc_io_pipe_phv_out_data_116; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_117 = proc_io_pipe_phv_out_data_117; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_118 = proc_io_pipe_phv_out_data_118; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_119 = proc_io_pipe_phv_out_data_119; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_120 = proc_io_pipe_phv_out_data_120; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_121 = proc_io_pipe_phv_out_data_121; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_122 = proc_io_pipe_phv_out_data_122; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_123 = proc_io_pipe_phv_out_data_123; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_124 = proc_io_pipe_phv_out_data_124; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_125 = proc_io_pipe_phv_out_data_125; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_126 = proc_io_pipe_phv_out_data_126; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_127 = proc_io_pipe_phv_out_data_127; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_128 = proc_io_pipe_phv_out_data_128; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_129 = proc_io_pipe_phv_out_data_129; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_130 = proc_io_pipe_phv_out_data_130; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_131 = proc_io_pipe_phv_out_data_131; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_132 = proc_io_pipe_phv_out_data_132; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_133 = proc_io_pipe_phv_out_data_133; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_134 = proc_io_pipe_phv_out_data_134; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_135 = proc_io_pipe_phv_out_data_135; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_136 = proc_io_pipe_phv_out_data_136; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_137 = proc_io_pipe_phv_out_data_137; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_138 = proc_io_pipe_phv_out_data_138; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_139 = proc_io_pipe_phv_out_data_139; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_140 = proc_io_pipe_phv_out_data_140; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_141 = proc_io_pipe_phv_out_data_141; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_142 = proc_io_pipe_phv_out_data_142; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_143 = proc_io_pipe_phv_out_data_143; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_144 = proc_io_pipe_phv_out_data_144; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_145 = proc_io_pipe_phv_out_data_145; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_146 = proc_io_pipe_phv_out_data_146; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_147 = proc_io_pipe_phv_out_data_147; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_148 = proc_io_pipe_phv_out_data_148; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_149 = proc_io_pipe_phv_out_data_149; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_150 = proc_io_pipe_phv_out_data_150; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_151 = proc_io_pipe_phv_out_data_151; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_152 = proc_io_pipe_phv_out_data_152; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_153 = proc_io_pipe_phv_out_data_153; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_154 = proc_io_pipe_phv_out_data_154; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_155 = proc_io_pipe_phv_out_data_155; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_156 = proc_io_pipe_phv_out_data_156; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_157 = proc_io_pipe_phv_out_data_157; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_158 = proc_io_pipe_phv_out_data_158; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_159 = proc_io_pipe_phv_out_data_159; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_160 = proc_io_pipe_phv_out_data_160; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_161 = proc_io_pipe_phv_out_data_161; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_162 = proc_io_pipe_phv_out_data_162; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_163 = proc_io_pipe_phv_out_data_163; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_164 = proc_io_pipe_phv_out_data_164; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_165 = proc_io_pipe_phv_out_data_165; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_166 = proc_io_pipe_phv_out_data_166; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_167 = proc_io_pipe_phv_out_data_167; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_168 = proc_io_pipe_phv_out_data_168; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_169 = proc_io_pipe_phv_out_data_169; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_170 = proc_io_pipe_phv_out_data_170; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_171 = proc_io_pipe_phv_out_data_171; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_172 = proc_io_pipe_phv_out_data_172; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_173 = proc_io_pipe_phv_out_data_173; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_174 = proc_io_pipe_phv_out_data_174; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_175 = proc_io_pipe_phv_out_data_175; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_176 = proc_io_pipe_phv_out_data_176; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_177 = proc_io_pipe_phv_out_data_177; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_178 = proc_io_pipe_phv_out_data_178; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_179 = proc_io_pipe_phv_out_data_179; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_180 = proc_io_pipe_phv_out_data_180; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_181 = proc_io_pipe_phv_out_data_181; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_182 = proc_io_pipe_phv_out_data_182; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_183 = proc_io_pipe_phv_out_data_183; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_184 = proc_io_pipe_phv_out_data_184; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_185 = proc_io_pipe_phv_out_data_185; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_186 = proc_io_pipe_phv_out_data_186; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_187 = proc_io_pipe_phv_out_data_187; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_188 = proc_io_pipe_phv_out_data_188; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_189 = proc_io_pipe_phv_out_data_189; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_190 = proc_io_pipe_phv_out_data_190; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_191 = proc_io_pipe_phv_out_data_191; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_192 = proc_io_pipe_phv_out_data_192; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_193 = proc_io_pipe_phv_out_data_193; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_194 = proc_io_pipe_phv_out_data_194; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_195 = proc_io_pipe_phv_out_data_195; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_196 = proc_io_pipe_phv_out_data_196; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_197 = proc_io_pipe_phv_out_data_197; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_198 = proc_io_pipe_phv_out_data_198; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_199 = proc_io_pipe_phv_out_data_199; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_200 = proc_io_pipe_phv_out_data_200; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_201 = proc_io_pipe_phv_out_data_201; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_202 = proc_io_pipe_phv_out_data_202; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_203 = proc_io_pipe_phv_out_data_203; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_204 = proc_io_pipe_phv_out_data_204; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_205 = proc_io_pipe_phv_out_data_205; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_206 = proc_io_pipe_phv_out_data_206; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_207 = proc_io_pipe_phv_out_data_207; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_208 = proc_io_pipe_phv_out_data_208; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_209 = proc_io_pipe_phv_out_data_209; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_210 = proc_io_pipe_phv_out_data_210; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_211 = proc_io_pipe_phv_out_data_211; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_212 = proc_io_pipe_phv_out_data_212; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_213 = proc_io_pipe_phv_out_data_213; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_214 = proc_io_pipe_phv_out_data_214; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_215 = proc_io_pipe_phv_out_data_215; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_216 = proc_io_pipe_phv_out_data_216; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_217 = proc_io_pipe_phv_out_data_217; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_218 = proc_io_pipe_phv_out_data_218; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_219 = proc_io_pipe_phv_out_data_219; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_220 = proc_io_pipe_phv_out_data_220; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_221 = proc_io_pipe_phv_out_data_221; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_222 = proc_io_pipe_phv_out_data_222; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_223 = proc_io_pipe_phv_out_data_223; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_224 = proc_io_pipe_phv_out_data_224; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_225 = proc_io_pipe_phv_out_data_225; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_226 = proc_io_pipe_phv_out_data_226; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_227 = proc_io_pipe_phv_out_data_227; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_228 = proc_io_pipe_phv_out_data_228; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_229 = proc_io_pipe_phv_out_data_229; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_230 = proc_io_pipe_phv_out_data_230; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_231 = proc_io_pipe_phv_out_data_231; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_232 = proc_io_pipe_phv_out_data_232; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_233 = proc_io_pipe_phv_out_data_233; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_234 = proc_io_pipe_phv_out_data_234; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_235 = proc_io_pipe_phv_out_data_235; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_236 = proc_io_pipe_phv_out_data_236; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_237 = proc_io_pipe_phv_out_data_237; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_238 = proc_io_pipe_phv_out_data_238; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_239 = proc_io_pipe_phv_out_data_239; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_240 = proc_io_pipe_phv_out_data_240; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_241 = proc_io_pipe_phv_out_data_241; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_242 = proc_io_pipe_phv_out_data_242; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_243 = proc_io_pipe_phv_out_data_243; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_244 = proc_io_pipe_phv_out_data_244; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_245 = proc_io_pipe_phv_out_data_245; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_246 = proc_io_pipe_phv_out_data_246; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_247 = proc_io_pipe_phv_out_data_247; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_248 = proc_io_pipe_phv_out_data_248; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_249 = proc_io_pipe_phv_out_data_249; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_250 = proc_io_pipe_phv_out_data_250; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_251 = proc_io_pipe_phv_out_data_251; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_252 = proc_io_pipe_phv_out_data_252; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_253 = proc_io_pipe_phv_out_data_253; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_254 = proc_io_pipe_phv_out_data_254; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_data_255 = proc_io_pipe_phv_out_data_255; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_header_0 = proc_io_pipe_phv_out_header_0; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_header_1 = proc_io_pipe_phv_out_header_1; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_header_2 = proc_io_pipe_phv_out_header_2; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_header_3 = proc_io_pipe_phv_out_header_3; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_header_4 = proc_io_pipe_phv_out_header_4; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_header_5 = proc_io_pipe_phv_out_header_5; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_header_6 = proc_io_pipe_phv_out_header_6; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_header_7 = proc_io_pipe_phv_out_header_7; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_header_8 = proc_io_pipe_phv_out_header_8; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_header_9 = proc_io_pipe_phv_out_header_9; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_header_10 = proc_io_pipe_phv_out_header_10; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_header_11 = proc_io_pipe_phv_out_header_11; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_header_12 = proc_io_pipe_phv_out_header_12; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_header_13 = proc_io_pipe_phv_out_header_13; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_header_14 = proc_io_pipe_phv_out_header_14; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_header_15 = proc_io_pipe_phv_out_header_15; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_parse_current_state = proc_io_pipe_phv_out_parse_current_state; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_parse_current_offset = proc_io_pipe_phv_out_parse_current_offset; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_parse_transition_field = proc_io_pipe_phv_out_parse_transition_field; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_next_processor_id = proc_io_pipe_phv_out_next_processor_id; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_next_config_id = proc_io_pipe_phv_out_next_config_id; // @[ipsa_single_processor.scala 16:26]
  assign io_pipe_phv_out_is_valid_processor = proc_io_pipe_phv_out_is_valid_processor; // @[ipsa_single_processor.scala 16:26]
  assign proc_clock = clock;
  assign proc_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_96 = io_pipe_phv_in_data_96; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_97 = io_pipe_phv_in_data_97; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_98 = io_pipe_phv_in_data_98; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_99 = io_pipe_phv_in_data_99; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_100 = io_pipe_phv_in_data_100; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_101 = io_pipe_phv_in_data_101; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_102 = io_pipe_phv_in_data_102; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_103 = io_pipe_phv_in_data_103; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_104 = io_pipe_phv_in_data_104; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_105 = io_pipe_phv_in_data_105; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_106 = io_pipe_phv_in_data_106; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_107 = io_pipe_phv_in_data_107; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_108 = io_pipe_phv_in_data_108; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_109 = io_pipe_phv_in_data_109; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_110 = io_pipe_phv_in_data_110; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_111 = io_pipe_phv_in_data_111; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_112 = io_pipe_phv_in_data_112; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_113 = io_pipe_phv_in_data_113; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_114 = io_pipe_phv_in_data_114; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_115 = io_pipe_phv_in_data_115; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_116 = io_pipe_phv_in_data_116; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_117 = io_pipe_phv_in_data_117; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_118 = io_pipe_phv_in_data_118; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_119 = io_pipe_phv_in_data_119; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_120 = io_pipe_phv_in_data_120; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_121 = io_pipe_phv_in_data_121; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_122 = io_pipe_phv_in_data_122; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_123 = io_pipe_phv_in_data_123; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_124 = io_pipe_phv_in_data_124; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_125 = io_pipe_phv_in_data_125; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_126 = io_pipe_phv_in_data_126; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_127 = io_pipe_phv_in_data_127; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_128 = io_pipe_phv_in_data_128; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_129 = io_pipe_phv_in_data_129; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_130 = io_pipe_phv_in_data_130; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_131 = io_pipe_phv_in_data_131; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_132 = io_pipe_phv_in_data_132; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_133 = io_pipe_phv_in_data_133; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_134 = io_pipe_phv_in_data_134; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_135 = io_pipe_phv_in_data_135; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_136 = io_pipe_phv_in_data_136; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_137 = io_pipe_phv_in_data_137; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_138 = io_pipe_phv_in_data_138; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_139 = io_pipe_phv_in_data_139; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_140 = io_pipe_phv_in_data_140; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_141 = io_pipe_phv_in_data_141; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_142 = io_pipe_phv_in_data_142; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_143 = io_pipe_phv_in_data_143; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_144 = io_pipe_phv_in_data_144; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_145 = io_pipe_phv_in_data_145; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_146 = io_pipe_phv_in_data_146; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_147 = io_pipe_phv_in_data_147; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_148 = io_pipe_phv_in_data_148; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_149 = io_pipe_phv_in_data_149; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_150 = io_pipe_phv_in_data_150; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_151 = io_pipe_phv_in_data_151; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_152 = io_pipe_phv_in_data_152; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_153 = io_pipe_phv_in_data_153; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_154 = io_pipe_phv_in_data_154; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_155 = io_pipe_phv_in_data_155; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_156 = io_pipe_phv_in_data_156; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_157 = io_pipe_phv_in_data_157; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_158 = io_pipe_phv_in_data_158; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_159 = io_pipe_phv_in_data_159; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_160 = io_pipe_phv_in_data_160; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_161 = io_pipe_phv_in_data_161; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_162 = io_pipe_phv_in_data_162; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_163 = io_pipe_phv_in_data_163; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_164 = io_pipe_phv_in_data_164; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_165 = io_pipe_phv_in_data_165; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_166 = io_pipe_phv_in_data_166; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_167 = io_pipe_phv_in_data_167; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_168 = io_pipe_phv_in_data_168; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_169 = io_pipe_phv_in_data_169; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_170 = io_pipe_phv_in_data_170; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_171 = io_pipe_phv_in_data_171; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_172 = io_pipe_phv_in_data_172; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_173 = io_pipe_phv_in_data_173; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_174 = io_pipe_phv_in_data_174; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_175 = io_pipe_phv_in_data_175; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_176 = io_pipe_phv_in_data_176; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_177 = io_pipe_phv_in_data_177; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_178 = io_pipe_phv_in_data_178; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_179 = io_pipe_phv_in_data_179; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_180 = io_pipe_phv_in_data_180; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_181 = io_pipe_phv_in_data_181; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_182 = io_pipe_phv_in_data_182; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_183 = io_pipe_phv_in_data_183; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_184 = io_pipe_phv_in_data_184; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_185 = io_pipe_phv_in_data_185; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_186 = io_pipe_phv_in_data_186; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_187 = io_pipe_phv_in_data_187; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_188 = io_pipe_phv_in_data_188; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_189 = io_pipe_phv_in_data_189; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_190 = io_pipe_phv_in_data_190; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_191 = io_pipe_phv_in_data_191; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_192 = io_pipe_phv_in_data_192; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_193 = io_pipe_phv_in_data_193; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_194 = io_pipe_phv_in_data_194; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_195 = io_pipe_phv_in_data_195; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_196 = io_pipe_phv_in_data_196; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_197 = io_pipe_phv_in_data_197; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_198 = io_pipe_phv_in_data_198; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_199 = io_pipe_phv_in_data_199; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_200 = io_pipe_phv_in_data_200; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_201 = io_pipe_phv_in_data_201; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_202 = io_pipe_phv_in_data_202; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_203 = io_pipe_phv_in_data_203; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_204 = io_pipe_phv_in_data_204; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_205 = io_pipe_phv_in_data_205; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_206 = io_pipe_phv_in_data_206; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_207 = io_pipe_phv_in_data_207; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_208 = io_pipe_phv_in_data_208; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_209 = io_pipe_phv_in_data_209; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_210 = io_pipe_phv_in_data_210; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_211 = io_pipe_phv_in_data_211; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_212 = io_pipe_phv_in_data_212; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_213 = io_pipe_phv_in_data_213; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_214 = io_pipe_phv_in_data_214; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_215 = io_pipe_phv_in_data_215; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_216 = io_pipe_phv_in_data_216; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_217 = io_pipe_phv_in_data_217; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_218 = io_pipe_phv_in_data_218; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_219 = io_pipe_phv_in_data_219; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_220 = io_pipe_phv_in_data_220; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_221 = io_pipe_phv_in_data_221; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_222 = io_pipe_phv_in_data_222; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_223 = io_pipe_phv_in_data_223; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_224 = io_pipe_phv_in_data_224; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_225 = io_pipe_phv_in_data_225; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_226 = io_pipe_phv_in_data_226; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_227 = io_pipe_phv_in_data_227; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_228 = io_pipe_phv_in_data_228; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_229 = io_pipe_phv_in_data_229; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_230 = io_pipe_phv_in_data_230; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_231 = io_pipe_phv_in_data_231; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_232 = io_pipe_phv_in_data_232; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_233 = io_pipe_phv_in_data_233; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_234 = io_pipe_phv_in_data_234; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_235 = io_pipe_phv_in_data_235; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_236 = io_pipe_phv_in_data_236; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_237 = io_pipe_phv_in_data_237; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_238 = io_pipe_phv_in_data_238; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_239 = io_pipe_phv_in_data_239; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_240 = io_pipe_phv_in_data_240; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_241 = io_pipe_phv_in_data_241; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_242 = io_pipe_phv_in_data_242; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_243 = io_pipe_phv_in_data_243; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_244 = io_pipe_phv_in_data_244; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_245 = io_pipe_phv_in_data_245; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_246 = io_pipe_phv_in_data_246; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_247 = io_pipe_phv_in_data_247; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_248 = io_pipe_phv_in_data_248; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_249 = io_pipe_phv_in_data_249; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_250 = io_pipe_phv_in_data_250; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_251 = io_pipe_phv_in_data_251; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_252 = io_pipe_phv_in_data_252; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_253 = io_pipe_phv_in_data_253; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_254 = io_pipe_phv_in_data_254; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_data_255 = io_pipe_phv_in_data_255; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_header_0 = io_pipe_phv_in_header_0; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_header_1 = io_pipe_phv_in_header_1; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_header_2 = io_pipe_phv_in_header_2; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_header_3 = io_pipe_phv_in_header_3; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_header_4 = io_pipe_phv_in_header_4; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_header_5 = io_pipe_phv_in_header_5; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_header_6 = io_pipe_phv_in_header_6; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_header_7 = io_pipe_phv_in_header_7; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_header_8 = io_pipe_phv_in_header_8; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_header_9 = io_pipe_phv_in_header_9; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_header_10 = io_pipe_phv_in_header_10; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_header_11 = io_pipe_phv_in_header_11; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_header_12 = io_pipe_phv_in_header_12; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_header_13 = io_pipe_phv_in_header_13; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_header_14 = io_pipe_phv_in_header_14; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_header_15 = io_pipe_phv_in_header_15; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_parse_current_state = io_pipe_phv_in_parse_current_state; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_parse_current_offset = io_pipe_phv_in_parse_current_offset; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_parse_transition_field = io_pipe_phv_in_parse_transition_field; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_next_processor_id = io_pipe_phv_in_next_processor_id; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_next_config_id = io_pipe_phv_in_next_config_id; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_pipe_phv_in_is_valid_processor = io_pipe_phv_in_is_valid_processor; // @[ipsa_single_processor.scala 15:25]
  assign proc_io_mod_par_mod_en = io_mod_par_mod_en; // @[ipsa_single_processor.scala 17:17]
  assign proc_io_mod_par_mod_last_mau_id_mod = io_mod_par_mod_last_mau_id_mod; // @[ipsa_single_processor.scala 17:17]
  assign proc_io_mod_par_mod_last_mau_id = io_mod_par_mod_last_mau_id; // @[ipsa_single_processor.scala 17:17]
  assign proc_io_mod_par_mod_cs = io_mod_par_mod_cs; // @[ipsa_single_processor.scala 17:17]
  assign proc_io_mod_par_mod_module_mod_state_id_mod = io_mod_par_mod_module_mod_state_id_mod; // @[ipsa_single_processor.scala 17:17]
  assign proc_io_mod_par_mod_module_mod_state_id = io_mod_par_mod_module_mod_state_id; // @[ipsa_single_processor.scala 17:17]
  assign proc_io_mod_par_mod_module_mod_sram_w_cs = io_mod_par_mod_module_mod_sram_w_cs; // @[ipsa_single_processor.scala 17:17]
  assign proc_io_mod_par_mod_module_mod_sram_w_en = io_mod_par_mod_module_mod_sram_w_en; // @[ipsa_single_processor.scala 17:17]
  assign proc_io_mod_par_mod_module_mod_sram_w_addr = io_mod_par_mod_module_mod_sram_w_addr; // @[ipsa_single_processor.scala 17:17]
  assign proc_io_mod_par_mod_module_mod_sram_w_data = io_mod_par_mod_module_mod_sram_w_data; // @[ipsa_single_processor.scala 17:17]
  assign proc_io_mod_mat_mod_en = io_mod_mat_mod_en; // @[ipsa_single_processor.scala 17:17]
  assign proc_io_mod_mat_mod_config_id = io_mod_mat_mod_config_id; // @[ipsa_single_processor.scala 17:17]
  assign proc_io_mod_mat_mod_key_mod_header_id = io_mod_mat_mod_key_mod_header_id; // @[ipsa_single_processor.scala 17:17]
  assign proc_io_mod_mat_mod_key_mod_internal_offset = io_mod_mat_mod_key_mod_internal_offset; // @[ipsa_single_processor.scala 17:17]
  assign proc_io_mod_mat_mod_key_mod_key_length = io_mod_mat_mod_key_mod_key_length; // @[ipsa_single_processor.scala 17:17]
  assign proc_io_mod_mat_mod_table_mod_table_width = io_mod_mat_mod_table_mod_table_width; // @[ipsa_single_processor.scala 17:17]
  assign proc_io_mod_mat_mod_table_mod_table_depth = io_mod_mat_mod_table_mod_table_depth; // @[ipsa_single_processor.scala 17:17]
  assign proc_io_mod_act_mod_en_0 = io_mod_act_mod_en_0; // @[ipsa_single_processor.scala 17:17]
  assign proc_io_mod_act_mod_en_1 = io_mod_act_mod_en_1; // @[ipsa_single_processor.scala 17:17]
  assign proc_io_mod_act_mod_addr = io_mod_act_mod_addr; // @[ipsa_single_processor.scala 17:17]
  assign proc_io_mod_act_mod_data_0 = io_mod_act_mod_data_0; // @[ipsa_single_processor.scala 17:17]
  assign proc_io_mod_act_mod_data_1 = io_mod_act_mod_data_1; // @[ipsa_single_processor.scala 17:17]
  assign proc_io_mem_cluster_0_data = sram_cluster_io_r_0_cluster_0_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_1_data = sram_cluster_io_r_0_cluster_1_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_2_data = sram_cluster_io_r_0_cluster_2_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_3_data = sram_cluster_io_r_0_cluster_3_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_4_data = sram_cluster_io_r_0_cluster_4_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_5_data = sram_cluster_io_r_0_cluster_5_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_6_data = sram_cluster_io_r_0_cluster_6_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_7_data = sram_cluster_io_r_0_cluster_7_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_8_data = sram_cluster_io_r_0_cluster_8_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_9_data = sram_cluster_io_r_0_cluster_9_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_10_data = sram_cluster_io_r_0_cluster_10_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_11_data = sram_cluster_io_r_0_cluster_11_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_12_data = sram_cluster_io_r_0_cluster_12_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_13_data = sram_cluster_io_r_0_cluster_13_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_14_data = sram_cluster_io_r_0_cluster_14_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_15_data = sram_cluster_io_r_0_cluster_15_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_16_data = sram_cluster_io_r_0_cluster_16_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_17_data = sram_cluster_io_r_0_cluster_17_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_18_data = sram_cluster_io_r_0_cluster_18_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_19_data = sram_cluster_io_r_0_cluster_19_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_20_data = sram_cluster_io_r_0_cluster_20_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_21_data = sram_cluster_io_r_0_cluster_21_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_22_data = sram_cluster_io_r_0_cluster_22_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_23_data = sram_cluster_io_r_0_cluster_23_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_24_data = sram_cluster_io_r_0_cluster_24_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_25_data = sram_cluster_io_r_0_cluster_25_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_26_data = sram_cluster_io_r_0_cluster_26_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_27_data = sram_cluster_io_r_0_cluster_27_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_28_data = sram_cluster_io_r_0_cluster_28_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_29_data = sram_cluster_io_r_0_cluster_29_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_30_data = sram_cluster_io_r_0_cluster_30_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_31_data = sram_cluster_io_r_0_cluster_31_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_32_data = sram_cluster_io_r_0_cluster_32_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_33_data = sram_cluster_io_r_0_cluster_33_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_34_data = sram_cluster_io_r_0_cluster_34_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_35_data = sram_cluster_io_r_0_cluster_35_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_36_data = sram_cluster_io_r_0_cluster_36_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_37_data = sram_cluster_io_r_0_cluster_37_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_38_data = sram_cluster_io_r_0_cluster_38_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_39_data = sram_cluster_io_r_0_cluster_39_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_40_data = sram_cluster_io_r_0_cluster_40_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_41_data = sram_cluster_io_r_0_cluster_41_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_42_data = sram_cluster_io_r_0_cluster_42_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_43_data = sram_cluster_io_r_0_cluster_43_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_44_data = sram_cluster_io_r_0_cluster_44_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_45_data = sram_cluster_io_r_0_cluster_45_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_46_data = sram_cluster_io_r_0_cluster_46_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_47_data = sram_cluster_io_r_0_cluster_47_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_48_data = sram_cluster_io_r_0_cluster_48_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_49_data = sram_cluster_io_r_0_cluster_49_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_50_data = sram_cluster_io_r_0_cluster_50_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_51_data = sram_cluster_io_r_0_cluster_51_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_52_data = sram_cluster_io_r_0_cluster_52_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_53_data = sram_cluster_io_r_0_cluster_53_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_54_data = sram_cluster_io_r_0_cluster_54_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_55_data = sram_cluster_io_r_0_cluster_55_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_56_data = sram_cluster_io_r_0_cluster_56_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_57_data = sram_cluster_io_r_0_cluster_57_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_58_data = sram_cluster_io_r_0_cluster_58_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_59_data = sram_cluster_io_r_0_cluster_59_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_60_data = sram_cluster_io_r_0_cluster_60_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_61_data = sram_cluster_io_r_0_cluster_61_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_62_data = sram_cluster_io_r_0_cluster_62_data; // @[ipsa_single_processor.scala 21:26]
  assign proc_io_mem_cluster_63_data = sram_cluster_io_r_0_cluster_63_data; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_clock = clock;
  assign sram_cluster_io_w_wcs = io_w_wcs; // @[ipsa_single_processor.scala 20:23]
  assign sram_cluster_io_w_w_en = io_w_w_en; // @[ipsa_single_processor.scala 20:23]
  assign sram_cluster_io_w_w_addr = io_w_w_addr; // @[ipsa_single_processor.scala 20:23]
  assign sram_cluster_io_w_w_data = io_w_w_data; // @[ipsa_single_processor.scala 20:23]
  assign sram_cluster_io_r_0_cluster_0_en = proc_io_mem_cluster_0_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_0_addr = proc_io_mem_cluster_0_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_1_en = proc_io_mem_cluster_1_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_1_addr = proc_io_mem_cluster_1_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_2_en = proc_io_mem_cluster_2_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_2_addr = proc_io_mem_cluster_2_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_3_en = proc_io_mem_cluster_3_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_3_addr = proc_io_mem_cluster_3_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_4_en = proc_io_mem_cluster_4_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_4_addr = proc_io_mem_cluster_4_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_5_en = proc_io_mem_cluster_5_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_5_addr = proc_io_mem_cluster_5_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_6_en = proc_io_mem_cluster_6_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_6_addr = proc_io_mem_cluster_6_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_7_en = proc_io_mem_cluster_7_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_7_addr = proc_io_mem_cluster_7_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_8_en = proc_io_mem_cluster_8_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_8_addr = proc_io_mem_cluster_8_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_9_en = proc_io_mem_cluster_9_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_9_addr = proc_io_mem_cluster_9_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_10_en = proc_io_mem_cluster_10_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_10_addr = proc_io_mem_cluster_10_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_11_en = proc_io_mem_cluster_11_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_11_addr = proc_io_mem_cluster_11_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_12_en = proc_io_mem_cluster_12_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_12_addr = proc_io_mem_cluster_12_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_13_en = proc_io_mem_cluster_13_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_13_addr = proc_io_mem_cluster_13_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_14_en = proc_io_mem_cluster_14_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_14_addr = proc_io_mem_cluster_14_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_15_en = proc_io_mem_cluster_15_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_15_addr = proc_io_mem_cluster_15_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_16_en = proc_io_mem_cluster_16_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_16_addr = proc_io_mem_cluster_16_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_17_en = proc_io_mem_cluster_17_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_17_addr = proc_io_mem_cluster_17_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_18_en = proc_io_mem_cluster_18_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_18_addr = proc_io_mem_cluster_18_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_19_en = proc_io_mem_cluster_19_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_19_addr = proc_io_mem_cluster_19_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_20_en = proc_io_mem_cluster_20_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_20_addr = proc_io_mem_cluster_20_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_21_en = proc_io_mem_cluster_21_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_21_addr = proc_io_mem_cluster_21_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_22_en = proc_io_mem_cluster_22_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_22_addr = proc_io_mem_cluster_22_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_23_en = proc_io_mem_cluster_23_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_23_addr = proc_io_mem_cluster_23_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_24_en = proc_io_mem_cluster_24_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_24_addr = proc_io_mem_cluster_24_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_25_en = proc_io_mem_cluster_25_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_25_addr = proc_io_mem_cluster_25_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_26_en = proc_io_mem_cluster_26_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_26_addr = proc_io_mem_cluster_26_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_27_en = proc_io_mem_cluster_27_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_27_addr = proc_io_mem_cluster_27_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_28_en = proc_io_mem_cluster_28_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_28_addr = proc_io_mem_cluster_28_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_29_en = proc_io_mem_cluster_29_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_29_addr = proc_io_mem_cluster_29_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_30_en = proc_io_mem_cluster_30_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_30_addr = proc_io_mem_cluster_30_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_31_en = proc_io_mem_cluster_31_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_31_addr = proc_io_mem_cluster_31_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_32_en = proc_io_mem_cluster_32_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_32_addr = proc_io_mem_cluster_32_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_33_en = proc_io_mem_cluster_33_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_33_addr = proc_io_mem_cluster_33_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_34_en = proc_io_mem_cluster_34_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_34_addr = proc_io_mem_cluster_34_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_35_en = proc_io_mem_cluster_35_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_35_addr = proc_io_mem_cluster_35_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_36_en = proc_io_mem_cluster_36_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_36_addr = proc_io_mem_cluster_36_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_37_en = proc_io_mem_cluster_37_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_37_addr = proc_io_mem_cluster_37_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_38_en = proc_io_mem_cluster_38_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_38_addr = proc_io_mem_cluster_38_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_39_en = proc_io_mem_cluster_39_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_39_addr = proc_io_mem_cluster_39_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_40_en = proc_io_mem_cluster_40_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_40_addr = proc_io_mem_cluster_40_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_41_en = proc_io_mem_cluster_41_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_41_addr = proc_io_mem_cluster_41_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_42_en = proc_io_mem_cluster_42_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_42_addr = proc_io_mem_cluster_42_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_43_en = proc_io_mem_cluster_43_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_43_addr = proc_io_mem_cluster_43_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_44_en = proc_io_mem_cluster_44_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_44_addr = proc_io_mem_cluster_44_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_45_en = proc_io_mem_cluster_45_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_45_addr = proc_io_mem_cluster_45_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_46_en = proc_io_mem_cluster_46_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_46_addr = proc_io_mem_cluster_46_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_47_en = proc_io_mem_cluster_47_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_47_addr = proc_io_mem_cluster_47_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_48_en = proc_io_mem_cluster_48_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_48_addr = proc_io_mem_cluster_48_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_49_en = proc_io_mem_cluster_49_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_49_addr = proc_io_mem_cluster_49_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_50_en = proc_io_mem_cluster_50_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_50_addr = proc_io_mem_cluster_50_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_51_en = proc_io_mem_cluster_51_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_51_addr = proc_io_mem_cluster_51_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_52_en = proc_io_mem_cluster_52_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_52_addr = proc_io_mem_cluster_52_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_53_en = proc_io_mem_cluster_53_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_53_addr = proc_io_mem_cluster_53_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_54_en = proc_io_mem_cluster_54_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_54_addr = proc_io_mem_cluster_54_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_55_en = proc_io_mem_cluster_55_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_55_addr = proc_io_mem_cluster_55_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_56_en = proc_io_mem_cluster_56_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_56_addr = proc_io_mem_cluster_56_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_57_en = proc_io_mem_cluster_57_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_57_addr = proc_io_mem_cluster_57_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_58_en = proc_io_mem_cluster_58_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_58_addr = proc_io_mem_cluster_58_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_59_en = proc_io_mem_cluster_59_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_59_addr = proc_io_mem_cluster_59_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_60_en = proc_io_mem_cluster_60_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_60_addr = proc_io_mem_cluster_60_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_61_en = proc_io_mem_cluster_61_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_61_addr = proc_io_mem_cluster_61_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_62_en = proc_io_mem_cluster_62_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_62_addr = proc_io_mem_cluster_62_addr; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_63_en = proc_io_mem_cluster_63_en; // @[ipsa_single_processor.scala 21:26]
  assign sram_cluster_io_r_0_cluster_63_addr = proc_io_mem_cluster_63_addr; // @[ipsa_single_processor.scala 21:26]
endmodule
