module ProcessorPISA(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [7:0]  io_pipe_phv_in_data_160,
  input  [7:0]  io_pipe_phv_in_data_161,
  input  [7:0]  io_pipe_phv_in_data_162,
  input  [7:0]  io_pipe_phv_in_data_163,
  input  [7:0]  io_pipe_phv_in_data_164,
  input  [7:0]  io_pipe_phv_in_data_165,
  input  [7:0]  io_pipe_phv_in_data_166,
  input  [7:0]  io_pipe_phv_in_data_167,
  input  [7:0]  io_pipe_phv_in_data_168,
  input  [7:0]  io_pipe_phv_in_data_169,
  input  [7:0]  io_pipe_phv_in_data_170,
  input  [7:0]  io_pipe_phv_in_data_171,
  input  [7:0]  io_pipe_phv_in_data_172,
  input  [7:0]  io_pipe_phv_in_data_173,
  input  [7:0]  io_pipe_phv_in_data_174,
  input  [7:0]  io_pipe_phv_in_data_175,
  input  [7:0]  io_pipe_phv_in_data_176,
  input  [7:0]  io_pipe_phv_in_data_177,
  input  [7:0]  io_pipe_phv_in_data_178,
  input  [7:0]  io_pipe_phv_in_data_179,
  input  [7:0]  io_pipe_phv_in_data_180,
  input  [7:0]  io_pipe_phv_in_data_181,
  input  [7:0]  io_pipe_phv_in_data_182,
  input  [7:0]  io_pipe_phv_in_data_183,
  input  [7:0]  io_pipe_phv_in_data_184,
  input  [7:0]  io_pipe_phv_in_data_185,
  input  [7:0]  io_pipe_phv_in_data_186,
  input  [7:0]  io_pipe_phv_in_data_187,
  input  [7:0]  io_pipe_phv_in_data_188,
  input  [7:0]  io_pipe_phv_in_data_189,
  input  [7:0]  io_pipe_phv_in_data_190,
  input  [7:0]  io_pipe_phv_in_data_191,
  input  [7:0]  io_pipe_phv_in_data_192,
  input  [7:0]  io_pipe_phv_in_data_193,
  input  [7:0]  io_pipe_phv_in_data_194,
  input  [7:0]  io_pipe_phv_in_data_195,
  input  [7:0]  io_pipe_phv_in_data_196,
  input  [7:0]  io_pipe_phv_in_data_197,
  input  [7:0]  io_pipe_phv_in_data_198,
  input  [7:0]  io_pipe_phv_in_data_199,
  input  [7:0]  io_pipe_phv_in_data_200,
  input  [7:0]  io_pipe_phv_in_data_201,
  input  [7:0]  io_pipe_phv_in_data_202,
  input  [7:0]  io_pipe_phv_in_data_203,
  input  [7:0]  io_pipe_phv_in_data_204,
  input  [7:0]  io_pipe_phv_in_data_205,
  input  [7:0]  io_pipe_phv_in_data_206,
  input  [7:0]  io_pipe_phv_in_data_207,
  input  [7:0]  io_pipe_phv_in_data_208,
  input  [7:0]  io_pipe_phv_in_data_209,
  input  [7:0]  io_pipe_phv_in_data_210,
  input  [7:0]  io_pipe_phv_in_data_211,
  input  [7:0]  io_pipe_phv_in_data_212,
  input  [7:0]  io_pipe_phv_in_data_213,
  input  [7:0]  io_pipe_phv_in_data_214,
  input  [7:0]  io_pipe_phv_in_data_215,
  input  [7:0]  io_pipe_phv_in_data_216,
  input  [7:0]  io_pipe_phv_in_data_217,
  input  [7:0]  io_pipe_phv_in_data_218,
  input  [7:0]  io_pipe_phv_in_data_219,
  input  [7:0]  io_pipe_phv_in_data_220,
  input  [7:0]  io_pipe_phv_in_data_221,
  input  [7:0]  io_pipe_phv_in_data_222,
  input  [7:0]  io_pipe_phv_in_data_223,
  input  [7:0]  io_pipe_phv_in_data_224,
  input  [7:0]  io_pipe_phv_in_data_225,
  input  [7:0]  io_pipe_phv_in_data_226,
  input  [7:0]  io_pipe_phv_in_data_227,
  input  [7:0]  io_pipe_phv_in_data_228,
  input  [7:0]  io_pipe_phv_in_data_229,
  input  [7:0]  io_pipe_phv_in_data_230,
  input  [7:0]  io_pipe_phv_in_data_231,
  input  [7:0]  io_pipe_phv_in_data_232,
  input  [7:0]  io_pipe_phv_in_data_233,
  input  [7:0]  io_pipe_phv_in_data_234,
  input  [7:0]  io_pipe_phv_in_data_235,
  input  [7:0]  io_pipe_phv_in_data_236,
  input  [7:0]  io_pipe_phv_in_data_237,
  input  [7:0]  io_pipe_phv_in_data_238,
  input  [7:0]  io_pipe_phv_in_data_239,
  input  [7:0]  io_pipe_phv_in_data_240,
  input  [7:0]  io_pipe_phv_in_data_241,
  input  [7:0]  io_pipe_phv_in_data_242,
  input  [7:0]  io_pipe_phv_in_data_243,
  input  [7:0]  io_pipe_phv_in_data_244,
  input  [7:0]  io_pipe_phv_in_data_245,
  input  [7:0]  io_pipe_phv_in_data_246,
  input  [7:0]  io_pipe_phv_in_data_247,
  input  [7:0]  io_pipe_phv_in_data_248,
  input  [7:0]  io_pipe_phv_in_data_249,
  input  [7:0]  io_pipe_phv_in_data_250,
  input  [7:0]  io_pipe_phv_in_data_251,
  input  [7:0]  io_pipe_phv_in_data_252,
  input  [7:0]  io_pipe_phv_in_data_253,
  input  [7:0]  io_pipe_phv_in_data_254,
  input  [7:0]  io_pipe_phv_in_data_255,
  input  [3:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [7:0]  io_pipe_phv_out_data_160,
  output [7:0]  io_pipe_phv_out_data_161,
  output [7:0]  io_pipe_phv_out_data_162,
  output [7:0]  io_pipe_phv_out_data_163,
  output [7:0]  io_pipe_phv_out_data_164,
  output [7:0]  io_pipe_phv_out_data_165,
  output [7:0]  io_pipe_phv_out_data_166,
  output [7:0]  io_pipe_phv_out_data_167,
  output [7:0]  io_pipe_phv_out_data_168,
  output [7:0]  io_pipe_phv_out_data_169,
  output [7:0]  io_pipe_phv_out_data_170,
  output [7:0]  io_pipe_phv_out_data_171,
  output [7:0]  io_pipe_phv_out_data_172,
  output [7:0]  io_pipe_phv_out_data_173,
  output [7:0]  io_pipe_phv_out_data_174,
  output [7:0]  io_pipe_phv_out_data_175,
  output [7:0]  io_pipe_phv_out_data_176,
  output [7:0]  io_pipe_phv_out_data_177,
  output [7:0]  io_pipe_phv_out_data_178,
  output [7:0]  io_pipe_phv_out_data_179,
  output [7:0]  io_pipe_phv_out_data_180,
  output [7:0]  io_pipe_phv_out_data_181,
  output [7:0]  io_pipe_phv_out_data_182,
  output [7:0]  io_pipe_phv_out_data_183,
  output [7:0]  io_pipe_phv_out_data_184,
  output [7:0]  io_pipe_phv_out_data_185,
  output [7:0]  io_pipe_phv_out_data_186,
  output [7:0]  io_pipe_phv_out_data_187,
  output [7:0]  io_pipe_phv_out_data_188,
  output [7:0]  io_pipe_phv_out_data_189,
  output [7:0]  io_pipe_phv_out_data_190,
  output [7:0]  io_pipe_phv_out_data_191,
  output [7:0]  io_pipe_phv_out_data_192,
  output [7:0]  io_pipe_phv_out_data_193,
  output [7:0]  io_pipe_phv_out_data_194,
  output [7:0]  io_pipe_phv_out_data_195,
  output [7:0]  io_pipe_phv_out_data_196,
  output [7:0]  io_pipe_phv_out_data_197,
  output [7:0]  io_pipe_phv_out_data_198,
  output [7:0]  io_pipe_phv_out_data_199,
  output [7:0]  io_pipe_phv_out_data_200,
  output [7:0]  io_pipe_phv_out_data_201,
  output [7:0]  io_pipe_phv_out_data_202,
  output [7:0]  io_pipe_phv_out_data_203,
  output [7:0]  io_pipe_phv_out_data_204,
  output [7:0]  io_pipe_phv_out_data_205,
  output [7:0]  io_pipe_phv_out_data_206,
  output [7:0]  io_pipe_phv_out_data_207,
  output [7:0]  io_pipe_phv_out_data_208,
  output [7:0]  io_pipe_phv_out_data_209,
  output [7:0]  io_pipe_phv_out_data_210,
  output [7:0]  io_pipe_phv_out_data_211,
  output [7:0]  io_pipe_phv_out_data_212,
  output [7:0]  io_pipe_phv_out_data_213,
  output [7:0]  io_pipe_phv_out_data_214,
  output [7:0]  io_pipe_phv_out_data_215,
  output [7:0]  io_pipe_phv_out_data_216,
  output [7:0]  io_pipe_phv_out_data_217,
  output [7:0]  io_pipe_phv_out_data_218,
  output [7:0]  io_pipe_phv_out_data_219,
  output [7:0]  io_pipe_phv_out_data_220,
  output [7:0]  io_pipe_phv_out_data_221,
  output [7:0]  io_pipe_phv_out_data_222,
  output [7:0]  io_pipe_phv_out_data_223,
  output [7:0]  io_pipe_phv_out_data_224,
  output [7:0]  io_pipe_phv_out_data_225,
  output [7:0]  io_pipe_phv_out_data_226,
  output [7:0]  io_pipe_phv_out_data_227,
  output [7:0]  io_pipe_phv_out_data_228,
  output [7:0]  io_pipe_phv_out_data_229,
  output [7:0]  io_pipe_phv_out_data_230,
  output [7:0]  io_pipe_phv_out_data_231,
  output [7:0]  io_pipe_phv_out_data_232,
  output [7:0]  io_pipe_phv_out_data_233,
  output [7:0]  io_pipe_phv_out_data_234,
  output [7:0]  io_pipe_phv_out_data_235,
  output [7:0]  io_pipe_phv_out_data_236,
  output [7:0]  io_pipe_phv_out_data_237,
  output [7:0]  io_pipe_phv_out_data_238,
  output [7:0]  io_pipe_phv_out_data_239,
  output [7:0]  io_pipe_phv_out_data_240,
  output [7:0]  io_pipe_phv_out_data_241,
  output [7:0]  io_pipe_phv_out_data_242,
  output [7:0]  io_pipe_phv_out_data_243,
  output [7:0]  io_pipe_phv_out_data_244,
  output [7:0]  io_pipe_phv_out_data_245,
  output [7:0]  io_pipe_phv_out_data_246,
  output [7:0]  io_pipe_phv_out_data_247,
  output [7:0]  io_pipe_phv_out_data_248,
  output [7:0]  io_pipe_phv_out_data_249,
  output [7:0]  io_pipe_phv_out_data_250,
  output [7:0]  io_pipe_phv_out_data_251,
  output [7:0]  io_pipe_phv_out_data_252,
  output [7:0]  io_pipe_phv_out_data_253,
  output [7:0]  io_pipe_phv_out_data_254,
  output [7:0]  io_pipe_phv_out_data_255,
  output [3:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  input         io_mod_mat_mod_en,
  input         io_mod_mat_mod_config_id,
  input         io_mod_mat_mod_key_mod_en,
  input  [2:0]  io_mod_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_mat_mod_key_mod_group_config,
  input         io_mod_mat_mod_key_mod_group_mask_0,
  input         io_mod_mat_mod_key_mod_group_mask_1,
  input         io_mod_mat_mod_key_mod_group_mask_2,
  input         io_mod_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_mat_mod_table_mod_table_width,
  input         io_mod_mat_mod_w_en,
  input  [3:0]  io_mod_mat_mod_w_sram_id,
  input  [7:0]  io_mod_mat_mod_w_addr,
  input  [63:0] io_mod_mat_mod_w_data,
  input         io_mod_exe_mod_en_0,
  input         io_mod_exe_mod_en_1,
  input  [7:0]  io_mod_exe_mod_addr,
  input  [63:0] io_mod_exe_mod_data_0,
  input  [63:0] io_mod_exe_mod_data_1
);
  wire  MAT_clock; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_0; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_1; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_2; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_3; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_4; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_5; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_6; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_7; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_8; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_9; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_10; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_11; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_12; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_13; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_14; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_15; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_16; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_17; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_18; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_19; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_20; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_21; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_22; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_23; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_24; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_25; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_26; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_27; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_28; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_29; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_30; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_31; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_32; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_33; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_34; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_35; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_36; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_37; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_38; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_39; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_40; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_41; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_42; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_43; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_44; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_45; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_46; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_47; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_48; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_49; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_50; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_51; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_52; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_53; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_54; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_55; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_56; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_57; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_58; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_59; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_60; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_61; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_62; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_63; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_64; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_65; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_66; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_67; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_68; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_69; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_70; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_71; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_72; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_73; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_74; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_75; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_76; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_77; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_78; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_79; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_80; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_81; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_82; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_83; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_84; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_85; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_86; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_87; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_88; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_89; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_90; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_91; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_92; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_93; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_94; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_95; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_96; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_97; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_98; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_99; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_100; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_101; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_102; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_103; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_104; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_105; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_106; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_107; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_108; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_109; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_110; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_111; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_112; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_113; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_114; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_115; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_116; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_117; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_118; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_119; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_120; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_121; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_122; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_123; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_124; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_125; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_126; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_127; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_128; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_129; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_130; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_131; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_132; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_133; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_134; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_135; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_136; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_137; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_138; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_139; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_140; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_141; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_142; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_143; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_144; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_145; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_146; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_147; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_148; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_149; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_150; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_151; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_152; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_153; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_154; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_155; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_156; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_157; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_158; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_159; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_160; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_161; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_162; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_163; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_164; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_165; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_166; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_167; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_168; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_169; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_170; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_171; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_172; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_173; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_174; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_175; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_176; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_177; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_178; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_179; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_180; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_181; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_182; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_183; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_184; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_185; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_186; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_187; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_188; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_189; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_190; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_191; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_192; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_193; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_194; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_195; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_196; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_197; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_198; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_199; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_200; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_201; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_202; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_203; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_204; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_205; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_206; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_207; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_208; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_209; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_210; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_211; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_212; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_213; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_214; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_215; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_216; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_217; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_218; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_219; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_220; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_221; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_222; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_223; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_224; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_225; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_226; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_227; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_228; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_229; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_230; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_231; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_232; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_233; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_234; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_235; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_236; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_237; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_238; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_239; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_240; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_241; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_242; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_243; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_244; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_245; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_246; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_247; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_248; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_249; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_250; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_251; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_252; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_253; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_254; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_in_data_255; // @[processor_pisa.scala 19:21]
  wire [3:0] MAT_io_pipe_phv_in_next_processor_id; // @[processor_pisa.scala 19:21]
  wire  MAT_io_pipe_phv_in_next_config_id; // @[processor_pisa.scala 19:21]
  wire  MAT_io_pipe_phv_in_is_valid_processor; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_0; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_1; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_2; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_3; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_4; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_5; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_6; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_7; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_8; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_9; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_10; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_11; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_12; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_13; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_14; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_15; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_16; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_17; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_18; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_19; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_20; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_21; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_22; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_23; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_24; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_25; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_26; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_27; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_28; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_29; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_30; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_31; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_32; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_33; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_34; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_35; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_36; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_37; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_38; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_39; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_40; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_41; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_42; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_43; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_44; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_45; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_46; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_47; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_48; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_49; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_50; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_51; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_52; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_53; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_54; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_55; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_56; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_57; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_58; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_59; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_60; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_61; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_62; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_63; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_64; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_65; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_66; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_67; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_68; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_69; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_70; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_71; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_72; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_73; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_74; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_75; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_76; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_77; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_78; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_79; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_80; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_81; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_82; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_83; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_84; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_85; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_86; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_87; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_88; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_89; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_90; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_91; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_92; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_93; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_94; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_95; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_96; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_97; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_98; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_99; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_100; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_101; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_102; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_103; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_104; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_105; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_106; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_107; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_108; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_109; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_110; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_111; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_112; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_113; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_114; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_115; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_116; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_117; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_118; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_119; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_120; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_121; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_122; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_123; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_124; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_125; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_126; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_127; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_128; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_129; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_130; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_131; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_132; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_133; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_134; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_135; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_136; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_137; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_138; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_139; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_140; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_141; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_142; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_143; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_144; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_145; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_146; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_147; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_148; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_149; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_150; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_151; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_152; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_153; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_154; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_155; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_156; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_157; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_158; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_159; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_160; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_161; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_162; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_163; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_164; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_165; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_166; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_167; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_168; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_169; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_170; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_171; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_172; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_173; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_174; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_175; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_176; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_177; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_178; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_179; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_180; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_181; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_182; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_183; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_184; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_185; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_186; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_187; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_188; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_189; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_190; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_191; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_192; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_193; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_194; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_195; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_196; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_197; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_198; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_199; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_200; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_201; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_202; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_203; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_204; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_205; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_206; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_207; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_208; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_209; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_210; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_211; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_212; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_213; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_214; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_215; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_216; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_217; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_218; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_219; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_220; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_221; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_222; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_223; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_224; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_225; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_226; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_227; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_228; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_229; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_230; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_231; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_232; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_233; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_234; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_235; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_236; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_237; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_238; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_239; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_240; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_241; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_242; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_243; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_244; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_245; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_246; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_247; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_248; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_249; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_250; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_251; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_252; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_253; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_254; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_pipe_phv_out_data_255; // @[processor_pisa.scala 19:21]
  wire [3:0] MAT_io_pipe_phv_out_next_processor_id; // @[processor_pisa.scala 19:21]
  wire  MAT_io_pipe_phv_out_next_config_id; // @[processor_pisa.scala 19:21]
  wire  MAT_io_pipe_phv_out_is_valid_processor; // @[processor_pisa.scala 19:21]
  wire  MAT_io_mod_en; // @[processor_pisa.scala 19:21]
  wire  MAT_io_mod_config_id; // @[processor_pisa.scala 19:21]
  wire  MAT_io_mod_key_mod_en; // @[processor_pisa.scala 19:21]
  wire [2:0] MAT_io_mod_key_mod_group_index; // @[processor_pisa.scala 19:21]
  wire [1:0] MAT_io_mod_key_mod_group_config; // @[processor_pisa.scala 19:21]
  wire  MAT_io_mod_key_mod_group_mask_0; // @[processor_pisa.scala 19:21]
  wire  MAT_io_mod_key_mod_group_mask_1; // @[processor_pisa.scala 19:21]
  wire  MAT_io_mod_key_mod_group_mask_2; // @[processor_pisa.scala 19:21]
  wire  MAT_io_mod_key_mod_group_mask_3; // @[processor_pisa.scala 19:21]
  wire [6:0] MAT_io_mod_key_mod_group_id_0; // @[processor_pisa.scala 19:21]
  wire [6:0] MAT_io_mod_key_mod_group_id_1; // @[processor_pisa.scala 19:21]
  wire [6:0] MAT_io_mod_key_mod_group_id_2; // @[processor_pisa.scala 19:21]
  wire [6:0] MAT_io_mod_key_mod_group_id_3; // @[processor_pisa.scala 19:21]
  wire [4:0] MAT_io_mod_table_mod_table_depth; // @[processor_pisa.scala 19:21]
  wire [4:0] MAT_io_mod_table_mod_table_width; // @[processor_pisa.scala 19:21]
  wire  MAT_io_mod_w_en; // @[processor_pisa.scala 19:21]
  wire [3:0] MAT_io_mod_w_sram_id; // @[processor_pisa.scala 19:21]
  wire [7:0] MAT_io_mod_w_addr; // @[processor_pisa.scala 19:21]
  wire [63:0] MAT_io_mod_w_data; // @[processor_pisa.scala 19:21]
  wire  MAT_io_hit; // @[processor_pisa.scala 19:21]
  wire [63:0] MAT_io_match_value; // @[processor_pisa.scala 19:21]
  wire  EXE_clock; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_0; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_1; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_2; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_3; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_4; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_5; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_6; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_7; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_8; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_9; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_10; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_11; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_12; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_13; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_14; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_15; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_16; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_17; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_18; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_19; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_20; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_21; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_22; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_23; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_24; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_25; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_26; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_27; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_28; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_29; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_30; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_31; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_32; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_33; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_34; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_35; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_36; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_37; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_38; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_39; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_40; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_41; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_42; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_43; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_44; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_45; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_46; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_47; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_48; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_49; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_50; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_51; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_52; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_53; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_54; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_55; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_56; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_57; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_58; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_59; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_60; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_61; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_62; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_63; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_64; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_65; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_66; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_67; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_68; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_69; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_70; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_71; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_72; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_73; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_74; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_75; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_76; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_77; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_78; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_79; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_80; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_81; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_82; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_83; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_84; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_85; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_86; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_87; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_88; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_89; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_90; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_91; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_92; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_93; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_94; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_95; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_96; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_97; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_98; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_99; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_100; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_101; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_102; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_103; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_104; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_105; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_106; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_107; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_108; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_109; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_110; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_111; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_112; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_113; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_114; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_115; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_116; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_117; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_118; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_119; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_120; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_121; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_122; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_123; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_124; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_125; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_126; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_127; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_128; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_129; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_130; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_131; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_132; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_133; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_134; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_135; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_136; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_137; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_138; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_139; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_140; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_141; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_142; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_143; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_144; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_145; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_146; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_147; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_148; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_149; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_150; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_151; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_152; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_153; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_154; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_155; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_156; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_157; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_158; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_159; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_160; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_161; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_162; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_163; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_164; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_165; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_166; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_167; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_168; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_169; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_170; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_171; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_172; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_173; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_174; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_175; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_176; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_177; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_178; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_179; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_180; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_181; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_182; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_183; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_184; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_185; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_186; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_187; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_188; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_189; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_190; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_191; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_192; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_193; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_194; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_195; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_196; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_197; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_198; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_199; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_200; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_201; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_202; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_203; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_204; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_205; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_206; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_207; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_208; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_209; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_210; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_211; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_212; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_213; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_214; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_215; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_216; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_217; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_218; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_219; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_220; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_221; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_222; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_223; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_224; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_225; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_226; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_227; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_228; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_229; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_230; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_231; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_232; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_233; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_234; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_235; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_236; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_237; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_238; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_239; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_240; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_241; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_242; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_243; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_244; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_245; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_246; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_247; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_248; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_249; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_250; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_251; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_252; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_253; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_254; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_in_data_255; // @[processor_pisa.scala 20:21]
  wire [3:0] EXE_io_pipe_phv_in_next_processor_id; // @[processor_pisa.scala 20:21]
  wire  EXE_io_pipe_phv_in_next_config_id; // @[processor_pisa.scala 20:21]
  wire  EXE_io_pipe_phv_in_is_valid_processor; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_0; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_1; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_2; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_3; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_4; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_5; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_6; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_7; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_8; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_9; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_10; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_11; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_12; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_13; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_14; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_15; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_16; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_17; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_18; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_19; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_20; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_21; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_22; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_23; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_24; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_25; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_26; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_27; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_28; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_29; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_30; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_31; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_32; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_33; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_34; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_35; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_36; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_37; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_38; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_39; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_40; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_41; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_42; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_43; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_44; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_45; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_46; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_47; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_48; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_49; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_50; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_51; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_52; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_53; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_54; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_55; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_56; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_57; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_58; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_59; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_60; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_61; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_62; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_63; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_64; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_65; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_66; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_67; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_68; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_69; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_70; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_71; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_72; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_73; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_74; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_75; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_76; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_77; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_78; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_79; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_80; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_81; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_82; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_83; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_84; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_85; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_86; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_87; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_88; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_89; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_90; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_91; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_92; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_93; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_94; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_95; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_96; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_97; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_98; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_99; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_100; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_101; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_102; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_103; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_104; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_105; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_106; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_107; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_108; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_109; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_110; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_111; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_112; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_113; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_114; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_115; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_116; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_117; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_118; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_119; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_120; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_121; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_122; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_123; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_124; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_125; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_126; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_127; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_128; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_129; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_130; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_131; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_132; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_133; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_134; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_135; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_136; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_137; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_138; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_139; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_140; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_141; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_142; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_143; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_144; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_145; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_146; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_147; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_148; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_149; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_150; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_151; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_152; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_153; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_154; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_155; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_156; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_157; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_158; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_159; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_160; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_161; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_162; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_163; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_164; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_165; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_166; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_167; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_168; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_169; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_170; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_171; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_172; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_173; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_174; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_175; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_176; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_177; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_178; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_179; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_180; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_181; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_182; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_183; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_184; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_185; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_186; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_187; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_188; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_189; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_190; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_191; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_192; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_193; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_194; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_195; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_196; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_197; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_198; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_199; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_200; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_201; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_202; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_203; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_204; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_205; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_206; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_207; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_208; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_209; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_210; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_211; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_212; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_213; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_214; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_215; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_216; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_217; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_218; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_219; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_220; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_221; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_222; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_223; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_224; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_225; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_226; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_227; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_228; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_229; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_230; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_231; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_232; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_233; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_234; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_235; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_236; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_237; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_238; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_239; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_240; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_241; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_242; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_243; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_244; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_245; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_246; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_247; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_248; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_249; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_250; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_251; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_252; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_253; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_254; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_pipe_phv_out_data_255; // @[processor_pisa.scala 20:21]
  wire [3:0] EXE_io_pipe_phv_out_next_processor_id; // @[processor_pisa.scala 20:21]
  wire  EXE_io_pipe_phv_out_next_config_id; // @[processor_pisa.scala 20:21]
  wire  EXE_io_hit; // @[processor_pisa.scala 20:21]
  wire [63:0] EXE_io_match_value; // @[processor_pisa.scala 20:21]
  wire  EXE_io_action_mod_en_0; // @[processor_pisa.scala 20:21]
  wire  EXE_io_action_mod_en_1; // @[processor_pisa.scala 20:21]
  wire [7:0] EXE_io_action_mod_addr; // @[processor_pisa.scala 20:21]
  wire [63:0] EXE_io_action_mod_data_0; // @[processor_pisa.scala 20:21]
  wire [63:0] EXE_io_action_mod_data_1; // @[processor_pisa.scala 20:21]
  MatcherPISA MAT ( // @[processor_pisa.scala 19:21]
    .clock(MAT_clock),
    .io_pipe_phv_in_data_0(MAT_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(MAT_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(MAT_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(MAT_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(MAT_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(MAT_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(MAT_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(MAT_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(MAT_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(MAT_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(MAT_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(MAT_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(MAT_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(MAT_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(MAT_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(MAT_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(MAT_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(MAT_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(MAT_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(MAT_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(MAT_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(MAT_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(MAT_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(MAT_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(MAT_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(MAT_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(MAT_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(MAT_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(MAT_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(MAT_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(MAT_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(MAT_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(MAT_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(MAT_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(MAT_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(MAT_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(MAT_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(MAT_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(MAT_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(MAT_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(MAT_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(MAT_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(MAT_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(MAT_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(MAT_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(MAT_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(MAT_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(MAT_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(MAT_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(MAT_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(MAT_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(MAT_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(MAT_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(MAT_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(MAT_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(MAT_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(MAT_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(MAT_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(MAT_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(MAT_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(MAT_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(MAT_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(MAT_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(MAT_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(MAT_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(MAT_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(MAT_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(MAT_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(MAT_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(MAT_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(MAT_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(MAT_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(MAT_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(MAT_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(MAT_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(MAT_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(MAT_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(MAT_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(MAT_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(MAT_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(MAT_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(MAT_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(MAT_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(MAT_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(MAT_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(MAT_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(MAT_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(MAT_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(MAT_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(MAT_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(MAT_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(MAT_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(MAT_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(MAT_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(MAT_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(MAT_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(MAT_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(MAT_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(MAT_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(MAT_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(MAT_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(MAT_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(MAT_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(MAT_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(MAT_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(MAT_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(MAT_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(MAT_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(MAT_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(MAT_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(MAT_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(MAT_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(MAT_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(MAT_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(MAT_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(MAT_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(MAT_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(MAT_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(MAT_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(MAT_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(MAT_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(MAT_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(MAT_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(MAT_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(MAT_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(MAT_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(MAT_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(MAT_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(MAT_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(MAT_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(MAT_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(MAT_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(MAT_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(MAT_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(MAT_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(MAT_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(MAT_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(MAT_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(MAT_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(MAT_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(MAT_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(MAT_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(MAT_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(MAT_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(MAT_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(MAT_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(MAT_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(MAT_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(MAT_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(MAT_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(MAT_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(MAT_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(MAT_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(MAT_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(MAT_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(MAT_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(MAT_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(MAT_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(MAT_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(MAT_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(MAT_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(MAT_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(MAT_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(MAT_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(MAT_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(MAT_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(MAT_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(MAT_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(MAT_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(MAT_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(MAT_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(MAT_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(MAT_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(MAT_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(MAT_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(MAT_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(MAT_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(MAT_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(MAT_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(MAT_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(MAT_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(MAT_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(MAT_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(MAT_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(MAT_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(MAT_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(MAT_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(MAT_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(MAT_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(MAT_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(MAT_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(MAT_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(MAT_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(MAT_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(MAT_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(MAT_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(MAT_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(MAT_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(MAT_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(MAT_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(MAT_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(MAT_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(MAT_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(MAT_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(MAT_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(MAT_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(MAT_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(MAT_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(MAT_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(MAT_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(MAT_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(MAT_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(MAT_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(MAT_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(MAT_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(MAT_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(MAT_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(MAT_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(MAT_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(MAT_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(MAT_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(MAT_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(MAT_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(MAT_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(MAT_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(MAT_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(MAT_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(MAT_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(MAT_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(MAT_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(MAT_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(MAT_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(MAT_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(MAT_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(MAT_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(MAT_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(MAT_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(MAT_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(MAT_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(MAT_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(MAT_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(MAT_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(MAT_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(MAT_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(MAT_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(MAT_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(MAT_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(MAT_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(MAT_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(MAT_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(MAT_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(MAT_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(MAT_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(MAT_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(MAT_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(MAT_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_next_processor_id(MAT_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(MAT_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(MAT_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(MAT_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(MAT_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(MAT_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(MAT_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(MAT_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(MAT_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(MAT_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(MAT_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(MAT_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(MAT_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(MAT_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(MAT_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(MAT_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(MAT_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(MAT_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(MAT_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(MAT_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(MAT_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(MAT_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(MAT_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(MAT_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(MAT_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(MAT_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(MAT_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(MAT_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(MAT_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(MAT_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(MAT_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(MAT_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(MAT_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(MAT_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(MAT_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(MAT_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(MAT_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(MAT_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(MAT_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(MAT_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(MAT_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(MAT_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(MAT_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(MAT_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(MAT_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(MAT_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(MAT_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(MAT_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(MAT_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(MAT_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(MAT_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(MAT_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(MAT_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(MAT_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(MAT_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(MAT_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(MAT_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(MAT_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(MAT_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(MAT_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(MAT_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(MAT_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(MAT_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(MAT_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(MAT_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(MAT_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(MAT_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(MAT_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(MAT_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(MAT_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(MAT_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(MAT_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(MAT_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(MAT_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(MAT_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(MAT_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(MAT_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(MAT_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(MAT_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(MAT_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(MAT_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(MAT_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(MAT_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(MAT_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(MAT_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(MAT_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(MAT_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(MAT_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(MAT_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(MAT_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(MAT_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(MAT_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(MAT_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(MAT_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(MAT_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(MAT_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(MAT_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(MAT_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(MAT_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(MAT_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(MAT_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(MAT_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(MAT_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(MAT_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(MAT_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(MAT_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(MAT_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(MAT_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(MAT_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(MAT_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(MAT_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(MAT_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(MAT_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(MAT_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(MAT_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(MAT_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(MAT_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(MAT_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(MAT_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(MAT_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(MAT_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(MAT_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(MAT_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(MAT_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(MAT_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(MAT_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(MAT_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(MAT_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(MAT_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(MAT_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(MAT_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(MAT_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(MAT_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(MAT_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(MAT_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(MAT_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(MAT_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(MAT_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(MAT_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(MAT_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(MAT_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(MAT_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(MAT_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(MAT_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(MAT_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(MAT_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(MAT_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(MAT_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(MAT_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(MAT_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(MAT_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(MAT_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(MAT_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(MAT_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(MAT_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(MAT_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(MAT_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(MAT_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(MAT_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(MAT_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(MAT_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(MAT_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(MAT_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(MAT_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(MAT_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(MAT_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(MAT_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(MAT_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(MAT_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(MAT_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(MAT_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(MAT_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(MAT_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(MAT_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(MAT_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(MAT_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(MAT_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(MAT_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(MAT_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(MAT_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(MAT_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(MAT_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(MAT_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(MAT_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(MAT_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(MAT_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(MAT_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(MAT_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(MAT_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(MAT_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(MAT_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(MAT_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(MAT_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(MAT_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(MAT_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(MAT_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(MAT_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(MAT_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(MAT_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(MAT_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(MAT_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(MAT_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(MAT_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(MAT_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(MAT_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(MAT_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(MAT_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(MAT_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(MAT_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(MAT_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(MAT_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(MAT_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(MAT_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(MAT_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(MAT_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(MAT_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(MAT_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(MAT_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(MAT_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(MAT_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(MAT_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(MAT_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(MAT_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(MAT_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(MAT_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(MAT_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(MAT_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(MAT_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(MAT_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(MAT_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(MAT_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(MAT_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(MAT_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(MAT_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(MAT_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(MAT_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(MAT_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(MAT_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(MAT_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(MAT_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(MAT_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(MAT_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(MAT_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(MAT_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(MAT_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(MAT_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(MAT_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(MAT_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(MAT_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(MAT_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(MAT_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(MAT_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(MAT_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(MAT_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(MAT_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(MAT_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(MAT_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(MAT_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(MAT_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_next_processor_id(MAT_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(MAT_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(MAT_io_pipe_phv_out_is_valid_processor),
    .io_mod_en(MAT_io_mod_en),
    .io_mod_config_id(MAT_io_mod_config_id),
    .io_mod_key_mod_en(MAT_io_mod_key_mod_en),
    .io_mod_key_mod_group_index(MAT_io_mod_key_mod_group_index),
    .io_mod_key_mod_group_config(MAT_io_mod_key_mod_group_config),
    .io_mod_key_mod_group_mask_0(MAT_io_mod_key_mod_group_mask_0),
    .io_mod_key_mod_group_mask_1(MAT_io_mod_key_mod_group_mask_1),
    .io_mod_key_mod_group_mask_2(MAT_io_mod_key_mod_group_mask_2),
    .io_mod_key_mod_group_mask_3(MAT_io_mod_key_mod_group_mask_3),
    .io_mod_key_mod_group_id_0(MAT_io_mod_key_mod_group_id_0),
    .io_mod_key_mod_group_id_1(MAT_io_mod_key_mod_group_id_1),
    .io_mod_key_mod_group_id_2(MAT_io_mod_key_mod_group_id_2),
    .io_mod_key_mod_group_id_3(MAT_io_mod_key_mod_group_id_3),
    .io_mod_table_mod_table_depth(MAT_io_mod_table_mod_table_depth),
    .io_mod_table_mod_table_width(MAT_io_mod_table_mod_table_width),
    .io_mod_w_en(MAT_io_mod_w_en),
    .io_mod_w_sram_id(MAT_io_mod_w_sram_id),
    .io_mod_w_addr(MAT_io_mod_w_addr),
    .io_mod_w_data(MAT_io_mod_w_data),
    .io_hit(MAT_io_hit),
    .io_match_value(MAT_io_match_value)
  );
  ExecutorPISA EXE ( // @[processor_pisa.scala 20:21]
    .clock(EXE_clock),
    .io_pipe_phv_in_data_0(EXE_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(EXE_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(EXE_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(EXE_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(EXE_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(EXE_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(EXE_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(EXE_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(EXE_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(EXE_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(EXE_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(EXE_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(EXE_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(EXE_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(EXE_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(EXE_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(EXE_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(EXE_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(EXE_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(EXE_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(EXE_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(EXE_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(EXE_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(EXE_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(EXE_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(EXE_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(EXE_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(EXE_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(EXE_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(EXE_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(EXE_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(EXE_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(EXE_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(EXE_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(EXE_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(EXE_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(EXE_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(EXE_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(EXE_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(EXE_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(EXE_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(EXE_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(EXE_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(EXE_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(EXE_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(EXE_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(EXE_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(EXE_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(EXE_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(EXE_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(EXE_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(EXE_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(EXE_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(EXE_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(EXE_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(EXE_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(EXE_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(EXE_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(EXE_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(EXE_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(EXE_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(EXE_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(EXE_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(EXE_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(EXE_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(EXE_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(EXE_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(EXE_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(EXE_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(EXE_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(EXE_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(EXE_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(EXE_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(EXE_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(EXE_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(EXE_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(EXE_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(EXE_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(EXE_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(EXE_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(EXE_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(EXE_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(EXE_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(EXE_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(EXE_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(EXE_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(EXE_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(EXE_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(EXE_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(EXE_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(EXE_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(EXE_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(EXE_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(EXE_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(EXE_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(EXE_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(EXE_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(EXE_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(EXE_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(EXE_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(EXE_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(EXE_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(EXE_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(EXE_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(EXE_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(EXE_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(EXE_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(EXE_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(EXE_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(EXE_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(EXE_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(EXE_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(EXE_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(EXE_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(EXE_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(EXE_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(EXE_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(EXE_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(EXE_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(EXE_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(EXE_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(EXE_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(EXE_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(EXE_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(EXE_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(EXE_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(EXE_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(EXE_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(EXE_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(EXE_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(EXE_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(EXE_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(EXE_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(EXE_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(EXE_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(EXE_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(EXE_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(EXE_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(EXE_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(EXE_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(EXE_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(EXE_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(EXE_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(EXE_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(EXE_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(EXE_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(EXE_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(EXE_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(EXE_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(EXE_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(EXE_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(EXE_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(EXE_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(EXE_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(EXE_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(EXE_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(EXE_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(EXE_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(EXE_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(EXE_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(EXE_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(EXE_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(EXE_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(EXE_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(EXE_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(EXE_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(EXE_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(EXE_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(EXE_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(EXE_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(EXE_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(EXE_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(EXE_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(EXE_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(EXE_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(EXE_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(EXE_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(EXE_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(EXE_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(EXE_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(EXE_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(EXE_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(EXE_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(EXE_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(EXE_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(EXE_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(EXE_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(EXE_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(EXE_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(EXE_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(EXE_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(EXE_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(EXE_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(EXE_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(EXE_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(EXE_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(EXE_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(EXE_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(EXE_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(EXE_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(EXE_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(EXE_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(EXE_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(EXE_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(EXE_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(EXE_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(EXE_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(EXE_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(EXE_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(EXE_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(EXE_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(EXE_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(EXE_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(EXE_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(EXE_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(EXE_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(EXE_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(EXE_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(EXE_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(EXE_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(EXE_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(EXE_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(EXE_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(EXE_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(EXE_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(EXE_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(EXE_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(EXE_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(EXE_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(EXE_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(EXE_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(EXE_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(EXE_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(EXE_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(EXE_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(EXE_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(EXE_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(EXE_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(EXE_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(EXE_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(EXE_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(EXE_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(EXE_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(EXE_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(EXE_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(EXE_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(EXE_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(EXE_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(EXE_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(EXE_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(EXE_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(EXE_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(EXE_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(EXE_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(EXE_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(EXE_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_next_processor_id(EXE_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(EXE_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(EXE_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(EXE_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(EXE_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(EXE_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(EXE_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(EXE_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(EXE_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(EXE_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(EXE_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(EXE_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(EXE_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(EXE_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(EXE_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(EXE_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(EXE_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(EXE_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(EXE_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(EXE_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(EXE_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(EXE_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(EXE_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(EXE_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(EXE_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(EXE_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(EXE_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(EXE_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(EXE_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(EXE_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(EXE_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(EXE_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(EXE_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(EXE_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(EXE_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(EXE_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(EXE_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(EXE_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(EXE_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(EXE_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(EXE_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(EXE_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(EXE_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(EXE_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(EXE_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(EXE_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(EXE_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(EXE_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(EXE_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(EXE_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(EXE_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(EXE_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(EXE_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(EXE_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(EXE_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(EXE_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(EXE_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(EXE_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(EXE_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(EXE_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(EXE_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(EXE_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(EXE_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(EXE_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(EXE_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(EXE_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(EXE_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(EXE_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(EXE_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(EXE_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(EXE_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(EXE_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(EXE_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(EXE_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(EXE_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(EXE_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(EXE_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(EXE_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(EXE_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(EXE_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(EXE_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(EXE_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(EXE_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(EXE_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(EXE_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(EXE_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(EXE_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(EXE_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(EXE_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(EXE_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(EXE_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(EXE_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(EXE_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(EXE_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(EXE_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(EXE_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(EXE_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(EXE_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(EXE_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(EXE_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(EXE_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(EXE_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(EXE_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(EXE_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(EXE_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(EXE_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(EXE_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(EXE_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(EXE_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(EXE_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(EXE_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(EXE_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(EXE_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(EXE_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(EXE_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(EXE_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(EXE_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(EXE_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(EXE_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(EXE_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(EXE_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(EXE_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(EXE_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(EXE_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(EXE_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(EXE_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(EXE_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(EXE_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(EXE_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(EXE_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(EXE_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(EXE_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(EXE_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(EXE_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(EXE_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(EXE_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(EXE_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(EXE_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(EXE_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(EXE_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(EXE_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(EXE_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(EXE_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(EXE_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(EXE_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(EXE_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(EXE_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(EXE_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(EXE_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(EXE_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(EXE_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(EXE_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(EXE_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(EXE_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(EXE_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(EXE_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(EXE_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(EXE_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(EXE_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(EXE_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(EXE_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(EXE_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(EXE_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(EXE_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(EXE_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(EXE_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(EXE_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(EXE_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(EXE_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(EXE_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(EXE_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(EXE_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(EXE_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(EXE_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(EXE_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(EXE_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(EXE_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(EXE_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(EXE_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(EXE_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(EXE_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(EXE_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(EXE_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(EXE_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(EXE_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(EXE_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(EXE_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(EXE_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(EXE_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(EXE_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(EXE_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(EXE_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(EXE_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(EXE_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(EXE_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(EXE_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(EXE_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(EXE_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(EXE_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(EXE_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(EXE_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(EXE_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(EXE_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(EXE_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(EXE_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(EXE_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(EXE_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(EXE_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(EXE_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(EXE_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(EXE_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(EXE_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(EXE_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(EXE_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(EXE_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(EXE_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(EXE_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(EXE_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(EXE_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(EXE_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(EXE_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(EXE_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(EXE_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(EXE_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(EXE_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(EXE_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(EXE_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(EXE_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(EXE_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(EXE_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(EXE_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(EXE_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(EXE_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(EXE_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(EXE_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(EXE_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(EXE_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(EXE_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(EXE_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(EXE_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(EXE_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(EXE_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(EXE_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(EXE_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(EXE_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(EXE_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(EXE_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(EXE_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(EXE_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(EXE_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(EXE_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(EXE_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(EXE_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(EXE_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(EXE_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(EXE_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(EXE_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(EXE_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(EXE_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_next_processor_id(EXE_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(EXE_io_pipe_phv_out_next_config_id),
    .io_hit(EXE_io_hit),
    .io_match_value(EXE_io_match_value),
    .io_action_mod_en_0(EXE_io_action_mod_en_0),
    .io_action_mod_en_1(EXE_io_action_mod_en_1),
    .io_action_mod_addr(EXE_io_action_mod_addr),
    .io_action_mod_data_0(EXE_io_action_mod_data_0),
    .io_action_mod_data_1(EXE_io_action_mod_data_1)
  );
  assign io_pipe_phv_out_data_0 = EXE_io_pipe_phv_out_data_0; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_1 = EXE_io_pipe_phv_out_data_1; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_2 = EXE_io_pipe_phv_out_data_2; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_3 = EXE_io_pipe_phv_out_data_3; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_4 = EXE_io_pipe_phv_out_data_4; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_5 = EXE_io_pipe_phv_out_data_5; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_6 = EXE_io_pipe_phv_out_data_6; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_7 = EXE_io_pipe_phv_out_data_7; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_8 = EXE_io_pipe_phv_out_data_8; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_9 = EXE_io_pipe_phv_out_data_9; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_10 = EXE_io_pipe_phv_out_data_10; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_11 = EXE_io_pipe_phv_out_data_11; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_12 = EXE_io_pipe_phv_out_data_12; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_13 = EXE_io_pipe_phv_out_data_13; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_14 = EXE_io_pipe_phv_out_data_14; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_15 = EXE_io_pipe_phv_out_data_15; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_16 = EXE_io_pipe_phv_out_data_16; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_17 = EXE_io_pipe_phv_out_data_17; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_18 = EXE_io_pipe_phv_out_data_18; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_19 = EXE_io_pipe_phv_out_data_19; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_20 = EXE_io_pipe_phv_out_data_20; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_21 = EXE_io_pipe_phv_out_data_21; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_22 = EXE_io_pipe_phv_out_data_22; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_23 = EXE_io_pipe_phv_out_data_23; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_24 = EXE_io_pipe_phv_out_data_24; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_25 = EXE_io_pipe_phv_out_data_25; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_26 = EXE_io_pipe_phv_out_data_26; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_27 = EXE_io_pipe_phv_out_data_27; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_28 = EXE_io_pipe_phv_out_data_28; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_29 = EXE_io_pipe_phv_out_data_29; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_30 = EXE_io_pipe_phv_out_data_30; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_31 = EXE_io_pipe_phv_out_data_31; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_32 = EXE_io_pipe_phv_out_data_32; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_33 = EXE_io_pipe_phv_out_data_33; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_34 = EXE_io_pipe_phv_out_data_34; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_35 = EXE_io_pipe_phv_out_data_35; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_36 = EXE_io_pipe_phv_out_data_36; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_37 = EXE_io_pipe_phv_out_data_37; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_38 = EXE_io_pipe_phv_out_data_38; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_39 = EXE_io_pipe_phv_out_data_39; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_40 = EXE_io_pipe_phv_out_data_40; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_41 = EXE_io_pipe_phv_out_data_41; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_42 = EXE_io_pipe_phv_out_data_42; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_43 = EXE_io_pipe_phv_out_data_43; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_44 = EXE_io_pipe_phv_out_data_44; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_45 = EXE_io_pipe_phv_out_data_45; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_46 = EXE_io_pipe_phv_out_data_46; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_47 = EXE_io_pipe_phv_out_data_47; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_48 = EXE_io_pipe_phv_out_data_48; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_49 = EXE_io_pipe_phv_out_data_49; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_50 = EXE_io_pipe_phv_out_data_50; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_51 = EXE_io_pipe_phv_out_data_51; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_52 = EXE_io_pipe_phv_out_data_52; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_53 = EXE_io_pipe_phv_out_data_53; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_54 = EXE_io_pipe_phv_out_data_54; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_55 = EXE_io_pipe_phv_out_data_55; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_56 = EXE_io_pipe_phv_out_data_56; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_57 = EXE_io_pipe_phv_out_data_57; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_58 = EXE_io_pipe_phv_out_data_58; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_59 = EXE_io_pipe_phv_out_data_59; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_60 = EXE_io_pipe_phv_out_data_60; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_61 = EXE_io_pipe_phv_out_data_61; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_62 = EXE_io_pipe_phv_out_data_62; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_63 = EXE_io_pipe_phv_out_data_63; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_64 = EXE_io_pipe_phv_out_data_64; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_65 = EXE_io_pipe_phv_out_data_65; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_66 = EXE_io_pipe_phv_out_data_66; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_67 = EXE_io_pipe_phv_out_data_67; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_68 = EXE_io_pipe_phv_out_data_68; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_69 = EXE_io_pipe_phv_out_data_69; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_70 = EXE_io_pipe_phv_out_data_70; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_71 = EXE_io_pipe_phv_out_data_71; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_72 = EXE_io_pipe_phv_out_data_72; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_73 = EXE_io_pipe_phv_out_data_73; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_74 = EXE_io_pipe_phv_out_data_74; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_75 = EXE_io_pipe_phv_out_data_75; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_76 = EXE_io_pipe_phv_out_data_76; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_77 = EXE_io_pipe_phv_out_data_77; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_78 = EXE_io_pipe_phv_out_data_78; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_79 = EXE_io_pipe_phv_out_data_79; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_80 = EXE_io_pipe_phv_out_data_80; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_81 = EXE_io_pipe_phv_out_data_81; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_82 = EXE_io_pipe_phv_out_data_82; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_83 = EXE_io_pipe_phv_out_data_83; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_84 = EXE_io_pipe_phv_out_data_84; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_85 = EXE_io_pipe_phv_out_data_85; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_86 = EXE_io_pipe_phv_out_data_86; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_87 = EXE_io_pipe_phv_out_data_87; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_88 = EXE_io_pipe_phv_out_data_88; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_89 = EXE_io_pipe_phv_out_data_89; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_90 = EXE_io_pipe_phv_out_data_90; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_91 = EXE_io_pipe_phv_out_data_91; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_92 = EXE_io_pipe_phv_out_data_92; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_93 = EXE_io_pipe_phv_out_data_93; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_94 = EXE_io_pipe_phv_out_data_94; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_95 = EXE_io_pipe_phv_out_data_95; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_96 = EXE_io_pipe_phv_out_data_96; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_97 = EXE_io_pipe_phv_out_data_97; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_98 = EXE_io_pipe_phv_out_data_98; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_99 = EXE_io_pipe_phv_out_data_99; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_100 = EXE_io_pipe_phv_out_data_100; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_101 = EXE_io_pipe_phv_out_data_101; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_102 = EXE_io_pipe_phv_out_data_102; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_103 = EXE_io_pipe_phv_out_data_103; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_104 = EXE_io_pipe_phv_out_data_104; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_105 = EXE_io_pipe_phv_out_data_105; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_106 = EXE_io_pipe_phv_out_data_106; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_107 = EXE_io_pipe_phv_out_data_107; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_108 = EXE_io_pipe_phv_out_data_108; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_109 = EXE_io_pipe_phv_out_data_109; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_110 = EXE_io_pipe_phv_out_data_110; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_111 = EXE_io_pipe_phv_out_data_111; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_112 = EXE_io_pipe_phv_out_data_112; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_113 = EXE_io_pipe_phv_out_data_113; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_114 = EXE_io_pipe_phv_out_data_114; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_115 = EXE_io_pipe_phv_out_data_115; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_116 = EXE_io_pipe_phv_out_data_116; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_117 = EXE_io_pipe_phv_out_data_117; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_118 = EXE_io_pipe_phv_out_data_118; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_119 = EXE_io_pipe_phv_out_data_119; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_120 = EXE_io_pipe_phv_out_data_120; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_121 = EXE_io_pipe_phv_out_data_121; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_122 = EXE_io_pipe_phv_out_data_122; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_123 = EXE_io_pipe_phv_out_data_123; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_124 = EXE_io_pipe_phv_out_data_124; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_125 = EXE_io_pipe_phv_out_data_125; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_126 = EXE_io_pipe_phv_out_data_126; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_127 = EXE_io_pipe_phv_out_data_127; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_128 = EXE_io_pipe_phv_out_data_128; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_129 = EXE_io_pipe_phv_out_data_129; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_130 = EXE_io_pipe_phv_out_data_130; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_131 = EXE_io_pipe_phv_out_data_131; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_132 = EXE_io_pipe_phv_out_data_132; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_133 = EXE_io_pipe_phv_out_data_133; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_134 = EXE_io_pipe_phv_out_data_134; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_135 = EXE_io_pipe_phv_out_data_135; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_136 = EXE_io_pipe_phv_out_data_136; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_137 = EXE_io_pipe_phv_out_data_137; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_138 = EXE_io_pipe_phv_out_data_138; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_139 = EXE_io_pipe_phv_out_data_139; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_140 = EXE_io_pipe_phv_out_data_140; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_141 = EXE_io_pipe_phv_out_data_141; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_142 = EXE_io_pipe_phv_out_data_142; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_143 = EXE_io_pipe_phv_out_data_143; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_144 = EXE_io_pipe_phv_out_data_144; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_145 = EXE_io_pipe_phv_out_data_145; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_146 = EXE_io_pipe_phv_out_data_146; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_147 = EXE_io_pipe_phv_out_data_147; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_148 = EXE_io_pipe_phv_out_data_148; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_149 = EXE_io_pipe_phv_out_data_149; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_150 = EXE_io_pipe_phv_out_data_150; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_151 = EXE_io_pipe_phv_out_data_151; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_152 = EXE_io_pipe_phv_out_data_152; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_153 = EXE_io_pipe_phv_out_data_153; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_154 = EXE_io_pipe_phv_out_data_154; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_155 = EXE_io_pipe_phv_out_data_155; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_156 = EXE_io_pipe_phv_out_data_156; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_157 = EXE_io_pipe_phv_out_data_157; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_158 = EXE_io_pipe_phv_out_data_158; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_159 = EXE_io_pipe_phv_out_data_159; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_160 = EXE_io_pipe_phv_out_data_160; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_161 = EXE_io_pipe_phv_out_data_161; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_162 = EXE_io_pipe_phv_out_data_162; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_163 = EXE_io_pipe_phv_out_data_163; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_164 = EXE_io_pipe_phv_out_data_164; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_165 = EXE_io_pipe_phv_out_data_165; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_166 = EXE_io_pipe_phv_out_data_166; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_167 = EXE_io_pipe_phv_out_data_167; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_168 = EXE_io_pipe_phv_out_data_168; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_169 = EXE_io_pipe_phv_out_data_169; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_170 = EXE_io_pipe_phv_out_data_170; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_171 = EXE_io_pipe_phv_out_data_171; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_172 = EXE_io_pipe_phv_out_data_172; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_173 = EXE_io_pipe_phv_out_data_173; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_174 = EXE_io_pipe_phv_out_data_174; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_175 = EXE_io_pipe_phv_out_data_175; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_176 = EXE_io_pipe_phv_out_data_176; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_177 = EXE_io_pipe_phv_out_data_177; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_178 = EXE_io_pipe_phv_out_data_178; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_179 = EXE_io_pipe_phv_out_data_179; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_180 = EXE_io_pipe_phv_out_data_180; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_181 = EXE_io_pipe_phv_out_data_181; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_182 = EXE_io_pipe_phv_out_data_182; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_183 = EXE_io_pipe_phv_out_data_183; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_184 = EXE_io_pipe_phv_out_data_184; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_185 = EXE_io_pipe_phv_out_data_185; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_186 = EXE_io_pipe_phv_out_data_186; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_187 = EXE_io_pipe_phv_out_data_187; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_188 = EXE_io_pipe_phv_out_data_188; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_189 = EXE_io_pipe_phv_out_data_189; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_190 = EXE_io_pipe_phv_out_data_190; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_191 = EXE_io_pipe_phv_out_data_191; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_192 = EXE_io_pipe_phv_out_data_192; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_193 = EXE_io_pipe_phv_out_data_193; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_194 = EXE_io_pipe_phv_out_data_194; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_195 = EXE_io_pipe_phv_out_data_195; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_196 = EXE_io_pipe_phv_out_data_196; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_197 = EXE_io_pipe_phv_out_data_197; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_198 = EXE_io_pipe_phv_out_data_198; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_199 = EXE_io_pipe_phv_out_data_199; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_200 = EXE_io_pipe_phv_out_data_200; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_201 = EXE_io_pipe_phv_out_data_201; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_202 = EXE_io_pipe_phv_out_data_202; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_203 = EXE_io_pipe_phv_out_data_203; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_204 = EXE_io_pipe_phv_out_data_204; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_205 = EXE_io_pipe_phv_out_data_205; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_206 = EXE_io_pipe_phv_out_data_206; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_207 = EXE_io_pipe_phv_out_data_207; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_208 = EXE_io_pipe_phv_out_data_208; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_209 = EXE_io_pipe_phv_out_data_209; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_210 = EXE_io_pipe_phv_out_data_210; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_211 = EXE_io_pipe_phv_out_data_211; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_212 = EXE_io_pipe_phv_out_data_212; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_213 = EXE_io_pipe_phv_out_data_213; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_214 = EXE_io_pipe_phv_out_data_214; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_215 = EXE_io_pipe_phv_out_data_215; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_216 = EXE_io_pipe_phv_out_data_216; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_217 = EXE_io_pipe_phv_out_data_217; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_218 = EXE_io_pipe_phv_out_data_218; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_219 = EXE_io_pipe_phv_out_data_219; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_220 = EXE_io_pipe_phv_out_data_220; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_221 = EXE_io_pipe_phv_out_data_221; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_222 = EXE_io_pipe_phv_out_data_222; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_223 = EXE_io_pipe_phv_out_data_223; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_224 = EXE_io_pipe_phv_out_data_224; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_225 = EXE_io_pipe_phv_out_data_225; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_226 = EXE_io_pipe_phv_out_data_226; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_227 = EXE_io_pipe_phv_out_data_227; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_228 = EXE_io_pipe_phv_out_data_228; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_229 = EXE_io_pipe_phv_out_data_229; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_230 = EXE_io_pipe_phv_out_data_230; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_231 = EXE_io_pipe_phv_out_data_231; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_232 = EXE_io_pipe_phv_out_data_232; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_233 = EXE_io_pipe_phv_out_data_233; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_234 = EXE_io_pipe_phv_out_data_234; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_235 = EXE_io_pipe_phv_out_data_235; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_236 = EXE_io_pipe_phv_out_data_236; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_237 = EXE_io_pipe_phv_out_data_237; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_238 = EXE_io_pipe_phv_out_data_238; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_239 = EXE_io_pipe_phv_out_data_239; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_240 = EXE_io_pipe_phv_out_data_240; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_241 = EXE_io_pipe_phv_out_data_241; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_242 = EXE_io_pipe_phv_out_data_242; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_243 = EXE_io_pipe_phv_out_data_243; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_244 = EXE_io_pipe_phv_out_data_244; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_245 = EXE_io_pipe_phv_out_data_245; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_246 = EXE_io_pipe_phv_out_data_246; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_247 = EXE_io_pipe_phv_out_data_247; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_248 = EXE_io_pipe_phv_out_data_248; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_249 = EXE_io_pipe_phv_out_data_249; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_250 = EXE_io_pipe_phv_out_data_250; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_251 = EXE_io_pipe_phv_out_data_251; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_252 = EXE_io_pipe_phv_out_data_252; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_253 = EXE_io_pipe_phv_out_data_253; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_254 = EXE_io_pipe_phv_out_data_254; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_data_255 = EXE_io_pipe_phv_out_data_255; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_next_processor_id = EXE_io_pipe_phv_out_next_processor_id; // @[processor_pisa.scala 33:24]
  assign io_pipe_phv_out_next_config_id = EXE_io_pipe_phv_out_next_config_id; // @[processor_pisa.scala 33:24]
  assign MAT_clock = clock;
  assign MAT_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_96 = io_pipe_phv_in_data_96; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_97 = io_pipe_phv_in_data_97; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_98 = io_pipe_phv_in_data_98; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_99 = io_pipe_phv_in_data_99; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_100 = io_pipe_phv_in_data_100; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_101 = io_pipe_phv_in_data_101; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_102 = io_pipe_phv_in_data_102; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_103 = io_pipe_phv_in_data_103; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_104 = io_pipe_phv_in_data_104; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_105 = io_pipe_phv_in_data_105; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_106 = io_pipe_phv_in_data_106; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_107 = io_pipe_phv_in_data_107; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_108 = io_pipe_phv_in_data_108; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_109 = io_pipe_phv_in_data_109; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_110 = io_pipe_phv_in_data_110; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_111 = io_pipe_phv_in_data_111; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_112 = io_pipe_phv_in_data_112; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_113 = io_pipe_phv_in_data_113; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_114 = io_pipe_phv_in_data_114; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_115 = io_pipe_phv_in_data_115; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_116 = io_pipe_phv_in_data_116; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_117 = io_pipe_phv_in_data_117; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_118 = io_pipe_phv_in_data_118; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_119 = io_pipe_phv_in_data_119; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_120 = io_pipe_phv_in_data_120; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_121 = io_pipe_phv_in_data_121; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_122 = io_pipe_phv_in_data_122; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_123 = io_pipe_phv_in_data_123; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_124 = io_pipe_phv_in_data_124; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_125 = io_pipe_phv_in_data_125; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_126 = io_pipe_phv_in_data_126; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_127 = io_pipe_phv_in_data_127; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_128 = io_pipe_phv_in_data_128; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_129 = io_pipe_phv_in_data_129; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_130 = io_pipe_phv_in_data_130; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_131 = io_pipe_phv_in_data_131; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_132 = io_pipe_phv_in_data_132; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_133 = io_pipe_phv_in_data_133; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_134 = io_pipe_phv_in_data_134; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_135 = io_pipe_phv_in_data_135; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_136 = io_pipe_phv_in_data_136; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_137 = io_pipe_phv_in_data_137; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_138 = io_pipe_phv_in_data_138; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_139 = io_pipe_phv_in_data_139; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_140 = io_pipe_phv_in_data_140; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_141 = io_pipe_phv_in_data_141; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_142 = io_pipe_phv_in_data_142; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_143 = io_pipe_phv_in_data_143; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_144 = io_pipe_phv_in_data_144; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_145 = io_pipe_phv_in_data_145; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_146 = io_pipe_phv_in_data_146; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_147 = io_pipe_phv_in_data_147; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_148 = io_pipe_phv_in_data_148; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_149 = io_pipe_phv_in_data_149; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_150 = io_pipe_phv_in_data_150; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_151 = io_pipe_phv_in_data_151; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_152 = io_pipe_phv_in_data_152; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_153 = io_pipe_phv_in_data_153; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_154 = io_pipe_phv_in_data_154; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_155 = io_pipe_phv_in_data_155; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_156 = io_pipe_phv_in_data_156; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_157 = io_pipe_phv_in_data_157; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_158 = io_pipe_phv_in_data_158; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_159 = io_pipe_phv_in_data_159; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_160 = io_pipe_phv_in_data_160; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_161 = io_pipe_phv_in_data_161; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_162 = io_pipe_phv_in_data_162; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_163 = io_pipe_phv_in_data_163; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_164 = io_pipe_phv_in_data_164; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_165 = io_pipe_phv_in_data_165; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_166 = io_pipe_phv_in_data_166; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_167 = io_pipe_phv_in_data_167; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_168 = io_pipe_phv_in_data_168; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_169 = io_pipe_phv_in_data_169; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_170 = io_pipe_phv_in_data_170; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_171 = io_pipe_phv_in_data_171; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_172 = io_pipe_phv_in_data_172; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_173 = io_pipe_phv_in_data_173; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_174 = io_pipe_phv_in_data_174; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_175 = io_pipe_phv_in_data_175; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_176 = io_pipe_phv_in_data_176; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_177 = io_pipe_phv_in_data_177; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_178 = io_pipe_phv_in_data_178; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_179 = io_pipe_phv_in_data_179; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_180 = io_pipe_phv_in_data_180; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_181 = io_pipe_phv_in_data_181; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_182 = io_pipe_phv_in_data_182; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_183 = io_pipe_phv_in_data_183; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_184 = io_pipe_phv_in_data_184; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_185 = io_pipe_phv_in_data_185; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_186 = io_pipe_phv_in_data_186; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_187 = io_pipe_phv_in_data_187; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_188 = io_pipe_phv_in_data_188; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_189 = io_pipe_phv_in_data_189; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_190 = io_pipe_phv_in_data_190; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_191 = io_pipe_phv_in_data_191; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_192 = io_pipe_phv_in_data_192; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_193 = io_pipe_phv_in_data_193; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_194 = io_pipe_phv_in_data_194; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_195 = io_pipe_phv_in_data_195; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_196 = io_pipe_phv_in_data_196; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_197 = io_pipe_phv_in_data_197; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_198 = io_pipe_phv_in_data_198; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_199 = io_pipe_phv_in_data_199; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_200 = io_pipe_phv_in_data_200; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_201 = io_pipe_phv_in_data_201; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_202 = io_pipe_phv_in_data_202; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_203 = io_pipe_phv_in_data_203; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_204 = io_pipe_phv_in_data_204; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_205 = io_pipe_phv_in_data_205; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_206 = io_pipe_phv_in_data_206; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_207 = io_pipe_phv_in_data_207; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_208 = io_pipe_phv_in_data_208; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_209 = io_pipe_phv_in_data_209; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_210 = io_pipe_phv_in_data_210; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_211 = io_pipe_phv_in_data_211; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_212 = io_pipe_phv_in_data_212; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_213 = io_pipe_phv_in_data_213; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_214 = io_pipe_phv_in_data_214; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_215 = io_pipe_phv_in_data_215; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_216 = io_pipe_phv_in_data_216; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_217 = io_pipe_phv_in_data_217; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_218 = io_pipe_phv_in_data_218; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_219 = io_pipe_phv_in_data_219; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_220 = io_pipe_phv_in_data_220; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_221 = io_pipe_phv_in_data_221; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_222 = io_pipe_phv_in_data_222; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_223 = io_pipe_phv_in_data_223; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_224 = io_pipe_phv_in_data_224; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_225 = io_pipe_phv_in_data_225; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_226 = io_pipe_phv_in_data_226; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_227 = io_pipe_phv_in_data_227; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_228 = io_pipe_phv_in_data_228; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_229 = io_pipe_phv_in_data_229; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_230 = io_pipe_phv_in_data_230; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_231 = io_pipe_phv_in_data_231; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_232 = io_pipe_phv_in_data_232; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_233 = io_pipe_phv_in_data_233; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_234 = io_pipe_phv_in_data_234; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_235 = io_pipe_phv_in_data_235; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_236 = io_pipe_phv_in_data_236; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_237 = io_pipe_phv_in_data_237; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_238 = io_pipe_phv_in_data_238; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_239 = io_pipe_phv_in_data_239; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_240 = io_pipe_phv_in_data_240; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_241 = io_pipe_phv_in_data_241; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_242 = io_pipe_phv_in_data_242; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_243 = io_pipe_phv_in_data_243; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_244 = io_pipe_phv_in_data_244; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_245 = io_pipe_phv_in_data_245; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_246 = io_pipe_phv_in_data_246; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_247 = io_pipe_phv_in_data_247; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_248 = io_pipe_phv_in_data_248; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_249 = io_pipe_phv_in_data_249; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_250 = io_pipe_phv_in_data_250; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_251 = io_pipe_phv_in_data_251; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_252 = io_pipe_phv_in_data_252; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_253 = io_pipe_phv_in_data_253; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_254 = io_pipe_phv_in_data_254; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_data_255 = io_pipe_phv_in_data_255; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_next_processor_id = io_pipe_phv_in_next_processor_id; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_next_config_id = io_pipe_phv_in_next_config_id; // @[processor_pisa.scala 25:24]
  assign MAT_io_pipe_phv_in_is_valid_processor = io_pipe_phv_in_is_valid_processor; // @[processor_pisa.scala 25:24]
  assign MAT_io_mod_en = io_mod_mat_mod_en; // @[processor_pisa.scala 26:24]
  assign MAT_io_mod_config_id = io_mod_mat_mod_config_id; // @[processor_pisa.scala 26:24]
  assign MAT_io_mod_key_mod_en = io_mod_mat_mod_key_mod_en; // @[processor_pisa.scala 26:24]
  assign MAT_io_mod_key_mod_group_index = io_mod_mat_mod_key_mod_group_index; // @[processor_pisa.scala 26:24]
  assign MAT_io_mod_key_mod_group_config = io_mod_mat_mod_key_mod_group_config; // @[processor_pisa.scala 26:24]
  assign MAT_io_mod_key_mod_group_mask_0 = io_mod_mat_mod_key_mod_group_mask_0; // @[processor_pisa.scala 26:24]
  assign MAT_io_mod_key_mod_group_mask_1 = io_mod_mat_mod_key_mod_group_mask_1; // @[processor_pisa.scala 26:24]
  assign MAT_io_mod_key_mod_group_mask_2 = io_mod_mat_mod_key_mod_group_mask_2; // @[processor_pisa.scala 26:24]
  assign MAT_io_mod_key_mod_group_mask_3 = io_mod_mat_mod_key_mod_group_mask_3; // @[processor_pisa.scala 26:24]
  assign MAT_io_mod_key_mod_group_id_0 = io_mod_mat_mod_key_mod_group_id_0; // @[processor_pisa.scala 26:24]
  assign MAT_io_mod_key_mod_group_id_1 = io_mod_mat_mod_key_mod_group_id_1; // @[processor_pisa.scala 26:24]
  assign MAT_io_mod_key_mod_group_id_2 = io_mod_mat_mod_key_mod_group_id_2; // @[processor_pisa.scala 26:24]
  assign MAT_io_mod_key_mod_group_id_3 = io_mod_mat_mod_key_mod_group_id_3; // @[processor_pisa.scala 26:24]
  assign MAT_io_mod_table_mod_table_depth = io_mod_mat_mod_table_mod_table_depth; // @[processor_pisa.scala 26:24]
  assign MAT_io_mod_table_mod_table_width = io_mod_mat_mod_table_mod_table_width; // @[processor_pisa.scala 26:24]
  assign MAT_io_mod_w_en = io_mod_mat_mod_w_en; // @[processor_pisa.scala 26:24]
  assign MAT_io_mod_w_sram_id = io_mod_mat_mod_w_sram_id; // @[processor_pisa.scala 26:24]
  assign MAT_io_mod_w_addr = io_mod_mat_mod_w_addr; // @[processor_pisa.scala 26:24]
  assign MAT_io_mod_w_data = io_mod_mat_mod_w_data; // @[processor_pisa.scala 26:24]
  assign EXE_clock = clock;
  assign EXE_io_pipe_phv_in_data_0 = MAT_io_pipe_phv_out_data_0; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_1 = MAT_io_pipe_phv_out_data_1; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_2 = MAT_io_pipe_phv_out_data_2; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_3 = MAT_io_pipe_phv_out_data_3; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_4 = MAT_io_pipe_phv_out_data_4; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_5 = MAT_io_pipe_phv_out_data_5; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_6 = MAT_io_pipe_phv_out_data_6; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_7 = MAT_io_pipe_phv_out_data_7; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_8 = MAT_io_pipe_phv_out_data_8; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_9 = MAT_io_pipe_phv_out_data_9; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_10 = MAT_io_pipe_phv_out_data_10; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_11 = MAT_io_pipe_phv_out_data_11; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_12 = MAT_io_pipe_phv_out_data_12; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_13 = MAT_io_pipe_phv_out_data_13; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_14 = MAT_io_pipe_phv_out_data_14; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_15 = MAT_io_pipe_phv_out_data_15; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_16 = MAT_io_pipe_phv_out_data_16; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_17 = MAT_io_pipe_phv_out_data_17; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_18 = MAT_io_pipe_phv_out_data_18; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_19 = MAT_io_pipe_phv_out_data_19; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_20 = MAT_io_pipe_phv_out_data_20; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_21 = MAT_io_pipe_phv_out_data_21; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_22 = MAT_io_pipe_phv_out_data_22; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_23 = MAT_io_pipe_phv_out_data_23; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_24 = MAT_io_pipe_phv_out_data_24; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_25 = MAT_io_pipe_phv_out_data_25; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_26 = MAT_io_pipe_phv_out_data_26; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_27 = MAT_io_pipe_phv_out_data_27; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_28 = MAT_io_pipe_phv_out_data_28; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_29 = MAT_io_pipe_phv_out_data_29; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_30 = MAT_io_pipe_phv_out_data_30; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_31 = MAT_io_pipe_phv_out_data_31; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_32 = MAT_io_pipe_phv_out_data_32; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_33 = MAT_io_pipe_phv_out_data_33; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_34 = MAT_io_pipe_phv_out_data_34; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_35 = MAT_io_pipe_phv_out_data_35; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_36 = MAT_io_pipe_phv_out_data_36; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_37 = MAT_io_pipe_phv_out_data_37; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_38 = MAT_io_pipe_phv_out_data_38; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_39 = MAT_io_pipe_phv_out_data_39; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_40 = MAT_io_pipe_phv_out_data_40; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_41 = MAT_io_pipe_phv_out_data_41; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_42 = MAT_io_pipe_phv_out_data_42; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_43 = MAT_io_pipe_phv_out_data_43; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_44 = MAT_io_pipe_phv_out_data_44; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_45 = MAT_io_pipe_phv_out_data_45; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_46 = MAT_io_pipe_phv_out_data_46; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_47 = MAT_io_pipe_phv_out_data_47; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_48 = MAT_io_pipe_phv_out_data_48; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_49 = MAT_io_pipe_phv_out_data_49; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_50 = MAT_io_pipe_phv_out_data_50; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_51 = MAT_io_pipe_phv_out_data_51; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_52 = MAT_io_pipe_phv_out_data_52; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_53 = MAT_io_pipe_phv_out_data_53; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_54 = MAT_io_pipe_phv_out_data_54; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_55 = MAT_io_pipe_phv_out_data_55; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_56 = MAT_io_pipe_phv_out_data_56; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_57 = MAT_io_pipe_phv_out_data_57; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_58 = MAT_io_pipe_phv_out_data_58; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_59 = MAT_io_pipe_phv_out_data_59; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_60 = MAT_io_pipe_phv_out_data_60; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_61 = MAT_io_pipe_phv_out_data_61; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_62 = MAT_io_pipe_phv_out_data_62; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_63 = MAT_io_pipe_phv_out_data_63; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_64 = MAT_io_pipe_phv_out_data_64; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_65 = MAT_io_pipe_phv_out_data_65; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_66 = MAT_io_pipe_phv_out_data_66; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_67 = MAT_io_pipe_phv_out_data_67; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_68 = MAT_io_pipe_phv_out_data_68; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_69 = MAT_io_pipe_phv_out_data_69; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_70 = MAT_io_pipe_phv_out_data_70; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_71 = MAT_io_pipe_phv_out_data_71; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_72 = MAT_io_pipe_phv_out_data_72; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_73 = MAT_io_pipe_phv_out_data_73; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_74 = MAT_io_pipe_phv_out_data_74; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_75 = MAT_io_pipe_phv_out_data_75; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_76 = MAT_io_pipe_phv_out_data_76; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_77 = MAT_io_pipe_phv_out_data_77; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_78 = MAT_io_pipe_phv_out_data_78; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_79 = MAT_io_pipe_phv_out_data_79; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_80 = MAT_io_pipe_phv_out_data_80; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_81 = MAT_io_pipe_phv_out_data_81; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_82 = MAT_io_pipe_phv_out_data_82; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_83 = MAT_io_pipe_phv_out_data_83; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_84 = MAT_io_pipe_phv_out_data_84; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_85 = MAT_io_pipe_phv_out_data_85; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_86 = MAT_io_pipe_phv_out_data_86; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_87 = MAT_io_pipe_phv_out_data_87; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_88 = MAT_io_pipe_phv_out_data_88; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_89 = MAT_io_pipe_phv_out_data_89; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_90 = MAT_io_pipe_phv_out_data_90; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_91 = MAT_io_pipe_phv_out_data_91; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_92 = MAT_io_pipe_phv_out_data_92; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_93 = MAT_io_pipe_phv_out_data_93; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_94 = MAT_io_pipe_phv_out_data_94; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_95 = MAT_io_pipe_phv_out_data_95; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_96 = MAT_io_pipe_phv_out_data_96; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_97 = MAT_io_pipe_phv_out_data_97; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_98 = MAT_io_pipe_phv_out_data_98; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_99 = MAT_io_pipe_phv_out_data_99; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_100 = MAT_io_pipe_phv_out_data_100; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_101 = MAT_io_pipe_phv_out_data_101; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_102 = MAT_io_pipe_phv_out_data_102; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_103 = MAT_io_pipe_phv_out_data_103; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_104 = MAT_io_pipe_phv_out_data_104; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_105 = MAT_io_pipe_phv_out_data_105; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_106 = MAT_io_pipe_phv_out_data_106; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_107 = MAT_io_pipe_phv_out_data_107; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_108 = MAT_io_pipe_phv_out_data_108; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_109 = MAT_io_pipe_phv_out_data_109; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_110 = MAT_io_pipe_phv_out_data_110; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_111 = MAT_io_pipe_phv_out_data_111; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_112 = MAT_io_pipe_phv_out_data_112; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_113 = MAT_io_pipe_phv_out_data_113; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_114 = MAT_io_pipe_phv_out_data_114; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_115 = MAT_io_pipe_phv_out_data_115; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_116 = MAT_io_pipe_phv_out_data_116; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_117 = MAT_io_pipe_phv_out_data_117; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_118 = MAT_io_pipe_phv_out_data_118; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_119 = MAT_io_pipe_phv_out_data_119; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_120 = MAT_io_pipe_phv_out_data_120; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_121 = MAT_io_pipe_phv_out_data_121; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_122 = MAT_io_pipe_phv_out_data_122; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_123 = MAT_io_pipe_phv_out_data_123; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_124 = MAT_io_pipe_phv_out_data_124; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_125 = MAT_io_pipe_phv_out_data_125; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_126 = MAT_io_pipe_phv_out_data_126; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_127 = MAT_io_pipe_phv_out_data_127; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_128 = MAT_io_pipe_phv_out_data_128; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_129 = MAT_io_pipe_phv_out_data_129; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_130 = MAT_io_pipe_phv_out_data_130; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_131 = MAT_io_pipe_phv_out_data_131; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_132 = MAT_io_pipe_phv_out_data_132; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_133 = MAT_io_pipe_phv_out_data_133; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_134 = MAT_io_pipe_phv_out_data_134; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_135 = MAT_io_pipe_phv_out_data_135; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_136 = MAT_io_pipe_phv_out_data_136; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_137 = MAT_io_pipe_phv_out_data_137; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_138 = MAT_io_pipe_phv_out_data_138; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_139 = MAT_io_pipe_phv_out_data_139; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_140 = MAT_io_pipe_phv_out_data_140; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_141 = MAT_io_pipe_phv_out_data_141; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_142 = MAT_io_pipe_phv_out_data_142; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_143 = MAT_io_pipe_phv_out_data_143; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_144 = MAT_io_pipe_phv_out_data_144; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_145 = MAT_io_pipe_phv_out_data_145; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_146 = MAT_io_pipe_phv_out_data_146; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_147 = MAT_io_pipe_phv_out_data_147; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_148 = MAT_io_pipe_phv_out_data_148; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_149 = MAT_io_pipe_phv_out_data_149; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_150 = MAT_io_pipe_phv_out_data_150; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_151 = MAT_io_pipe_phv_out_data_151; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_152 = MAT_io_pipe_phv_out_data_152; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_153 = MAT_io_pipe_phv_out_data_153; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_154 = MAT_io_pipe_phv_out_data_154; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_155 = MAT_io_pipe_phv_out_data_155; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_156 = MAT_io_pipe_phv_out_data_156; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_157 = MAT_io_pipe_phv_out_data_157; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_158 = MAT_io_pipe_phv_out_data_158; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_159 = MAT_io_pipe_phv_out_data_159; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_160 = MAT_io_pipe_phv_out_data_160; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_161 = MAT_io_pipe_phv_out_data_161; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_162 = MAT_io_pipe_phv_out_data_162; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_163 = MAT_io_pipe_phv_out_data_163; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_164 = MAT_io_pipe_phv_out_data_164; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_165 = MAT_io_pipe_phv_out_data_165; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_166 = MAT_io_pipe_phv_out_data_166; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_167 = MAT_io_pipe_phv_out_data_167; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_168 = MAT_io_pipe_phv_out_data_168; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_169 = MAT_io_pipe_phv_out_data_169; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_170 = MAT_io_pipe_phv_out_data_170; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_171 = MAT_io_pipe_phv_out_data_171; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_172 = MAT_io_pipe_phv_out_data_172; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_173 = MAT_io_pipe_phv_out_data_173; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_174 = MAT_io_pipe_phv_out_data_174; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_175 = MAT_io_pipe_phv_out_data_175; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_176 = MAT_io_pipe_phv_out_data_176; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_177 = MAT_io_pipe_phv_out_data_177; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_178 = MAT_io_pipe_phv_out_data_178; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_179 = MAT_io_pipe_phv_out_data_179; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_180 = MAT_io_pipe_phv_out_data_180; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_181 = MAT_io_pipe_phv_out_data_181; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_182 = MAT_io_pipe_phv_out_data_182; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_183 = MAT_io_pipe_phv_out_data_183; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_184 = MAT_io_pipe_phv_out_data_184; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_185 = MAT_io_pipe_phv_out_data_185; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_186 = MAT_io_pipe_phv_out_data_186; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_187 = MAT_io_pipe_phv_out_data_187; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_188 = MAT_io_pipe_phv_out_data_188; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_189 = MAT_io_pipe_phv_out_data_189; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_190 = MAT_io_pipe_phv_out_data_190; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_191 = MAT_io_pipe_phv_out_data_191; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_192 = MAT_io_pipe_phv_out_data_192; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_193 = MAT_io_pipe_phv_out_data_193; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_194 = MAT_io_pipe_phv_out_data_194; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_195 = MAT_io_pipe_phv_out_data_195; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_196 = MAT_io_pipe_phv_out_data_196; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_197 = MAT_io_pipe_phv_out_data_197; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_198 = MAT_io_pipe_phv_out_data_198; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_199 = MAT_io_pipe_phv_out_data_199; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_200 = MAT_io_pipe_phv_out_data_200; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_201 = MAT_io_pipe_phv_out_data_201; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_202 = MAT_io_pipe_phv_out_data_202; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_203 = MAT_io_pipe_phv_out_data_203; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_204 = MAT_io_pipe_phv_out_data_204; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_205 = MAT_io_pipe_phv_out_data_205; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_206 = MAT_io_pipe_phv_out_data_206; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_207 = MAT_io_pipe_phv_out_data_207; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_208 = MAT_io_pipe_phv_out_data_208; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_209 = MAT_io_pipe_phv_out_data_209; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_210 = MAT_io_pipe_phv_out_data_210; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_211 = MAT_io_pipe_phv_out_data_211; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_212 = MAT_io_pipe_phv_out_data_212; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_213 = MAT_io_pipe_phv_out_data_213; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_214 = MAT_io_pipe_phv_out_data_214; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_215 = MAT_io_pipe_phv_out_data_215; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_216 = MAT_io_pipe_phv_out_data_216; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_217 = MAT_io_pipe_phv_out_data_217; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_218 = MAT_io_pipe_phv_out_data_218; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_219 = MAT_io_pipe_phv_out_data_219; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_220 = MAT_io_pipe_phv_out_data_220; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_221 = MAT_io_pipe_phv_out_data_221; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_222 = MAT_io_pipe_phv_out_data_222; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_223 = MAT_io_pipe_phv_out_data_223; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_224 = MAT_io_pipe_phv_out_data_224; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_225 = MAT_io_pipe_phv_out_data_225; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_226 = MAT_io_pipe_phv_out_data_226; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_227 = MAT_io_pipe_phv_out_data_227; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_228 = MAT_io_pipe_phv_out_data_228; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_229 = MAT_io_pipe_phv_out_data_229; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_230 = MAT_io_pipe_phv_out_data_230; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_231 = MAT_io_pipe_phv_out_data_231; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_232 = MAT_io_pipe_phv_out_data_232; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_233 = MAT_io_pipe_phv_out_data_233; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_234 = MAT_io_pipe_phv_out_data_234; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_235 = MAT_io_pipe_phv_out_data_235; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_236 = MAT_io_pipe_phv_out_data_236; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_237 = MAT_io_pipe_phv_out_data_237; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_238 = MAT_io_pipe_phv_out_data_238; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_239 = MAT_io_pipe_phv_out_data_239; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_240 = MAT_io_pipe_phv_out_data_240; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_241 = MAT_io_pipe_phv_out_data_241; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_242 = MAT_io_pipe_phv_out_data_242; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_243 = MAT_io_pipe_phv_out_data_243; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_244 = MAT_io_pipe_phv_out_data_244; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_245 = MAT_io_pipe_phv_out_data_245; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_246 = MAT_io_pipe_phv_out_data_246; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_247 = MAT_io_pipe_phv_out_data_247; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_248 = MAT_io_pipe_phv_out_data_248; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_249 = MAT_io_pipe_phv_out_data_249; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_250 = MAT_io_pipe_phv_out_data_250; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_251 = MAT_io_pipe_phv_out_data_251; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_252 = MAT_io_pipe_phv_out_data_252; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_253 = MAT_io_pipe_phv_out_data_253; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_254 = MAT_io_pipe_phv_out_data_254; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_data_255 = MAT_io_pipe_phv_out_data_255; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_next_processor_id = MAT_io_pipe_phv_out_next_processor_id; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_next_config_id = MAT_io_pipe_phv_out_next_config_id; // @[processor_pisa.scala 28:24]
  assign EXE_io_pipe_phv_in_is_valid_processor = MAT_io_pipe_phv_out_is_valid_processor; // @[processor_pisa.scala 28:24]
  assign EXE_io_hit = MAT_io_hit; // @[processor_pisa.scala 29:24]
  assign EXE_io_match_value = MAT_io_match_value; // @[processor_pisa.scala 30:24]
  assign EXE_io_action_mod_en_0 = io_mod_exe_mod_en_0; // @[processor_pisa.scala 31:24]
  assign EXE_io_action_mod_en_1 = io_mod_exe_mod_en_1; // @[processor_pisa.scala 31:24]
  assign EXE_io_action_mod_addr = io_mod_exe_mod_addr; // @[processor_pisa.scala 31:24]
  assign EXE_io_action_mod_data_0 = io_mod_exe_mod_data_0; // @[processor_pisa.scala 31:24]
  assign EXE_io_action_mod_data_1 = io_mod_exe_mod_data_1; // @[processor_pisa.scala 31:24]
endmodule
