module MatchGetKeyRaw(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [3:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [3:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input  [7:0]  io_key_config_0_key_length,
  input  [7:0]  io_key_config_1_key_length,
  input  [7:0]  io_key_offset_in,
  output [1:0]  io_bias_out,
  output [7:0]  io_match_key_bytes_0,
  output [7:0]  io_match_key_bytes_1,
  output [7:0]  io_match_key_bytes_2,
  output [7:0]  io_match_key_bytes_3,
  output [7:0]  io_match_key_bytes_4,
  output [7:0]  io_match_key_bytes_5,
  output [7:0]  io_match_key_bytes_6,
  output [7:0]  io_match_key_bytes_7,
  output [7:0]  io_match_key_bytes_8,
  output [7:0]  io_match_key_bytes_9,
  output [7:0]  io_match_key_bytes_10,
  output [7:0]  io_match_key_bytes_11,
  output [7:0]  io_match_key_bytes_12,
  output [7:0]  io_match_key_bytes_13,
  output [7:0]  io_match_key_bytes_14,
  output [7:0]  io_match_key_bytes_15,
  output [7:0]  io_match_key_bytes_16,
  output [7:0]  io_match_key_bytes_17,
  output [7:0]  io_match_key_bytes_18,
  output [7:0]  io_match_key_bytes_19,
  output [7:0]  io_match_key_bytes_20,
  output [7:0]  io_match_key_bytes_21,
  output [7:0]  io_match_key_bytes_22,
  output [7:0]  io_match_key_bytes_23
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[matcher.scala 67:26]
  reg [7:0] phv_data_1; // @[matcher.scala 67:26]
  reg [7:0] phv_data_2; // @[matcher.scala 67:26]
  reg [7:0] phv_data_3; // @[matcher.scala 67:26]
  reg [7:0] phv_data_4; // @[matcher.scala 67:26]
  reg [7:0] phv_data_5; // @[matcher.scala 67:26]
  reg [7:0] phv_data_6; // @[matcher.scala 67:26]
  reg [7:0] phv_data_7; // @[matcher.scala 67:26]
  reg [7:0] phv_data_8; // @[matcher.scala 67:26]
  reg [7:0] phv_data_9; // @[matcher.scala 67:26]
  reg [7:0] phv_data_10; // @[matcher.scala 67:26]
  reg [7:0] phv_data_11; // @[matcher.scala 67:26]
  reg [7:0] phv_data_12; // @[matcher.scala 67:26]
  reg [7:0] phv_data_13; // @[matcher.scala 67:26]
  reg [7:0] phv_data_14; // @[matcher.scala 67:26]
  reg [7:0] phv_data_15; // @[matcher.scala 67:26]
  reg [7:0] phv_data_16; // @[matcher.scala 67:26]
  reg [7:0] phv_data_17; // @[matcher.scala 67:26]
  reg [7:0] phv_data_18; // @[matcher.scala 67:26]
  reg [7:0] phv_data_19; // @[matcher.scala 67:26]
  reg [7:0] phv_data_20; // @[matcher.scala 67:26]
  reg [7:0] phv_data_21; // @[matcher.scala 67:26]
  reg [7:0] phv_data_22; // @[matcher.scala 67:26]
  reg [7:0] phv_data_23; // @[matcher.scala 67:26]
  reg [7:0] phv_data_24; // @[matcher.scala 67:26]
  reg [7:0] phv_data_25; // @[matcher.scala 67:26]
  reg [7:0] phv_data_26; // @[matcher.scala 67:26]
  reg [7:0] phv_data_27; // @[matcher.scala 67:26]
  reg [7:0] phv_data_28; // @[matcher.scala 67:26]
  reg [7:0] phv_data_29; // @[matcher.scala 67:26]
  reg [7:0] phv_data_30; // @[matcher.scala 67:26]
  reg [7:0] phv_data_31; // @[matcher.scala 67:26]
  reg [7:0] phv_data_32; // @[matcher.scala 67:26]
  reg [7:0] phv_data_33; // @[matcher.scala 67:26]
  reg [7:0] phv_data_34; // @[matcher.scala 67:26]
  reg [7:0] phv_data_35; // @[matcher.scala 67:26]
  reg [7:0] phv_data_36; // @[matcher.scala 67:26]
  reg [7:0] phv_data_37; // @[matcher.scala 67:26]
  reg [7:0] phv_data_38; // @[matcher.scala 67:26]
  reg [7:0] phv_data_39; // @[matcher.scala 67:26]
  reg [7:0] phv_data_40; // @[matcher.scala 67:26]
  reg [7:0] phv_data_41; // @[matcher.scala 67:26]
  reg [7:0] phv_data_42; // @[matcher.scala 67:26]
  reg [7:0] phv_data_43; // @[matcher.scala 67:26]
  reg [7:0] phv_data_44; // @[matcher.scala 67:26]
  reg [7:0] phv_data_45; // @[matcher.scala 67:26]
  reg [7:0] phv_data_46; // @[matcher.scala 67:26]
  reg [7:0] phv_data_47; // @[matcher.scala 67:26]
  reg [7:0] phv_data_48; // @[matcher.scala 67:26]
  reg [7:0] phv_data_49; // @[matcher.scala 67:26]
  reg [7:0] phv_data_50; // @[matcher.scala 67:26]
  reg [7:0] phv_data_51; // @[matcher.scala 67:26]
  reg [7:0] phv_data_52; // @[matcher.scala 67:26]
  reg [7:0] phv_data_53; // @[matcher.scala 67:26]
  reg [7:0] phv_data_54; // @[matcher.scala 67:26]
  reg [7:0] phv_data_55; // @[matcher.scala 67:26]
  reg [7:0] phv_data_56; // @[matcher.scala 67:26]
  reg [7:0] phv_data_57; // @[matcher.scala 67:26]
  reg [7:0] phv_data_58; // @[matcher.scala 67:26]
  reg [7:0] phv_data_59; // @[matcher.scala 67:26]
  reg [7:0] phv_data_60; // @[matcher.scala 67:26]
  reg [7:0] phv_data_61; // @[matcher.scala 67:26]
  reg [7:0] phv_data_62; // @[matcher.scala 67:26]
  reg [7:0] phv_data_63; // @[matcher.scala 67:26]
  reg [7:0] phv_data_64; // @[matcher.scala 67:26]
  reg [7:0] phv_data_65; // @[matcher.scala 67:26]
  reg [7:0] phv_data_66; // @[matcher.scala 67:26]
  reg [7:0] phv_data_67; // @[matcher.scala 67:26]
  reg [7:0] phv_data_68; // @[matcher.scala 67:26]
  reg [7:0] phv_data_69; // @[matcher.scala 67:26]
  reg [7:0] phv_data_70; // @[matcher.scala 67:26]
  reg [7:0] phv_data_71; // @[matcher.scala 67:26]
  reg [7:0] phv_data_72; // @[matcher.scala 67:26]
  reg [7:0] phv_data_73; // @[matcher.scala 67:26]
  reg [7:0] phv_data_74; // @[matcher.scala 67:26]
  reg [7:0] phv_data_75; // @[matcher.scala 67:26]
  reg [7:0] phv_data_76; // @[matcher.scala 67:26]
  reg [7:0] phv_data_77; // @[matcher.scala 67:26]
  reg [7:0] phv_data_78; // @[matcher.scala 67:26]
  reg [7:0] phv_data_79; // @[matcher.scala 67:26]
  reg [7:0] phv_data_80; // @[matcher.scala 67:26]
  reg [7:0] phv_data_81; // @[matcher.scala 67:26]
  reg [7:0] phv_data_82; // @[matcher.scala 67:26]
  reg [7:0] phv_data_83; // @[matcher.scala 67:26]
  reg [7:0] phv_data_84; // @[matcher.scala 67:26]
  reg [7:0] phv_data_85; // @[matcher.scala 67:26]
  reg [7:0] phv_data_86; // @[matcher.scala 67:26]
  reg [7:0] phv_data_87; // @[matcher.scala 67:26]
  reg [7:0] phv_data_88; // @[matcher.scala 67:26]
  reg [7:0] phv_data_89; // @[matcher.scala 67:26]
  reg [7:0] phv_data_90; // @[matcher.scala 67:26]
  reg [7:0] phv_data_91; // @[matcher.scala 67:26]
  reg [7:0] phv_data_92; // @[matcher.scala 67:26]
  reg [7:0] phv_data_93; // @[matcher.scala 67:26]
  reg [7:0] phv_data_94; // @[matcher.scala 67:26]
  reg [7:0] phv_data_95; // @[matcher.scala 67:26]
  reg [7:0] phv_data_96; // @[matcher.scala 67:26]
  reg [7:0] phv_data_97; // @[matcher.scala 67:26]
  reg [7:0] phv_data_98; // @[matcher.scala 67:26]
  reg [7:0] phv_data_99; // @[matcher.scala 67:26]
  reg [7:0] phv_data_100; // @[matcher.scala 67:26]
  reg [7:0] phv_data_101; // @[matcher.scala 67:26]
  reg [7:0] phv_data_102; // @[matcher.scala 67:26]
  reg [7:0] phv_data_103; // @[matcher.scala 67:26]
  reg [7:0] phv_data_104; // @[matcher.scala 67:26]
  reg [7:0] phv_data_105; // @[matcher.scala 67:26]
  reg [7:0] phv_data_106; // @[matcher.scala 67:26]
  reg [7:0] phv_data_107; // @[matcher.scala 67:26]
  reg [7:0] phv_data_108; // @[matcher.scala 67:26]
  reg [7:0] phv_data_109; // @[matcher.scala 67:26]
  reg [7:0] phv_data_110; // @[matcher.scala 67:26]
  reg [7:0] phv_data_111; // @[matcher.scala 67:26]
  reg [7:0] phv_data_112; // @[matcher.scala 67:26]
  reg [7:0] phv_data_113; // @[matcher.scala 67:26]
  reg [7:0] phv_data_114; // @[matcher.scala 67:26]
  reg [7:0] phv_data_115; // @[matcher.scala 67:26]
  reg [7:0] phv_data_116; // @[matcher.scala 67:26]
  reg [7:0] phv_data_117; // @[matcher.scala 67:26]
  reg [7:0] phv_data_118; // @[matcher.scala 67:26]
  reg [7:0] phv_data_119; // @[matcher.scala 67:26]
  reg [7:0] phv_data_120; // @[matcher.scala 67:26]
  reg [7:0] phv_data_121; // @[matcher.scala 67:26]
  reg [7:0] phv_data_122; // @[matcher.scala 67:26]
  reg [7:0] phv_data_123; // @[matcher.scala 67:26]
  reg [7:0] phv_data_124; // @[matcher.scala 67:26]
  reg [7:0] phv_data_125; // @[matcher.scala 67:26]
  reg [7:0] phv_data_126; // @[matcher.scala 67:26]
  reg [7:0] phv_data_127; // @[matcher.scala 67:26]
  reg [7:0] phv_data_128; // @[matcher.scala 67:26]
  reg [7:0] phv_data_129; // @[matcher.scala 67:26]
  reg [7:0] phv_data_130; // @[matcher.scala 67:26]
  reg [7:0] phv_data_131; // @[matcher.scala 67:26]
  reg [7:0] phv_data_132; // @[matcher.scala 67:26]
  reg [7:0] phv_data_133; // @[matcher.scala 67:26]
  reg [7:0] phv_data_134; // @[matcher.scala 67:26]
  reg [7:0] phv_data_135; // @[matcher.scala 67:26]
  reg [7:0] phv_data_136; // @[matcher.scala 67:26]
  reg [7:0] phv_data_137; // @[matcher.scala 67:26]
  reg [7:0] phv_data_138; // @[matcher.scala 67:26]
  reg [7:0] phv_data_139; // @[matcher.scala 67:26]
  reg [7:0] phv_data_140; // @[matcher.scala 67:26]
  reg [7:0] phv_data_141; // @[matcher.scala 67:26]
  reg [7:0] phv_data_142; // @[matcher.scala 67:26]
  reg [7:0] phv_data_143; // @[matcher.scala 67:26]
  reg [7:0] phv_data_144; // @[matcher.scala 67:26]
  reg [7:0] phv_data_145; // @[matcher.scala 67:26]
  reg [7:0] phv_data_146; // @[matcher.scala 67:26]
  reg [7:0] phv_data_147; // @[matcher.scala 67:26]
  reg [7:0] phv_data_148; // @[matcher.scala 67:26]
  reg [7:0] phv_data_149; // @[matcher.scala 67:26]
  reg [7:0] phv_data_150; // @[matcher.scala 67:26]
  reg [7:0] phv_data_151; // @[matcher.scala 67:26]
  reg [7:0] phv_data_152; // @[matcher.scala 67:26]
  reg [7:0] phv_data_153; // @[matcher.scala 67:26]
  reg [7:0] phv_data_154; // @[matcher.scala 67:26]
  reg [7:0] phv_data_155; // @[matcher.scala 67:26]
  reg [7:0] phv_data_156; // @[matcher.scala 67:26]
  reg [7:0] phv_data_157; // @[matcher.scala 67:26]
  reg [7:0] phv_data_158; // @[matcher.scala 67:26]
  reg [7:0] phv_data_159; // @[matcher.scala 67:26]
  reg [15:0] phv_header_0; // @[matcher.scala 67:26]
  reg [15:0] phv_header_1; // @[matcher.scala 67:26]
  reg [15:0] phv_header_2; // @[matcher.scala 67:26]
  reg [15:0] phv_header_3; // @[matcher.scala 67:26]
  reg [15:0] phv_header_4; // @[matcher.scala 67:26]
  reg [15:0] phv_header_5; // @[matcher.scala 67:26]
  reg [15:0] phv_header_6; // @[matcher.scala 67:26]
  reg [15:0] phv_header_7; // @[matcher.scala 67:26]
  reg [15:0] phv_header_8; // @[matcher.scala 67:26]
  reg [15:0] phv_header_9; // @[matcher.scala 67:26]
  reg [15:0] phv_header_10; // @[matcher.scala 67:26]
  reg [15:0] phv_header_11; // @[matcher.scala 67:26]
  reg [15:0] phv_header_12; // @[matcher.scala 67:26]
  reg [15:0] phv_header_13; // @[matcher.scala 67:26]
  reg [15:0] phv_header_14; // @[matcher.scala 67:26]
  reg [15:0] phv_header_15; // @[matcher.scala 67:26]
  reg [7:0] phv_parse_current_state; // @[matcher.scala 67:26]
  reg [7:0] phv_parse_current_offset; // @[matcher.scala 67:26]
  reg [15:0] phv_parse_transition_field; // @[matcher.scala 67:26]
  reg [3:0] phv_next_processor_id; // @[matcher.scala 67:26]
  reg  phv_next_config_id; // @[matcher.scala 67:26]
  reg  phv_is_valid_processor; // @[matcher.scala 67:26]
  reg [7:0] key_offset; // @[matcher.scala 71:33]
  wire [5:0] read_key_offset_hi = key_offset[7:2]; // @[matcher.scala 73:49]
  wire [7:0] read_key_offset = {read_key_offset_hi,2'h0}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_6 = phv_next_config_id ? io_key_config_1_key_length : io_key_config_0_key_length; // @[matcher.scala 84:85 matcher.scala 84:85]
  wire [7:0] end_offset = _GEN_6 + key_offset; // @[matcher.scala 84:85]
  wire [8:0] _local_offset_T = {{1'd0}, read_key_offset}; // @[matcher.scala 87:77]
  wire [7:0] local_offset = _local_offset_T[7:0]; // @[matcher.scala 87:77]
  wire [5:0] match_key_qbytes_0_hi = local_offset[7:2]; // @[matcher.scala 91:54]
  wire [7:0] _match_key_qbytes_0_T = {match_key_qbytes_0_hi,2'h3}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_0_T_1 = {match_key_qbytes_0_hi,2'h2}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_0_T_2 = {match_key_qbytes_0_hi,2'h1}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_9 = 8'h1 == _match_key_qbytes_0_T_2 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10 = 8'h2 == _match_key_qbytes_0_T_2 ? phv_data_2 : _GEN_9; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11 = 8'h3 == _match_key_qbytes_0_T_2 ? phv_data_3 : _GEN_10; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12 = 8'h4 == _match_key_qbytes_0_T_2 ? phv_data_4 : _GEN_11; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_13 = 8'h5 == _match_key_qbytes_0_T_2 ? phv_data_5 : _GEN_12; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_14 = 8'h6 == _match_key_qbytes_0_T_2 ? phv_data_6 : _GEN_13; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_15 = 8'h7 == _match_key_qbytes_0_T_2 ? phv_data_7 : _GEN_14; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_16 = 8'h8 == _match_key_qbytes_0_T_2 ? phv_data_8 : _GEN_15; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_17 = 8'h9 == _match_key_qbytes_0_T_2 ? phv_data_9 : _GEN_16; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_18 = 8'ha == _match_key_qbytes_0_T_2 ? phv_data_10 : _GEN_17; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_19 = 8'hb == _match_key_qbytes_0_T_2 ? phv_data_11 : _GEN_18; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_20 = 8'hc == _match_key_qbytes_0_T_2 ? phv_data_12 : _GEN_19; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_21 = 8'hd == _match_key_qbytes_0_T_2 ? phv_data_13 : _GEN_20; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_22 = 8'he == _match_key_qbytes_0_T_2 ? phv_data_14 : _GEN_21; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_23 = 8'hf == _match_key_qbytes_0_T_2 ? phv_data_15 : _GEN_22; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_24 = 8'h10 == _match_key_qbytes_0_T_2 ? phv_data_16 : _GEN_23; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_25 = 8'h11 == _match_key_qbytes_0_T_2 ? phv_data_17 : _GEN_24; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_26 = 8'h12 == _match_key_qbytes_0_T_2 ? phv_data_18 : _GEN_25; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_27 = 8'h13 == _match_key_qbytes_0_T_2 ? phv_data_19 : _GEN_26; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_28 = 8'h14 == _match_key_qbytes_0_T_2 ? phv_data_20 : _GEN_27; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_29 = 8'h15 == _match_key_qbytes_0_T_2 ? phv_data_21 : _GEN_28; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_30 = 8'h16 == _match_key_qbytes_0_T_2 ? phv_data_22 : _GEN_29; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_31 = 8'h17 == _match_key_qbytes_0_T_2 ? phv_data_23 : _GEN_30; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_32 = 8'h18 == _match_key_qbytes_0_T_2 ? phv_data_24 : _GEN_31; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_33 = 8'h19 == _match_key_qbytes_0_T_2 ? phv_data_25 : _GEN_32; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_34 = 8'h1a == _match_key_qbytes_0_T_2 ? phv_data_26 : _GEN_33; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_35 = 8'h1b == _match_key_qbytes_0_T_2 ? phv_data_27 : _GEN_34; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_36 = 8'h1c == _match_key_qbytes_0_T_2 ? phv_data_28 : _GEN_35; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_37 = 8'h1d == _match_key_qbytes_0_T_2 ? phv_data_29 : _GEN_36; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_38 = 8'h1e == _match_key_qbytes_0_T_2 ? phv_data_30 : _GEN_37; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_39 = 8'h1f == _match_key_qbytes_0_T_2 ? phv_data_31 : _GEN_38; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_40 = 8'h20 == _match_key_qbytes_0_T_2 ? phv_data_32 : _GEN_39; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_41 = 8'h21 == _match_key_qbytes_0_T_2 ? phv_data_33 : _GEN_40; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_42 = 8'h22 == _match_key_qbytes_0_T_2 ? phv_data_34 : _GEN_41; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_43 = 8'h23 == _match_key_qbytes_0_T_2 ? phv_data_35 : _GEN_42; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_44 = 8'h24 == _match_key_qbytes_0_T_2 ? phv_data_36 : _GEN_43; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_45 = 8'h25 == _match_key_qbytes_0_T_2 ? phv_data_37 : _GEN_44; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_46 = 8'h26 == _match_key_qbytes_0_T_2 ? phv_data_38 : _GEN_45; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_47 = 8'h27 == _match_key_qbytes_0_T_2 ? phv_data_39 : _GEN_46; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_48 = 8'h28 == _match_key_qbytes_0_T_2 ? phv_data_40 : _GEN_47; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_49 = 8'h29 == _match_key_qbytes_0_T_2 ? phv_data_41 : _GEN_48; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_50 = 8'h2a == _match_key_qbytes_0_T_2 ? phv_data_42 : _GEN_49; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_51 = 8'h2b == _match_key_qbytes_0_T_2 ? phv_data_43 : _GEN_50; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_52 = 8'h2c == _match_key_qbytes_0_T_2 ? phv_data_44 : _GEN_51; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_53 = 8'h2d == _match_key_qbytes_0_T_2 ? phv_data_45 : _GEN_52; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_54 = 8'h2e == _match_key_qbytes_0_T_2 ? phv_data_46 : _GEN_53; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_55 = 8'h2f == _match_key_qbytes_0_T_2 ? phv_data_47 : _GEN_54; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_56 = 8'h30 == _match_key_qbytes_0_T_2 ? phv_data_48 : _GEN_55; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_57 = 8'h31 == _match_key_qbytes_0_T_2 ? phv_data_49 : _GEN_56; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_58 = 8'h32 == _match_key_qbytes_0_T_2 ? phv_data_50 : _GEN_57; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_59 = 8'h33 == _match_key_qbytes_0_T_2 ? phv_data_51 : _GEN_58; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_60 = 8'h34 == _match_key_qbytes_0_T_2 ? phv_data_52 : _GEN_59; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_61 = 8'h35 == _match_key_qbytes_0_T_2 ? phv_data_53 : _GEN_60; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_62 = 8'h36 == _match_key_qbytes_0_T_2 ? phv_data_54 : _GEN_61; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_63 = 8'h37 == _match_key_qbytes_0_T_2 ? phv_data_55 : _GEN_62; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_64 = 8'h38 == _match_key_qbytes_0_T_2 ? phv_data_56 : _GEN_63; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_65 = 8'h39 == _match_key_qbytes_0_T_2 ? phv_data_57 : _GEN_64; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_66 = 8'h3a == _match_key_qbytes_0_T_2 ? phv_data_58 : _GEN_65; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_67 = 8'h3b == _match_key_qbytes_0_T_2 ? phv_data_59 : _GEN_66; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_68 = 8'h3c == _match_key_qbytes_0_T_2 ? phv_data_60 : _GEN_67; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_69 = 8'h3d == _match_key_qbytes_0_T_2 ? phv_data_61 : _GEN_68; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_70 = 8'h3e == _match_key_qbytes_0_T_2 ? phv_data_62 : _GEN_69; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_71 = 8'h3f == _match_key_qbytes_0_T_2 ? phv_data_63 : _GEN_70; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_72 = 8'h40 == _match_key_qbytes_0_T_2 ? phv_data_64 : _GEN_71; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_73 = 8'h41 == _match_key_qbytes_0_T_2 ? phv_data_65 : _GEN_72; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_74 = 8'h42 == _match_key_qbytes_0_T_2 ? phv_data_66 : _GEN_73; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_75 = 8'h43 == _match_key_qbytes_0_T_2 ? phv_data_67 : _GEN_74; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_76 = 8'h44 == _match_key_qbytes_0_T_2 ? phv_data_68 : _GEN_75; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_77 = 8'h45 == _match_key_qbytes_0_T_2 ? phv_data_69 : _GEN_76; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_78 = 8'h46 == _match_key_qbytes_0_T_2 ? phv_data_70 : _GEN_77; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_79 = 8'h47 == _match_key_qbytes_0_T_2 ? phv_data_71 : _GEN_78; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_80 = 8'h48 == _match_key_qbytes_0_T_2 ? phv_data_72 : _GEN_79; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_81 = 8'h49 == _match_key_qbytes_0_T_2 ? phv_data_73 : _GEN_80; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_82 = 8'h4a == _match_key_qbytes_0_T_2 ? phv_data_74 : _GEN_81; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_83 = 8'h4b == _match_key_qbytes_0_T_2 ? phv_data_75 : _GEN_82; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_84 = 8'h4c == _match_key_qbytes_0_T_2 ? phv_data_76 : _GEN_83; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_85 = 8'h4d == _match_key_qbytes_0_T_2 ? phv_data_77 : _GEN_84; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_86 = 8'h4e == _match_key_qbytes_0_T_2 ? phv_data_78 : _GEN_85; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_87 = 8'h4f == _match_key_qbytes_0_T_2 ? phv_data_79 : _GEN_86; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_88 = 8'h50 == _match_key_qbytes_0_T_2 ? phv_data_80 : _GEN_87; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_89 = 8'h51 == _match_key_qbytes_0_T_2 ? phv_data_81 : _GEN_88; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_90 = 8'h52 == _match_key_qbytes_0_T_2 ? phv_data_82 : _GEN_89; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_91 = 8'h53 == _match_key_qbytes_0_T_2 ? phv_data_83 : _GEN_90; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_92 = 8'h54 == _match_key_qbytes_0_T_2 ? phv_data_84 : _GEN_91; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_93 = 8'h55 == _match_key_qbytes_0_T_2 ? phv_data_85 : _GEN_92; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_94 = 8'h56 == _match_key_qbytes_0_T_2 ? phv_data_86 : _GEN_93; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_95 = 8'h57 == _match_key_qbytes_0_T_2 ? phv_data_87 : _GEN_94; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_96 = 8'h58 == _match_key_qbytes_0_T_2 ? phv_data_88 : _GEN_95; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_97 = 8'h59 == _match_key_qbytes_0_T_2 ? phv_data_89 : _GEN_96; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_98 = 8'h5a == _match_key_qbytes_0_T_2 ? phv_data_90 : _GEN_97; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_99 = 8'h5b == _match_key_qbytes_0_T_2 ? phv_data_91 : _GEN_98; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_100 = 8'h5c == _match_key_qbytes_0_T_2 ? phv_data_92 : _GEN_99; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_101 = 8'h5d == _match_key_qbytes_0_T_2 ? phv_data_93 : _GEN_100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_102 = 8'h5e == _match_key_qbytes_0_T_2 ? phv_data_94 : _GEN_101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_103 = 8'h5f == _match_key_qbytes_0_T_2 ? phv_data_95 : _GEN_102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_104 = 8'h60 == _match_key_qbytes_0_T_2 ? phv_data_96 : _GEN_103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_105 = 8'h61 == _match_key_qbytes_0_T_2 ? phv_data_97 : _GEN_104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_106 = 8'h62 == _match_key_qbytes_0_T_2 ? phv_data_98 : _GEN_105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_107 = 8'h63 == _match_key_qbytes_0_T_2 ? phv_data_99 : _GEN_106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_108 = 8'h64 == _match_key_qbytes_0_T_2 ? phv_data_100 : _GEN_107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_109 = 8'h65 == _match_key_qbytes_0_T_2 ? phv_data_101 : _GEN_108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_110 = 8'h66 == _match_key_qbytes_0_T_2 ? phv_data_102 : _GEN_109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_111 = 8'h67 == _match_key_qbytes_0_T_2 ? phv_data_103 : _GEN_110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_112 = 8'h68 == _match_key_qbytes_0_T_2 ? phv_data_104 : _GEN_111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_113 = 8'h69 == _match_key_qbytes_0_T_2 ? phv_data_105 : _GEN_112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_114 = 8'h6a == _match_key_qbytes_0_T_2 ? phv_data_106 : _GEN_113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_115 = 8'h6b == _match_key_qbytes_0_T_2 ? phv_data_107 : _GEN_114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_116 = 8'h6c == _match_key_qbytes_0_T_2 ? phv_data_108 : _GEN_115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_117 = 8'h6d == _match_key_qbytes_0_T_2 ? phv_data_109 : _GEN_116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_118 = 8'h6e == _match_key_qbytes_0_T_2 ? phv_data_110 : _GEN_117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_119 = 8'h6f == _match_key_qbytes_0_T_2 ? phv_data_111 : _GEN_118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_120 = 8'h70 == _match_key_qbytes_0_T_2 ? phv_data_112 : _GEN_119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_121 = 8'h71 == _match_key_qbytes_0_T_2 ? phv_data_113 : _GEN_120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_122 = 8'h72 == _match_key_qbytes_0_T_2 ? phv_data_114 : _GEN_121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_123 = 8'h73 == _match_key_qbytes_0_T_2 ? phv_data_115 : _GEN_122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_124 = 8'h74 == _match_key_qbytes_0_T_2 ? phv_data_116 : _GEN_123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_125 = 8'h75 == _match_key_qbytes_0_T_2 ? phv_data_117 : _GEN_124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_126 = 8'h76 == _match_key_qbytes_0_T_2 ? phv_data_118 : _GEN_125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_127 = 8'h77 == _match_key_qbytes_0_T_2 ? phv_data_119 : _GEN_126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_128 = 8'h78 == _match_key_qbytes_0_T_2 ? phv_data_120 : _GEN_127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_129 = 8'h79 == _match_key_qbytes_0_T_2 ? phv_data_121 : _GEN_128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_130 = 8'h7a == _match_key_qbytes_0_T_2 ? phv_data_122 : _GEN_129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_131 = 8'h7b == _match_key_qbytes_0_T_2 ? phv_data_123 : _GEN_130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_132 = 8'h7c == _match_key_qbytes_0_T_2 ? phv_data_124 : _GEN_131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_133 = 8'h7d == _match_key_qbytes_0_T_2 ? phv_data_125 : _GEN_132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_134 = 8'h7e == _match_key_qbytes_0_T_2 ? phv_data_126 : _GEN_133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_135 = 8'h7f == _match_key_qbytes_0_T_2 ? phv_data_127 : _GEN_134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_136 = 8'h80 == _match_key_qbytes_0_T_2 ? phv_data_128 : _GEN_135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_137 = 8'h81 == _match_key_qbytes_0_T_2 ? phv_data_129 : _GEN_136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_138 = 8'h82 == _match_key_qbytes_0_T_2 ? phv_data_130 : _GEN_137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_139 = 8'h83 == _match_key_qbytes_0_T_2 ? phv_data_131 : _GEN_138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_140 = 8'h84 == _match_key_qbytes_0_T_2 ? phv_data_132 : _GEN_139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_141 = 8'h85 == _match_key_qbytes_0_T_2 ? phv_data_133 : _GEN_140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_142 = 8'h86 == _match_key_qbytes_0_T_2 ? phv_data_134 : _GEN_141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_143 = 8'h87 == _match_key_qbytes_0_T_2 ? phv_data_135 : _GEN_142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_144 = 8'h88 == _match_key_qbytes_0_T_2 ? phv_data_136 : _GEN_143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_145 = 8'h89 == _match_key_qbytes_0_T_2 ? phv_data_137 : _GEN_144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_146 = 8'h8a == _match_key_qbytes_0_T_2 ? phv_data_138 : _GEN_145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_147 = 8'h8b == _match_key_qbytes_0_T_2 ? phv_data_139 : _GEN_146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_148 = 8'h8c == _match_key_qbytes_0_T_2 ? phv_data_140 : _GEN_147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_149 = 8'h8d == _match_key_qbytes_0_T_2 ? phv_data_141 : _GEN_148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_150 = 8'h8e == _match_key_qbytes_0_T_2 ? phv_data_142 : _GEN_149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_151 = 8'h8f == _match_key_qbytes_0_T_2 ? phv_data_143 : _GEN_150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_152 = 8'h90 == _match_key_qbytes_0_T_2 ? phv_data_144 : _GEN_151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_153 = 8'h91 == _match_key_qbytes_0_T_2 ? phv_data_145 : _GEN_152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_154 = 8'h92 == _match_key_qbytes_0_T_2 ? phv_data_146 : _GEN_153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_155 = 8'h93 == _match_key_qbytes_0_T_2 ? phv_data_147 : _GEN_154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_156 = 8'h94 == _match_key_qbytes_0_T_2 ? phv_data_148 : _GEN_155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_157 = 8'h95 == _match_key_qbytes_0_T_2 ? phv_data_149 : _GEN_156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_158 = 8'h96 == _match_key_qbytes_0_T_2 ? phv_data_150 : _GEN_157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_159 = 8'h97 == _match_key_qbytes_0_T_2 ? phv_data_151 : _GEN_158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_160 = 8'h98 == _match_key_qbytes_0_T_2 ? phv_data_152 : _GEN_159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_161 = 8'h99 == _match_key_qbytes_0_T_2 ? phv_data_153 : _GEN_160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_162 = 8'h9a == _match_key_qbytes_0_T_2 ? phv_data_154 : _GEN_161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_163 = 8'h9b == _match_key_qbytes_0_T_2 ? phv_data_155 : _GEN_162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_164 = 8'h9c == _match_key_qbytes_0_T_2 ? phv_data_156 : _GEN_163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_165 = 8'h9d == _match_key_qbytes_0_T_2 ? phv_data_157 : _GEN_164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_166 = 8'h9e == _match_key_qbytes_0_T_2 ? phv_data_158 : _GEN_165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_167 = 8'h9f == _match_key_qbytes_0_T_2 ? phv_data_159 : _GEN_166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_169 = 8'h1 == local_offset ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_170 = 8'h2 == local_offset ? phv_data_2 : _GEN_169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_171 = 8'h3 == local_offset ? phv_data_3 : _GEN_170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_172 = 8'h4 == local_offset ? phv_data_4 : _GEN_171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_173 = 8'h5 == local_offset ? phv_data_5 : _GEN_172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_174 = 8'h6 == local_offset ? phv_data_6 : _GEN_173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_175 = 8'h7 == local_offset ? phv_data_7 : _GEN_174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_176 = 8'h8 == local_offset ? phv_data_8 : _GEN_175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_177 = 8'h9 == local_offset ? phv_data_9 : _GEN_176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_178 = 8'ha == local_offset ? phv_data_10 : _GEN_177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_179 = 8'hb == local_offset ? phv_data_11 : _GEN_178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_180 = 8'hc == local_offset ? phv_data_12 : _GEN_179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_181 = 8'hd == local_offset ? phv_data_13 : _GEN_180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_182 = 8'he == local_offset ? phv_data_14 : _GEN_181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_183 = 8'hf == local_offset ? phv_data_15 : _GEN_182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_184 = 8'h10 == local_offset ? phv_data_16 : _GEN_183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_185 = 8'h11 == local_offset ? phv_data_17 : _GEN_184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_186 = 8'h12 == local_offset ? phv_data_18 : _GEN_185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_187 = 8'h13 == local_offset ? phv_data_19 : _GEN_186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_188 = 8'h14 == local_offset ? phv_data_20 : _GEN_187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_189 = 8'h15 == local_offset ? phv_data_21 : _GEN_188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_190 = 8'h16 == local_offset ? phv_data_22 : _GEN_189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_191 = 8'h17 == local_offset ? phv_data_23 : _GEN_190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_192 = 8'h18 == local_offset ? phv_data_24 : _GEN_191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_193 = 8'h19 == local_offset ? phv_data_25 : _GEN_192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_194 = 8'h1a == local_offset ? phv_data_26 : _GEN_193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_195 = 8'h1b == local_offset ? phv_data_27 : _GEN_194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_196 = 8'h1c == local_offset ? phv_data_28 : _GEN_195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_197 = 8'h1d == local_offset ? phv_data_29 : _GEN_196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_198 = 8'h1e == local_offset ? phv_data_30 : _GEN_197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_199 = 8'h1f == local_offset ? phv_data_31 : _GEN_198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_200 = 8'h20 == local_offset ? phv_data_32 : _GEN_199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_201 = 8'h21 == local_offset ? phv_data_33 : _GEN_200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_202 = 8'h22 == local_offset ? phv_data_34 : _GEN_201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_203 = 8'h23 == local_offset ? phv_data_35 : _GEN_202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_204 = 8'h24 == local_offset ? phv_data_36 : _GEN_203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_205 = 8'h25 == local_offset ? phv_data_37 : _GEN_204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_206 = 8'h26 == local_offset ? phv_data_38 : _GEN_205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_207 = 8'h27 == local_offset ? phv_data_39 : _GEN_206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_208 = 8'h28 == local_offset ? phv_data_40 : _GEN_207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_209 = 8'h29 == local_offset ? phv_data_41 : _GEN_208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_210 = 8'h2a == local_offset ? phv_data_42 : _GEN_209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_211 = 8'h2b == local_offset ? phv_data_43 : _GEN_210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_212 = 8'h2c == local_offset ? phv_data_44 : _GEN_211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_213 = 8'h2d == local_offset ? phv_data_45 : _GEN_212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_214 = 8'h2e == local_offset ? phv_data_46 : _GEN_213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_215 = 8'h2f == local_offset ? phv_data_47 : _GEN_214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_216 = 8'h30 == local_offset ? phv_data_48 : _GEN_215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_217 = 8'h31 == local_offset ? phv_data_49 : _GEN_216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_218 = 8'h32 == local_offset ? phv_data_50 : _GEN_217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_219 = 8'h33 == local_offset ? phv_data_51 : _GEN_218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_220 = 8'h34 == local_offset ? phv_data_52 : _GEN_219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_221 = 8'h35 == local_offset ? phv_data_53 : _GEN_220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_222 = 8'h36 == local_offset ? phv_data_54 : _GEN_221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_223 = 8'h37 == local_offset ? phv_data_55 : _GEN_222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_224 = 8'h38 == local_offset ? phv_data_56 : _GEN_223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_225 = 8'h39 == local_offset ? phv_data_57 : _GEN_224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_226 = 8'h3a == local_offset ? phv_data_58 : _GEN_225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_227 = 8'h3b == local_offset ? phv_data_59 : _GEN_226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_228 = 8'h3c == local_offset ? phv_data_60 : _GEN_227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_229 = 8'h3d == local_offset ? phv_data_61 : _GEN_228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_230 = 8'h3e == local_offset ? phv_data_62 : _GEN_229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_231 = 8'h3f == local_offset ? phv_data_63 : _GEN_230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_232 = 8'h40 == local_offset ? phv_data_64 : _GEN_231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_233 = 8'h41 == local_offset ? phv_data_65 : _GEN_232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_234 = 8'h42 == local_offset ? phv_data_66 : _GEN_233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_235 = 8'h43 == local_offset ? phv_data_67 : _GEN_234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_236 = 8'h44 == local_offset ? phv_data_68 : _GEN_235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_237 = 8'h45 == local_offset ? phv_data_69 : _GEN_236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_238 = 8'h46 == local_offset ? phv_data_70 : _GEN_237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_239 = 8'h47 == local_offset ? phv_data_71 : _GEN_238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_240 = 8'h48 == local_offset ? phv_data_72 : _GEN_239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_241 = 8'h49 == local_offset ? phv_data_73 : _GEN_240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_242 = 8'h4a == local_offset ? phv_data_74 : _GEN_241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_243 = 8'h4b == local_offset ? phv_data_75 : _GEN_242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_244 = 8'h4c == local_offset ? phv_data_76 : _GEN_243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_245 = 8'h4d == local_offset ? phv_data_77 : _GEN_244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_246 = 8'h4e == local_offset ? phv_data_78 : _GEN_245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_247 = 8'h4f == local_offset ? phv_data_79 : _GEN_246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_248 = 8'h50 == local_offset ? phv_data_80 : _GEN_247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_249 = 8'h51 == local_offset ? phv_data_81 : _GEN_248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_250 = 8'h52 == local_offset ? phv_data_82 : _GEN_249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_251 = 8'h53 == local_offset ? phv_data_83 : _GEN_250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_252 = 8'h54 == local_offset ? phv_data_84 : _GEN_251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_253 = 8'h55 == local_offset ? phv_data_85 : _GEN_252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_254 = 8'h56 == local_offset ? phv_data_86 : _GEN_253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_255 = 8'h57 == local_offset ? phv_data_87 : _GEN_254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_256 = 8'h58 == local_offset ? phv_data_88 : _GEN_255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_257 = 8'h59 == local_offset ? phv_data_89 : _GEN_256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_258 = 8'h5a == local_offset ? phv_data_90 : _GEN_257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_259 = 8'h5b == local_offset ? phv_data_91 : _GEN_258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_260 = 8'h5c == local_offset ? phv_data_92 : _GEN_259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_261 = 8'h5d == local_offset ? phv_data_93 : _GEN_260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_262 = 8'h5e == local_offset ? phv_data_94 : _GEN_261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_263 = 8'h5f == local_offset ? phv_data_95 : _GEN_262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_264 = 8'h60 == local_offset ? phv_data_96 : _GEN_263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_265 = 8'h61 == local_offset ? phv_data_97 : _GEN_264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_266 = 8'h62 == local_offset ? phv_data_98 : _GEN_265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_267 = 8'h63 == local_offset ? phv_data_99 : _GEN_266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_268 = 8'h64 == local_offset ? phv_data_100 : _GEN_267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_269 = 8'h65 == local_offset ? phv_data_101 : _GEN_268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_270 = 8'h66 == local_offset ? phv_data_102 : _GEN_269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_271 = 8'h67 == local_offset ? phv_data_103 : _GEN_270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_272 = 8'h68 == local_offset ? phv_data_104 : _GEN_271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_273 = 8'h69 == local_offset ? phv_data_105 : _GEN_272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_274 = 8'h6a == local_offset ? phv_data_106 : _GEN_273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_275 = 8'h6b == local_offset ? phv_data_107 : _GEN_274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_276 = 8'h6c == local_offset ? phv_data_108 : _GEN_275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_277 = 8'h6d == local_offset ? phv_data_109 : _GEN_276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_278 = 8'h6e == local_offset ? phv_data_110 : _GEN_277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_279 = 8'h6f == local_offset ? phv_data_111 : _GEN_278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_280 = 8'h70 == local_offset ? phv_data_112 : _GEN_279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_281 = 8'h71 == local_offset ? phv_data_113 : _GEN_280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_282 = 8'h72 == local_offset ? phv_data_114 : _GEN_281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_283 = 8'h73 == local_offset ? phv_data_115 : _GEN_282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_284 = 8'h74 == local_offset ? phv_data_116 : _GEN_283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_285 = 8'h75 == local_offset ? phv_data_117 : _GEN_284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_286 = 8'h76 == local_offset ? phv_data_118 : _GEN_285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_287 = 8'h77 == local_offset ? phv_data_119 : _GEN_286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_288 = 8'h78 == local_offset ? phv_data_120 : _GEN_287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_289 = 8'h79 == local_offset ? phv_data_121 : _GEN_288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_290 = 8'h7a == local_offset ? phv_data_122 : _GEN_289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_291 = 8'h7b == local_offset ? phv_data_123 : _GEN_290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_292 = 8'h7c == local_offset ? phv_data_124 : _GEN_291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_293 = 8'h7d == local_offset ? phv_data_125 : _GEN_292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_294 = 8'h7e == local_offset ? phv_data_126 : _GEN_293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_295 = 8'h7f == local_offset ? phv_data_127 : _GEN_294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_296 = 8'h80 == local_offset ? phv_data_128 : _GEN_295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_297 = 8'h81 == local_offset ? phv_data_129 : _GEN_296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_298 = 8'h82 == local_offset ? phv_data_130 : _GEN_297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_299 = 8'h83 == local_offset ? phv_data_131 : _GEN_298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_300 = 8'h84 == local_offset ? phv_data_132 : _GEN_299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_301 = 8'h85 == local_offset ? phv_data_133 : _GEN_300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_302 = 8'h86 == local_offset ? phv_data_134 : _GEN_301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_303 = 8'h87 == local_offset ? phv_data_135 : _GEN_302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_304 = 8'h88 == local_offset ? phv_data_136 : _GEN_303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_305 = 8'h89 == local_offset ? phv_data_137 : _GEN_304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_306 = 8'h8a == local_offset ? phv_data_138 : _GEN_305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_307 = 8'h8b == local_offset ? phv_data_139 : _GEN_306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_308 = 8'h8c == local_offset ? phv_data_140 : _GEN_307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_309 = 8'h8d == local_offset ? phv_data_141 : _GEN_308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_310 = 8'h8e == local_offset ? phv_data_142 : _GEN_309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_311 = 8'h8f == local_offset ? phv_data_143 : _GEN_310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_312 = 8'h90 == local_offset ? phv_data_144 : _GEN_311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_313 = 8'h91 == local_offset ? phv_data_145 : _GEN_312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_314 = 8'h92 == local_offset ? phv_data_146 : _GEN_313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_315 = 8'h93 == local_offset ? phv_data_147 : _GEN_314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_316 = 8'h94 == local_offset ? phv_data_148 : _GEN_315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_317 = 8'h95 == local_offset ? phv_data_149 : _GEN_316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_318 = 8'h96 == local_offset ? phv_data_150 : _GEN_317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_319 = 8'h97 == local_offset ? phv_data_151 : _GEN_318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_320 = 8'h98 == local_offset ? phv_data_152 : _GEN_319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_321 = 8'h99 == local_offset ? phv_data_153 : _GEN_320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_322 = 8'h9a == local_offset ? phv_data_154 : _GEN_321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_323 = 8'h9b == local_offset ? phv_data_155 : _GEN_322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_324 = 8'h9c == local_offset ? phv_data_156 : _GEN_323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_325 = 8'h9d == local_offset ? phv_data_157 : _GEN_324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_326 = 8'h9e == local_offset ? phv_data_158 : _GEN_325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_327 = 8'h9f == local_offset ? phv_data_159 : _GEN_326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_329 = 8'h1 == _match_key_qbytes_0_T ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_330 = 8'h2 == _match_key_qbytes_0_T ? phv_data_2 : _GEN_329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_331 = 8'h3 == _match_key_qbytes_0_T ? phv_data_3 : _GEN_330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_332 = 8'h4 == _match_key_qbytes_0_T ? phv_data_4 : _GEN_331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_333 = 8'h5 == _match_key_qbytes_0_T ? phv_data_5 : _GEN_332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_334 = 8'h6 == _match_key_qbytes_0_T ? phv_data_6 : _GEN_333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_335 = 8'h7 == _match_key_qbytes_0_T ? phv_data_7 : _GEN_334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_336 = 8'h8 == _match_key_qbytes_0_T ? phv_data_8 : _GEN_335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_337 = 8'h9 == _match_key_qbytes_0_T ? phv_data_9 : _GEN_336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_338 = 8'ha == _match_key_qbytes_0_T ? phv_data_10 : _GEN_337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_339 = 8'hb == _match_key_qbytes_0_T ? phv_data_11 : _GEN_338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_340 = 8'hc == _match_key_qbytes_0_T ? phv_data_12 : _GEN_339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_341 = 8'hd == _match_key_qbytes_0_T ? phv_data_13 : _GEN_340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_342 = 8'he == _match_key_qbytes_0_T ? phv_data_14 : _GEN_341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_343 = 8'hf == _match_key_qbytes_0_T ? phv_data_15 : _GEN_342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_344 = 8'h10 == _match_key_qbytes_0_T ? phv_data_16 : _GEN_343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_345 = 8'h11 == _match_key_qbytes_0_T ? phv_data_17 : _GEN_344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_346 = 8'h12 == _match_key_qbytes_0_T ? phv_data_18 : _GEN_345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_347 = 8'h13 == _match_key_qbytes_0_T ? phv_data_19 : _GEN_346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_348 = 8'h14 == _match_key_qbytes_0_T ? phv_data_20 : _GEN_347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_349 = 8'h15 == _match_key_qbytes_0_T ? phv_data_21 : _GEN_348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_350 = 8'h16 == _match_key_qbytes_0_T ? phv_data_22 : _GEN_349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_351 = 8'h17 == _match_key_qbytes_0_T ? phv_data_23 : _GEN_350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_352 = 8'h18 == _match_key_qbytes_0_T ? phv_data_24 : _GEN_351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_353 = 8'h19 == _match_key_qbytes_0_T ? phv_data_25 : _GEN_352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_354 = 8'h1a == _match_key_qbytes_0_T ? phv_data_26 : _GEN_353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_355 = 8'h1b == _match_key_qbytes_0_T ? phv_data_27 : _GEN_354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_356 = 8'h1c == _match_key_qbytes_0_T ? phv_data_28 : _GEN_355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_357 = 8'h1d == _match_key_qbytes_0_T ? phv_data_29 : _GEN_356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_358 = 8'h1e == _match_key_qbytes_0_T ? phv_data_30 : _GEN_357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_359 = 8'h1f == _match_key_qbytes_0_T ? phv_data_31 : _GEN_358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_360 = 8'h20 == _match_key_qbytes_0_T ? phv_data_32 : _GEN_359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_361 = 8'h21 == _match_key_qbytes_0_T ? phv_data_33 : _GEN_360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_362 = 8'h22 == _match_key_qbytes_0_T ? phv_data_34 : _GEN_361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_363 = 8'h23 == _match_key_qbytes_0_T ? phv_data_35 : _GEN_362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_364 = 8'h24 == _match_key_qbytes_0_T ? phv_data_36 : _GEN_363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_365 = 8'h25 == _match_key_qbytes_0_T ? phv_data_37 : _GEN_364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_366 = 8'h26 == _match_key_qbytes_0_T ? phv_data_38 : _GEN_365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_367 = 8'h27 == _match_key_qbytes_0_T ? phv_data_39 : _GEN_366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_368 = 8'h28 == _match_key_qbytes_0_T ? phv_data_40 : _GEN_367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_369 = 8'h29 == _match_key_qbytes_0_T ? phv_data_41 : _GEN_368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_370 = 8'h2a == _match_key_qbytes_0_T ? phv_data_42 : _GEN_369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_371 = 8'h2b == _match_key_qbytes_0_T ? phv_data_43 : _GEN_370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_372 = 8'h2c == _match_key_qbytes_0_T ? phv_data_44 : _GEN_371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_373 = 8'h2d == _match_key_qbytes_0_T ? phv_data_45 : _GEN_372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_374 = 8'h2e == _match_key_qbytes_0_T ? phv_data_46 : _GEN_373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_375 = 8'h2f == _match_key_qbytes_0_T ? phv_data_47 : _GEN_374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_376 = 8'h30 == _match_key_qbytes_0_T ? phv_data_48 : _GEN_375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_377 = 8'h31 == _match_key_qbytes_0_T ? phv_data_49 : _GEN_376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_378 = 8'h32 == _match_key_qbytes_0_T ? phv_data_50 : _GEN_377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_379 = 8'h33 == _match_key_qbytes_0_T ? phv_data_51 : _GEN_378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_380 = 8'h34 == _match_key_qbytes_0_T ? phv_data_52 : _GEN_379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_381 = 8'h35 == _match_key_qbytes_0_T ? phv_data_53 : _GEN_380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_382 = 8'h36 == _match_key_qbytes_0_T ? phv_data_54 : _GEN_381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_383 = 8'h37 == _match_key_qbytes_0_T ? phv_data_55 : _GEN_382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_384 = 8'h38 == _match_key_qbytes_0_T ? phv_data_56 : _GEN_383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_385 = 8'h39 == _match_key_qbytes_0_T ? phv_data_57 : _GEN_384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_386 = 8'h3a == _match_key_qbytes_0_T ? phv_data_58 : _GEN_385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_387 = 8'h3b == _match_key_qbytes_0_T ? phv_data_59 : _GEN_386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_388 = 8'h3c == _match_key_qbytes_0_T ? phv_data_60 : _GEN_387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_389 = 8'h3d == _match_key_qbytes_0_T ? phv_data_61 : _GEN_388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_390 = 8'h3e == _match_key_qbytes_0_T ? phv_data_62 : _GEN_389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_391 = 8'h3f == _match_key_qbytes_0_T ? phv_data_63 : _GEN_390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_392 = 8'h40 == _match_key_qbytes_0_T ? phv_data_64 : _GEN_391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_393 = 8'h41 == _match_key_qbytes_0_T ? phv_data_65 : _GEN_392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_394 = 8'h42 == _match_key_qbytes_0_T ? phv_data_66 : _GEN_393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_395 = 8'h43 == _match_key_qbytes_0_T ? phv_data_67 : _GEN_394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_396 = 8'h44 == _match_key_qbytes_0_T ? phv_data_68 : _GEN_395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_397 = 8'h45 == _match_key_qbytes_0_T ? phv_data_69 : _GEN_396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_398 = 8'h46 == _match_key_qbytes_0_T ? phv_data_70 : _GEN_397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_399 = 8'h47 == _match_key_qbytes_0_T ? phv_data_71 : _GEN_398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_400 = 8'h48 == _match_key_qbytes_0_T ? phv_data_72 : _GEN_399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_401 = 8'h49 == _match_key_qbytes_0_T ? phv_data_73 : _GEN_400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_402 = 8'h4a == _match_key_qbytes_0_T ? phv_data_74 : _GEN_401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_403 = 8'h4b == _match_key_qbytes_0_T ? phv_data_75 : _GEN_402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_404 = 8'h4c == _match_key_qbytes_0_T ? phv_data_76 : _GEN_403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_405 = 8'h4d == _match_key_qbytes_0_T ? phv_data_77 : _GEN_404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_406 = 8'h4e == _match_key_qbytes_0_T ? phv_data_78 : _GEN_405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_407 = 8'h4f == _match_key_qbytes_0_T ? phv_data_79 : _GEN_406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_408 = 8'h50 == _match_key_qbytes_0_T ? phv_data_80 : _GEN_407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_409 = 8'h51 == _match_key_qbytes_0_T ? phv_data_81 : _GEN_408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_410 = 8'h52 == _match_key_qbytes_0_T ? phv_data_82 : _GEN_409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_411 = 8'h53 == _match_key_qbytes_0_T ? phv_data_83 : _GEN_410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_412 = 8'h54 == _match_key_qbytes_0_T ? phv_data_84 : _GEN_411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_413 = 8'h55 == _match_key_qbytes_0_T ? phv_data_85 : _GEN_412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_414 = 8'h56 == _match_key_qbytes_0_T ? phv_data_86 : _GEN_413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_415 = 8'h57 == _match_key_qbytes_0_T ? phv_data_87 : _GEN_414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_416 = 8'h58 == _match_key_qbytes_0_T ? phv_data_88 : _GEN_415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_417 = 8'h59 == _match_key_qbytes_0_T ? phv_data_89 : _GEN_416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_418 = 8'h5a == _match_key_qbytes_0_T ? phv_data_90 : _GEN_417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_419 = 8'h5b == _match_key_qbytes_0_T ? phv_data_91 : _GEN_418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_420 = 8'h5c == _match_key_qbytes_0_T ? phv_data_92 : _GEN_419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_421 = 8'h5d == _match_key_qbytes_0_T ? phv_data_93 : _GEN_420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_422 = 8'h5e == _match_key_qbytes_0_T ? phv_data_94 : _GEN_421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_423 = 8'h5f == _match_key_qbytes_0_T ? phv_data_95 : _GEN_422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_424 = 8'h60 == _match_key_qbytes_0_T ? phv_data_96 : _GEN_423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_425 = 8'h61 == _match_key_qbytes_0_T ? phv_data_97 : _GEN_424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_426 = 8'h62 == _match_key_qbytes_0_T ? phv_data_98 : _GEN_425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_427 = 8'h63 == _match_key_qbytes_0_T ? phv_data_99 : _GEN_426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_428 = 8'h64 == _match_key_qbytes_0_T ? phv_data_100 : _GEN_427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_429 = 8'h65 == _match_key_qbytes_0_T ? phv_data_101 : _GEN_428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_430 = 8'h66 == _match_key_qbytes_0_T ? phv_data_102 : _GEN_429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_431 = 8'h67 == _match_key_qbytes_0_T ? phv_data_103 : _GEN_430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_432 = 8'h68 == _match_key_qbytes_0_T ? phv_data_104 : _GEN_431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_433 = 8'h69 == _match_key_qbytes_0_T ? phv_data_105 : _GEN_432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_434 = 8'h6a == _match_key_qbytes_0_T ? phv_data_106 : _GEN_433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_435 = 8'h6b == _match_key_qbytes_0_T ? phv_data_107 : _GEN_434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_436 = 8'h6c == _match_key_qbytes_0_T ? phv_data_108 : _GEN_435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_437 = 8'h6d == _match_key_qbytes_0_T ? phv_data_109 : _GEN_436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_438 = 8'h6e == _match_key_qbytes_0_T ? phv_data_110 : _GEN_437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_439 = 8'h6f == _match_key_qbytes_0_T ? phv_data_111 : _GEN_438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_440 = 8'h70 == _match_key_qbytes_0_T ? phv_data_112 : _GEN_439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_441 = 8'h71 == _match_key_qbytes_0_T ? phv_data_113 : _GEN_440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_442 = 8'h72 == _match_key_qbytes_0_T ? phv_data_114 : _GEN_441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_443 = 8'h73 == _match_key_qbytes_0_T ? phv_data_115 : _GEN_442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_444 = 8'h74 == _match_key_qbytes_0_T ? phv_data_116 : _GEN_443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_445 = 8'h75 == _match_key_qbytes_0_T ? phv_data_117 : _GEN_444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_446 = 8'h76 == _match_key_qbytes_0_T ? phv_data_118 : _GEN_445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_447 = 8'h77 == _match_key_qbytes_0_T ? phv_data_119 : _GEN_446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_448 = 8'h78 == _match_key_qbytes_0_T ? phv_data_120 : _GEN_447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_449 = 8'h79 == _match_key_qbytes_0_T ? phv_data_121 : _GEN_448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_450 = 8'h7a == _match_key_qbytes_0_T ? phv_data_122 : _GEN_449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_451 = 8'h7b == _match_key_qbytes_0_T ? phv_data_123 : _GEN_450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_452 = 8'h7c == _match_key_qbytes_0_T ? phv_data_124 : _GEN_451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_453 = 8'h7d == _match_key_qbytes_0_T ? phv_data_125 : _GEN_452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_454 = 8'h7e == _match_key_qbytes_0_T ? phv_data_126 : _GEN_453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_455 = 8'h7f == _match_key_qbytes_0_T ? phv_data_127 : _GEN_454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_456 = 8'h80 == _match_key_qbytes_0_T ? phv_data_128 : _GEN_455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_457 = 8'h81 == _match_key_qbytes_0_T ? phv_data_129 : _GEN_456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_458 = 8'h82 == _match_key_qbytes_0_T ? phv_data_130 : _GEN_457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_459 = 8'h83 == _match_key_qbytes_0_T ? phv_data_131 : _GEN_458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_460 = 8'h84 == _match_key_qbytes_0_T ? phv_data_132 : _GEN_459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_461 = 8'h85 == _match_key_qbytes_0_T ? phv_data_133 : _GEN_460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_462 = 8'h86 == _match_key_qbytes_0_T ? phv_data_134 : _GEN_461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_463 = 8'h87 == _match_key_qbytes_0_T ? phv_data_135 : _GEN_462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_464 = 8'h88 == _match_key_qbytes_0_T ? phv_data_136 : _GEN_463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_465 = 8'h89 == _match_key_qbytes_0_T ? phv_data_137 : _GEN_464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_466 = 8'h8a == _match_key_qbytes_0_T ? phv_data_138 : _GEN_465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_467 = 8'h8b == _match_key_qbytes_0_T ? phv_data_139 : _GEN_466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_468 = 8'h8c == _match_key_qbytes_0_T ? phv_data_140 : _GEN_467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_469 = 8'h8d == _match_key_qbytes_0_T ? phv_data_141 : _GEN_468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_470 = 8'h8e == _match_key_qbytes_0_T ? phv_data_142 : _GEN_469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_471 = 8'h8f == _match_key_qbytes_0_T ? phv_data_143 : _GEN_470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_472 = 8'h90 == _match_key_qbytes_0_T ? phv_data_144 : _GEN_471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_473 = 8'h91 == _match_key_qbytes_0_T ? phv_data_145 : _GEN_472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_474 = 8'h92 == _match_key_qbytes_0_T ? phv_data_146 : _GEN_473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_475 = 8'h93 == _match_key_qbytes_0_T ? phv_data_147 : _GEN_474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_476 = 8'h94 == _match_key_qbytes_0_T ? phv_data_148 : _GEN_475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_477 = 8'h95 == _match_key_qbytes_0_T ? phv_data_149 : _GEN_476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_478 = 8'h96 == _match_key_qbytes_0_T ? phv_data_150 : _GEN_477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_479 = 8'h97 == _match_key_qbytes_0_T ? phv_data_151 : _GEN_478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_480 = 8'h98 == _match_key_qbytes_0_T ? phv_data_152 : _GEN_479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_481 = 8'h99 == _match_key_qbytes_0_T ? phv_data_153 : _GEN_480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_482 = 8'h9a == _match_key_qbytes_0_T ? phv_data_154 : _GEN_481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_483 = 8'h9b == _match_key_qbytes_0_T ? phv_data_155 : _GEN_482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_484 = 8'h9c == _match_key_qbytes_0_T ? phv_data_156 : _GEN_483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_485 = 8'h9d == _match_key_qbytes_0_T ? phv_data_157 : _GEN_484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_486 = 8'h9e == _match_key_qbytes_0_T ? phv_data_158 : _GEN_485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_487 = 8'h9f == _match_key_qbytes_0_T ? phv_data_159 : _GEN_486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_489 = 8'h1 == _match_key_qbytes_0_T_1 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_490 = 8'h2 == _match_key_qbytes_0_T_1 ? phv_data_2 : _GEN_489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_491 = 8'h3 == _match_key_qbytes_0_T_1 ? phv_data_3 : _GEN_490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_492 = 8'h4 == _match_key_qbytes_0_T_1 ? phv_data_4 : _GEN_491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_493 = 8'h5 == _match_key_qbytes_0_T_1 ? phv_data_5 : _GEN_492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_494 = 8'h6 == _match_key_qbytes_0_T_1 ? phv_data_6 : _GEN_493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_495 = 8'h7 == _match_key_qbytes_0_T_1 ? phv_data_7 : _GEN_494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_496 = 8'h8 == _match_key_qbytes_0_T_1 ? phv_data_8 : _GEN_495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_497 = 8'h9 == _match_key_qbytes_0_T_1 ? phv_data_9 : _GEN_496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_498 = 8'ha == _match_key_qbytes_0_T_1 ? phv_data_10 : _GEN_497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_499 = 8'hb == _match_key_qbytes_0_T_1 ? phv_data_11 : _GEN_498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_500 = 8'hc == _match_key_qbytes_0_T_1 ? phv_data_12 : _GEN_499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_501 = 8'hd == _match_key_qbytes_0_T_1 ? phv_data_13 : _GEN_500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_502 = 8'he == _match_key_qbytes_0_T_1 ? phv_data_14 : _GEN_501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_503 = 8'hf == _match_key_qbytes_0_T_1 ? phv_data_15 : _GEN_502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_504 = 8'h10 == _match_key_qbytes_0_T_1 ? phv_data_16 : _GEN_503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_505 = 8'h11 == _match_key_qbytes_0_T_1 ? phv_data_17 : _GEN_504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_506 = 8'h12 == _match_key_qbytes_0_T_1 ? phv_data_18 : _GEN_505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_507 = 8'h13 == _match_key_qbytes_0_T_1 ? phv_data_19 : _GEN_506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_508 = 8'h14 == _match_key_qbytes_0_T_1 ? phv_data_20 : _GEN_507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_509 = 8'h15 == _match_key_qbytes_0_T_1 ? phv_data_21 : _GEN_508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_510 = 8'h16 == _match_key_qbytes_0_T_1 ? phv_data_22 : _GEN_509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_511 = 8'h17 == _match_key_qbytes_0_T_1 ? phv_data_23 : _GEN_510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_512 = 8'h18 == _match_key_qbytes_0_T_1 ? phv_data_24 : _GEN_511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_513 = 8'h19 == _match_key_qbytes_0_T_1 ? phv_data_25 : _GEN_512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_514 = 8'h1a == _match_key_qbytes_0_T_1 ? phv_data_26 : _GEN_513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_515 = 8'h1b == _match_key_qbytes_0_T_1 ? phv_data_27 : _GEN_514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_516 = 8'h1c == _match_key_qbytes_0_T_1 ? phv_data_28 : _GEN_515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_517 = 8'h1d == _match_key_qbytes_0_T_1 ? phv_data_29 : _GEN_516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_518 = 8'h1e == _match_key_qbytes_0_T_1 ? phv_data_30 : _GEN_517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_519 = 8'h1f == _match_key_qbytes_0_T_1 ? phv_data_31 : _GEN_518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_520 = 8'h20 == _match_key_qbytes_0_T_1 ? phv_data_32 : _GEN_519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_521 = 8'h21 == _match_key_qbytes_0_T_1 ? phv_data_33 : _GEN_520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_522 = 8'h22 == _match_key_qbytes_0_T_1 ? phv_data_34 : _GEN_521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_523 = 8'h23 == _match_key_qbytes_0_T_1 ? phv_data_35 : _GEN_522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_524 = 8'h24 == _match_key_qbytes_0_T_1 ? phv_data_36 : _GEN_523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_525 = 8'h25 == _match_key_qbytes_0_T_1 ? phv_data_37 : _GEN_524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_526 = 8'h26 == _match_key_qbytes_0_T_1 ? phv_data_38 : _GEN_525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_527 = 8'h27 == _match_key_qbytes_0_T_1 ? phv_data_39 : _GEN_526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_528 = 8'h28 == _match_key_qbytes_0_T_1 ? phv_data_40 : _GEN_527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_529 = 8'h29 == _match_key_qbytes_0_T_1 ? phv_data_41 : _GEN_528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_530 = 8'h2a == _match_key_qbytes_0_T_1 ? phv_data_42 : _GEN_529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_531 = 8'h2b == _match_key_qbytes_0_T_1 ? phv_data_43 : _GEN_530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_532 = 8'h2c == _match_key_qbytes_0_T_1 ? phv_data_44 : _GEN_531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_533 = 8'h2d == _match_key_qbytes_0_T_1 ? phv_data_45 : _GEN_532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_534 = 8'h2e == _match_key_qbytes_0_T_1 ? phv_data_46 : _GEN_533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_535 = 8'h2f == _match_key_qbytes_0_T_1 ? phv_data_47 : _GEN_534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_536 = 8'h30 == _match_key_qbytes_0_T_1 ? phv_data_48 : _GEN_535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_537 = 8'h31 == _match_key_qbytes_0_T_1 ? phv_data_49 : _GEN_536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_538 = 8'h32 == _match_key_qbytes_0_T_1 ? phv_data_50 : _GEN_537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_539 = 8'h33 == _match_key_qbytes_0_T_1 ? phv_data_51 : _GEN_538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_540 = 8'h34 == _match_key_qbytes_0_T_1 ? phv_data_52 : _GEN_539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_541 = 8'h35 == _match_key_qbytes_0_T_1 ? phv_data_53 : _GEN_540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_542 = 8'h36 == _match_key_qbytes_0_T_1 ? phv_data_54 : _GEN_541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_543 = 8'h37 == _match_key_qbytes_0_T_1 ? phv_data_55 : _GEN_542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_544 = 8'h38 == _match_key_qbytes_0_T_1 ? phv_data_56 : _GEN_543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_545 = 8'h39 == _match_key_qbytes_0_T_1 ? phv_data_57 : _GEN_544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_546 = 8'h3a == _match_key_qbytes_0_T_1 ? phv_data_58 : _GEN_545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_547 = 8'h3b == _match_key_qbytes_0_T_1 ? phv_data_59 : _GEN_546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_548 = 8'h3c == _match_key_qbytes_0_T_1 ? phv_data_60 : _GEN_547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_549 = 8'h3d == _match_key_qbytes_0_T_1 ? phv_data_61 : _GEN_548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_550 = 8'h3e == _match_key_qbytes_0_T_1 ? phv_data_62 : _GEN_549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_551 = 8'h3f == _match_key_qbytes_0_T_1 ? phv_data_63 : _GEN_550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_552 = 8'h40 == _match_key_qbytes_0_T_1 ? phv_data_64 : _GEN_551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_553 = 8'h41 == _match_key_qbytes_0_T_1 ? phv_data_65 : _GEN_552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_554 = 8'h42 == _match_key_qbytes_0_T_1 ? phv_data_66 : _GEN_553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_555 = 8'h43 == _match_key_qbytes_0_T_1 ? phv_data_67 : _GEN_554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_556 = 8'h44 == _match_key_qbytes_0_T_1 ? phv_data_68 : _GEN_555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_557 = 8'h45 == _match_key_qbytes_0_T_1 ? phv_data_69 : _GEN_556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_558 = 8'h46 == _match_key_qbytes_0_T_1 ? phv_data_70 : _GEN_557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_559 = 8'h47 == _match_key_qbytes_0_T_1 ? phv_data_71 : _GEN_558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_560 = 8'h48 == _match_key_qbytes_0_T_1 ? phv_data_72 : _GEN_559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_561 = 8'h49 == _match_key_qbytes_0_T_1 ? phv_data_73 : _GEN_560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_562 = 8'h4a == _match_key_qbytes_0_T_1 ? phv_data_74 : _GEN_561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_563 = 8'h4b == _match_key_qbytes_0_T_1 ? phv_data_75 : _GEN_562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_564 = 8'h4c == _match_key_qbytes_0_T_1 ? phv_data_76 : _GEN_563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_565 = 8'h4d == _match_key_qbytes_0_T_1 ? phv_data_77 : _GEN_564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_566 = 8'h4e == _match_key_qbytes_0_T_1 ? phv_data_78 : _GEN_565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_567 = 8'h4f == _match_key_qbytes_0_T_1 ? phv_data_79 : _GEN_566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_568 = 8'h50 == _match_key_qbytes_0_T_1 ? phv_data_80 : _GEN_567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_569 = 8'h51 == _match_key_qbytes_0_T_1 ? phv_data_81 : _GEN_568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_570 = 8'h52 == _match_key_qbytes_0_T_1 ? phv_data_82 : _GEN_569; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_571 = 8'h53 == _match_key_qbytes_0_T_1 ? phv_data_83 : _GEN_570; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_572 = 8'h54 == _match_key_qbytes_0_T_1 ? phv_data_84 : _GEN_571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_573 = 8'h55 == _match_key_qbytes_0_T_1 ? phv_data_85 : _GEN_572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_574 = 8'h56 == _match_key_qbytes_0_T_1 ? phv_data_86 : _GEN_573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_575 = 8'h57 == _match_key_qbytes_0_T_1 ? phv_data_87 : _GEN_574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_576 = 8'h58 == _match_key_qbytes_0_T_1 ? phv_data_88 : _GEN_575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_577 = 8'h59 == _match_key_qbytes_0_T_1 ? phv_data_89 : _GEN_576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_578 = 8'h5a == _match_key_qbytes_0_T_1 ? phv_data_90 : _GEN_577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_579 = 8'h5b == _match_key_qbytes_0_T_1 ? phv_data_91 : _GEN_578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_580 = 8'h5c == _match_key_qbytes_0_T_1 ? phv_data_92 : _GEN_579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_581 = 8'h5d == _match_key_qbytes_0_T_1 ? phv_data_93 : _GEN_580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_582 = 8'h5e == _match_key_qbytes_0_T_1 ? phv_data_94 : _GEN_581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_583 = 8'h5f == _match_key_qbytes_0_T_1 ? phv_data_95 : _GEN_582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_584 = 8'h60 == _match_key_qbytes_0_T_1 ? phv_data_96 : _GEN_583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_585 = 8'h61 == _match_key_qbytes_0_T_1 ? phv_data_97 : _GEN_584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_586 = 8'h62 == _match_key_qbytes_0_T_1 ? phv_data_98 : _GEN_585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_587 = 8'h63 == _match_key_qbytes_0_T_1 ? phv_data_99 : _GEN_586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_588 = 8'h64 == _match_key_qbytes_0_T_1 ? phv_data_100 : _GEN_587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_589 = 8'h65 == _match_key_qbytes_0_T_1 ? phv_data_101 : _GEN_588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_590 = 8'h66 == _match_key_qbytes_0_T_1 ? phv_data_102 : _GEN_589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_591 = 8'h67 == _match_key_qbytes_0_T_1 ? phv_data_103 : _GEN_590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_592 = 8'h68 == _match_key_qbytes_0_T_1 ? phv_data_104 : _GEN_591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_593 = 8'h69 == _match_key_qbytes_0_T_1 ? phv_data_105 : _GEN_592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_594 = 8'h6a == _match_key_qbytes_0_T_1 ? phv_data_106 : _GEN_593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_595 = 8'h6b == _match_key_qbytes_0_T_1 ? phv_data_107 : _GEN_594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_596 = 8'h6c == _match_key_qbytes_0_T_1 ? phv_data_108 : _GEN_595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_597 = 8'h6d == _match_key_qbytes_0_T_1 ? phv_data_109 : _GEN_596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_598 = 8'h6e == _match_key_qbytes_0_T_1 ? phv_data_110 : _GEN_597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_599 = 8'h6f == _match_key_qbytes_0_T_1 ? phv_data_111 : _GEN_598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_600 = 8'h70 == _match_key_qbytes_0_T_1 ? phv_data_112 : _GEN_599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_601 = 8'h71 == _match_key_qbytes_0_T_1 ? phv_data_113 : _GEN_600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_602 = 8'h72 == _match_key_qbytes_0_T_1 ? phv_data_114 : _GEN_601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_603 = 8'h73 == _match_key_qbytes_0_T_1 ? phv_data_115 : _GEN_602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_604 = 8'h74 == _match_key_qbytes_0_T_1 ? phv_data_116 : _GEN_603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_605 = 8'h75 == _match_key_qbytes_0_T_1 ? phv_data_117 : _GEN_604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_606 = 8'h76 == _match_key_qbytes_0_T_1 ? phv_data_118 : _GEN_605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_607 = 8'h77 == _match_key_qbytes_0_T_1 ? phv_data_119 : _GEN_606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_608 = 8'h78 == _match_key_qbytes_0_T_1 ? phv_data_120 : _GEN_607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_609 = 8'h79 == _match_key_qbytes_0_T_1 ? phv_data_121 : _GEN_608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_610 = 8'h7a == _match_key_qbytes_0_T_1 ? phv_data_122 : _GEN_609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_611 = 8'h7b == _match_key_qbytes_0_T_1 ? phv_data_123 : _GEN_610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_612 = 8'h7c == _match_key_qbytes_0_T_1 ? phv_data_124 : _GEN_611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_613 = 8'h7d == _match_key_qbytes_0_T_1 ? phv_data_125 : _GEN_612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_614 = 8'h7e == _match_key_qbytes_0_T_1 ? phv_data_126 : _GEN_613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_615 = 8'h7f == _match_key_qbytes_0_T_1 ? phv_data_127 : _GEN_614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_616 = 8'h80 == _match_key_qbytes_0_T_1 ? phv_data_128 : _GEN_615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_617 = 8'h81 == _match_key_qbytes_0_T_1 ? phv_data_129 : _GEN_616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_618 = 8'h82 == _match_key_qbytes_0_T_1 ? phv_data_130 : _GEN_617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_619 = 8'h83 == _match_key_qbytes_0_T_1 ? phv_data_131 : _GEN_618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_620 = 8'h84 == _match_key_qbytes_0_T_1 ? phv_data_132 : _GEN_619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_621 = 8'h85 == _match_key_qbytes_0_T_1 ? phv_data_133 : _GEN_620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_622 = 8'h86 == _match_key_qbytes_0_T_1 ? phv_data_134 : _GEN_621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_623 = 8'h87 == _match_key_qbytes_0_T_1 ? phv_data_135 : _GEN_622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_624 = 8'h88 == _match_key_qbytes_0_T_1 ? phv_data_136 : _GEN_623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_625 = 8'h89 == _match_key_qbytes_0_T_1 ? phv_data_137 : _GEN_624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_626 = 8'h8a == _match_key_qbytes_0_T_1 ? phv_data_138 : _GEN_625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_627 = 8'h8b == _match_key_qbytes_0_T_1 ? phv_data_139 : _GEN_626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_628 = 8'h8c == _match_key_qbytes_0_T_1 ? phv_data_140 : _GEN_627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_629 = 8'h8d == _match_key_qbytes_0_T_1 ? phv_data_141 : _GEN_628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_630 = 8'h8e == _match_key_qbytes_0_T_1 ? phv_data_142 : _GEN_629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_631 = 8'h8f == _match_key_qbytes_0_T_1 ? phv_data_143 : _GEN_630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_632 = 8'h90 == _match_key_qbytes_0_T_1 ? phv_data_144 : _GEN_631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_633 = 8'h91 == _match_key_qbytes_0_T_1 ? phv_data_145 : _GEN_632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_634 = 8'h92 == _match_key_qbytes_0_T_1 ? phv_data_146 : _GEN_633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_635 = 8'h93 == _match_key_qbytes_0_T_1 ? phv_data_147 : _GEN_634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_636 = 8'h94 == _match_key_qbytes_0_T_1 ? phv_data_148 : _GEN_635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_637 = 8'h95 == _match_key_qbytes_0_T_1 ? phv_data_149 : _GEN_636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_638 = 8'h96 == _match_key_qbytes_0_T_1 ? phv_data_150 : _GEN_637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_639 = 8'h97 == _match_key_qbytes_0_T_1 ? phv_data_151 : _GEN_638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_640 = 8'h98 == _match_key_qbytes_0_T_1 ? phv_data_152 : _GEN_639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_641 = 8'h99 == _match_key_qbytes_0_T_1 ? phv_data_153 : _GEN_640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_642 = 8'h9a == _match_key_qbytes_0_T_1 ? phv_data_154 : _GEN_641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_643 = 8'h9b == _match_key_qbytes_0_T_1 ? phv_data_155 : _GEN_642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_644 = 8'h9c == _match_key_qbytes_0_T_1 ? phv_data_156 : _GEN_643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_645 = 8'h9d == _match_key_qbytes_0_T_1 ? phv_data_157 : _GEN_644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_646 = 8'h9e == _match_key_qbytes_0_T_1 ? phv_data_158 : _GEN_645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_647 = 8'h9f == _match_key_qbytes_0_T_1 ? phv_data_159 : _GEN_646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [31:0] _match_key_qbytes_0_T_3 = {_GEN_487,_GEN_647,_GEN_167,_GEN_327}; // @[Cat.scala 30:58]
  wire [31:0] match_key_qbytes_0 = local_offset < end_offset ? _match_key_qbytes_0_T_3 : 32'h0; // @[matcher.scala 88:54 matcher.scala 89:45 matcher.scala 97:45]
  wire [7:0] local_offset_1 = 8'h4 + read_key_offset; // @[matcher.scala 87:77]
  wire [5:0] match_key_qbytes_1_hi = local_offset_1[7:2]; // @[matcher.scala 91:54]
  wire [7:0] _match_key_qbytes_1_T = {match_key_qbytes_1_hi,2'h3}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_1_T_1 = {match_key_qbytes_1_hi,2'h2}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_1_T_2 = {match_key_qbytes_1_hi,2'h1}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_650 = 8'h1 == _match_key_qbytes_1_T_2 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_651 = 8'h2 == _match_key_qbytes_1_T_2 ? phv_data_2 : _GEN_650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_652 = 8'h3 == _match_key_qbytes_1_T_2 ? phv_data_3 : _GEN_651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_653 = 8'h4 == _match_key_qbytes_1_T_2 ? phv_data_4 : _GEN_652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_654 = 8'h5 == _match_key_qbytes_1_T_2 ? phv_data_5 : _GEN_653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_655 = 8'h6 == _match_key_qbytes_1_T_2 ? phv_data_6 : _GEN_654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_656 = 8'h7 == _match_key_qbytes_1_T_2 ? phv_data_7 : _GEN_655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_657 = 8'h8 == _match_key_qbytes_1_T_2 ? phv_data_8 : _GEN_656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_658 = 8'h9 == _match_key_qbytes_1_T_2 ? phv_data_9 : _GEN_657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_659 = 8'ha == _match_key_qbytes_1_T_2 ? phv_data_10 : _GEN_658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_660 = 8'hb == _match_key_qbytes_1_T_2 ? phv_data_11 : _GEN_659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_661 = 8'hc == _match_key_qbytes_1_T_2 ? phv_data_12 : _GEN_660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_662 = 8'hd == _match_key_qbytes_1_T_2 ? phv_data_13 : _GEN_661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_663 = 8'he == _match_key_qbytes_1_T_2 ? phv_data_14 : _GEN_662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_664 = 8'hf == _match_key_qbytes_1_T_2 ? phv_data_15 : _GEN_663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_665 = 8'h10 == _match_key_qbytes_1_T_2 ? phv_data_16 : _GEN_664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_666 = 8'h11 == _match_key_qbytes_1_T_2 ? phv_data_17 : _GEN_665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_667 = 8'h12 == _match_key_qbytes_1_T_2 ? phv_data_18 : _GEN_666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_668 = 8'h13 == _match_key_qbytes_1_T_2 ? phv_data_19 : _GEN_667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_669 = 8'h14 == _match_key_qbytes_1_T_2 ? phv_data_20 : _GEN_668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_670 = 8'h15 == _match_key_qbytes_1_T_2 ? phv_data_21 : _GEN_669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_671 = 8'h16 == _match_key_qbytes_1_T_2 ? phv_data_22 : _GEN_670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_672 = 8'h17 == _match_key_qbytes_1_T_2 ? phv_data_23 : _GEN_671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_673 = 8'h18 == _match_key_qbytes_1_T_2 ? phv_data_24 : _GEN_672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_674 = 8'h19 == _match_key_qbytes_1_T_2 ? phv_data_25 : _GEN_673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_675 = 8'h1a == _match_key_qbytes_1_T_2 ? phv_data_26 : _GEN_674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_676 = 8'h1b == _match_key_qbytes_1_T_2 ? phv_data_27 : _GEN_675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_677 = 8'h1c == _match_key_qbytes_1_T_2 ? phv_data_28 : _GEN_676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_678 = 8'h1d == _match_key_qbytes_1_T_2 ? phv_data_29 : _GEN_677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_679 = 8'h1e == _match_key_qbytes_1_T_2 ? phv_data_30 : _GEN_678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_680 = 8'h1f == _match_key_qbytes_1_T_2 ? phv_data_31 : _GEN_679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_681 = 8'h20 == _match_key_qbytes_1_T_2 ? phv_data_32 : _GEN_680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_682 = 8'h21 == _match_key_qbytes_1_T_2 ? phv_data_33 : _GEN_681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_683 = 8'h22 == _match_key_qbytes_1_T_2 ? phv_data_34 : _GEN_682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_684 = 8'h23 == _match_key_qbytes_1_T_2 ? phv_data_35 : _GEN_683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_685 = 8'h24 == _match_key_qbytes_1_T_2 ? phv_data_36 : _GEN_684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_686 = 8'h25 == _match_key_qbytes_1_T_2 ? phv_data_37 : _GEN_685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_687 = 8'h26 == _match_key_qbytes_1_T_2 ? phv_data_38 : _GEN_686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_688 = 8'h27 == _match_key_qbytes_1_T_2 ? phv_data_39 : _GEN_687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_689 = 8'h28 == _match_key_qbytes_1_T_2 ? phv_data_40 : _GEN_688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_690 = 8'h29 == _match_key_qbytes_1_T_2 ? phv_data_41 : _GEN_689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_691 = 8'h2a == _match_key_qbytes_1_T_2 ? phv_data_42 : _GEN_690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_692 = 8'h2b == _match_key_qbytes_1_T_2 ? phv_data_43 : _GEN_691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_693 = 8'h2c == _match_key_qbytes_1_T_2 ? phv_data_44 : _GEN_692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_694 = 8'h2d == _match_key_qbytes_1_T_2 ? phv_data_45 : _GEN_693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_695 = 8'h2e == _match_key_qbytes_1_T_2 ? phv_data_46 : _GEN_694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_696 = 8'h2f == _match_key_qbytes_1_T_2 ? phv_data_47 : _GEN_695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_697 = 8'h30 == _match_key_qbytes_1_T_2 ? phv_data_48 : _GEN_696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_698 = 8'h31 == _match_key_qbytes_1_T_2 ? phv_data_49 : _GEN_697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_699 = 8'h32 == _match_key_qbytes_1_T_2 ? phv_data_50 : _GEN_698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_700 = 8'h33 == _match_key_qbytes_1_T_2 ? phv_data_51 : _GEN_699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_701 = 8'h34 == _match_key_qbytes_1_T_2 ? phv_data_52 : _GEN_700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_702 = 8'h35 == _match_key_qbytes_1_T_2 ? phv_data_53 : _GEN_701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_703 = 8'h36 == _match_key_qbytes_1_T_2 ? phv_data_54 : _GEN_702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_704 = 8'h37 == _match_key_qbytes_1_T_2 ? phv_data_55 : _GEN_703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_705 = 8'h38 == _match_key_qbytes_1_T_2 ? phv_data_56 : _GEN_704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_706 = 8'h39 == _match_key_qbytes_1_T_2 ? phv_data_57 : _GEN_705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_707 = 8'h3a == _match_key_qbytes_1_T_2 ? phv_data_58 : _GEN_706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_708 = 8'h3b == _match_key_qbytes_1_T_2 ? phv_data_59 : _GEN_707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_709 = 8'h3c == _match_key_qbytes_1_T_2 ? phv_data_60 : _GEN_708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_710 = 8'h3d == _match_key_qbytes_1_T_2 ? phv_data_61 : _GEN_709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_711 = 8'h3e == _match_key_qbytes_1_T_2 ? phv_data_62 : _GEN_710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_712 = 8'h3f == _match_key_qbytes_1_T_2 ? phv_data_63 : _GEN_711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_713 = 8'h40 == _match_key_qbytes_1_T_2 ? phv_data_64 : _GEN_712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_714 = 8'h41 == _match_key_qbytes_1_T_2 ? phv_data_65 : _GEN_713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_715 = 8'h42 == _match_key_qbytes_1_T_2 ? phv_data_66 : _GEN_714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_716 = 8'h43 == _match_key_qbytes_1_T_2 ? phv_data_67 : _GEN_715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_717 = 8'h44 == _match_key_qbytes_1_T_2 ? phv_data_68 : _GEN_716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_718 = 8'h45 == _match_key_qbytes_1_T_2 ? phv_data_69 : _GEN_717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_719 = 8'h46 == _match_key_qbytes_1_T_2 ? phv_data_70 : _GEN_718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_720 = 8'h47 == _match_key_qbytes_1_T_2 ? phv_data_71 : _GEN_719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_721 = 8'h48 == _match_key_qbytes_1_T_2 ? phv_data_72 : _GEN_720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_722 = 8'h49 == _match_key_qbytes_1_T_2 ? phv_data_73 : _GEN_721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_723 = 8'h4a == _match_key_qbytes_1_T_2 ? phv_data_74 : _GEN_722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_724 = 8'h4b == _match_key_qbytes_1_T_2 ? phv_data_75 : _GEN_723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_725 = 8'h4c == _match_key_qbytes_1_T_2 ? phv_data_76 : _GEN_724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_726 = 8'h4d == _match_key_qbytes_1_T_2 ? phv_data_77 : _GEN_725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_727 = 8'h4e == _match_key_qbytes_1_T_2 ? phv_data_78 : _GEN_726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_728 = 8'h4f == _match_key_qbytes_1_T_2 ? phv_data_79 : _GEN_727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_729 = 8'h50 == _match_key_qbytes_1_T_2 ? phv_data_80 : _GEN_728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_730 = 8'h51 == _match_key_qbytes_1_T_2 ? phv_data_81 : _GEN_729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_731 = 8'h52 == _match_key_qbytes_1_T_2 ? phv_data_82 : _GEN_730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_732 = 8'h53 == _match_key_qbytes_1_T_2 ? phv_data_83 : _GEN_731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_733 = 8'h54 == _match_key_qbytes_1_T_2 ? phv_data_84 : _GEN_732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_734 = 8'h55 == _match_key_qbytes_1_T_2 ? phv_data_85 : _GEN_733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_735 = 8'h56 == _match_key_qbytes_1_T_2 ? phv_data_86 : _GEN_734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_736 = 8'h57 == _match_key_qbytes_1_T_2 ? phv_data_87 : _GEN_735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_737 = 8'h58 == _match_key_qbytes_1_T_2 ? phv_data_88 : _GEN_736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_738 = 8'h59 == _match_key_qbytes_1_T_2 ? phv_data_89 : _GEN_737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_739 = 8'h5a == _match_key_qbytes_1_T_2 ? phv_data_90 : _GEN_738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_740 = 8'h5b == _match_key_qbytes_1_T_2 ? phv_data_91 : _GEN_739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_741 = 8'h5c == _match_key_qbytes_1_T_2 ? phv_data_92 : _GEN_740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_742 = 8'h5d == _match_key_qbytes_1_T_2 ? phv_data_93 : _GEN_741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_743 = 8'h5e == _match_key_qbytes_1_T_2 ? phv_data_94 : _GEN_742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_744 = 8'h5f == _match_key_qbytes_1_T_2 ? phv_data_95 : _GEN_743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_745 = 8'h60 == _match_key_qbytes_1_T_2 ? phv_data_96 : _GEN_744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_746 = 8'h61 == _match_key_qbytes_1_T_2 ? phv_data_97 : _GEN_745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_747 = 8'h62 == _match_key_qbytes_1_T_2 ? phv_data_98 : _GEN_746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_748 = 8'h63 == _match_key_qbytes_1_T_2 ? phv_data_99 : _GEN_747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_749 = 8'h64 == _match_key_qbytes_1_T_2 ? phv_data_100 : _GEN_748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_750 = 8'h65 == _match_key_qbytes_1_T_2 ? phv_data_101 : _GEN_749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_751 = 8'h66 == _match_key_qbytes_1_T_2 ? phv_data_102 : _GEN_750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_752 = 8'h67 == _match_key_qbytes_1_T_2 ? phv_data_103 : _GEN_751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_753 = 8'h68 == _match_key_qbytes_1_T_2 ? phv_data_104 : _GEN_752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_754 = 8'h69 == _match_key_qbytes_1_T_2 ? phv_data_105 : _GEN_753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_755 = 8'h6a == _match_key_qbytes_1_T_2 ? phv_data_106 : _GEN_754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_756 = 8'h6b == _match_key_qbytes_1_T_2 ? phv_data_107 : _GEN_755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_757 = 8'h6c == _match_key_qbytes_1_T_2 ? phv_data_108 : _GEN_756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_758 = 8'h6d == _match_key_qbytes_1_T_2 ? phv_data_109 : _GEN_757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_759 = 8'h6e == _match_key_qbytes_1_T_2 ? phv_data_110 : _GEN_758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_760 = 8'h6f == _match_key_qbytes_1_T_2 ? phv_data_111 : _GEN_759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_761 = 8'h70 == _match_key_qbytes_1_T_2 ? phv_data_112 : _GEN_760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_762 = 8'h71 == _match_key_qbytes_1_T_2 ? phv_data_113 : _GEN_761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_763 = 8'h72 == _match_key_qbytes_1_T_2 ? phv_data_114 : _GEN_762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_764 = 8'h73 == _match_key_qbytes_1_T_2 ? phv_data_115 : _GEN_763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_765 = 8'h74 == _match_key_qbytes_1_T_2 ? phv_data_116 : _GEN_764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_766 = 8'h75 == _match_key_qbytes_1_T_2 ? phv_data_117 : _GEN_765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_767 = 8'h76 == _match_key_qbytes_1_T_2 ? phv_data_118 : _GEN_766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_768 = 8'h77 == _match_key_qbytes_1_T_2 ? phv_data_119 : _GEN_767; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_769 = 8'h78 == _match_key_qbytes_1_T_2 ? phv_data_120 : _GEN_768; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_770 = 8'h79 == _match_key_qbytes_1_T_2 ? phv_data_121 : _GEN_769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_771 = 8'h7a == _match_key_qbytes_1_T_2 ? phv_data_122 : _GEN_770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_772 = 8'h7b == _match_key_qbytes_1_T_2 ? phv_data_123 : _GEN_771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_773 = 8'h7c == _match_key_qbytes_1_T_2 ? phv_data_124 : _GEN_772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_774 = 8'h7d == _match_key_qbytes_1_T_2 ? phv_data_125 : _GEN_773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_775 = 8'h7e == _match_key_qbytes_1_T_2 ? phv_data_126 : _GEN_774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_776 = 8'h7f == _match_key_qbytes_1_T_2 ? phv_data_127 : _GEN_775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_777 = 8'h80 == _match_key_qbytes_1_T_2 ? phv_data_128 : _GEN_776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_778 = 8'h81 == _match_key_qbytes_1_T_2 ? phv_data_129 : _GEN_777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_779 = 8'h82 == _match_key_qbytes_1_T_2 ? phv_data_130 : _GEN_778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_780 = 8'h83 == _match_key_qbytes_1_T_2 ? phv_data_131 : _GEN_779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_781 = 8'h84 == _match_key_qbytes_1_T_2 ? phv_data_132 : _GEN_780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_782 = 8'h85 == _match_key_qbytes_1_T_2 ? phv_data_133 : _GEN_781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_783 = 8'h86 == _match_key_qbytes_1_T_2 ? phv_data_134 : _GEN_782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_784 = 8'h87 == _match_key_qbytes_1_T_2 ? phv_data_135 : _GEN_783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_785 = 8'h88 == _match_key_qbytes_1_T_2 ? phv_data_136 : _GEN_784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_786 = 8'h89 == _match_key_qbytes_1_T_2 ? phv_data_137 : _GEN_785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_787 = 8'h8a == _match_key_qbytes_1_T_2 ? phv_data_138 : _GEN_786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_788 = 8'h8b == _match_key_qbytes_1_T_2 ? phv_data_139 : _GEN_787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_789 = 8'h8c == _match_key_qbytes_1_T_2 ? phv_data_140 : _GEN_788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_790 = 8'h8d == _match_key_qbytes_1_T_2 ? phv_data_141 : _GEN_789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_791 = 8'h8e == _match_key_qbytes_1_T_2 ? phv_data_142 : _GEN_790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_792 = 8'h8f == _match_key_qbytes_1_T_2 ? phv_data_143 : _GEN_791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_793 = 8'h90 == _match_key_qbytes_1_T_2 ? phv_data_144 : _GEN_792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_794 = 8'h91 == _match_key_qbytes_1_T_2 ? phv_data_145 : _GEN_793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_795 = 8'h92 == _match_key_qbytes_1_T_2 ? phv_data_146 : _GEN_794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_796 = 8'h93 == _match_key_qbytes_1_T_2 ? phv_data_147 : _GEN_795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_797 = 8'h94 == _match_key_qbytes_1_T_2 ? phv_data_148 : _GEN_796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_798 = 8'h95 == _match_key_qbytes_1_T_2 ? phv_data_149 : _GEN_797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_799 = 8'h96 == _match_key_qbytes_1_T_2 ? phv_data_150 : _GEN_798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_800 = 8'h97 == _match_key_qbytes_1_T_2 ? phv_data_151 : _GEN_799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_801 = 8'h98 == _match_key_qbytes_1_T_2 ? phv_data_152 : _GEN_800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_802 = 8'h99 == _match_key_qbytes_1_T_2 ? phv_data_153 : _GEN_801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_803 = 8'h9a == _match_key_qbytes_1_T_2 ? phv_data_154 : _GEN_802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_804 = 8'h9b == _match_key_qbytes_1_T_2 ? phv_data_155 : _GEN_803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_805 = 8'h9c == _match_key_qbytes_1_T_2 ? phv_data_156 : _GEN_804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_806 = 8'h9d == _match_key_qbytes_1_T_2 ? phv_data_157 : _GEN_805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_807 = 8'h9e == _match_key_qbytes_1_T_2 ? phv_data_158 : _GEN_806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_808 = 8'h9f == _match_key_qbytes_1_T_2 ? phv_data_159 : _GEN_807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_810 = 8'h1 == local_offset_1 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_811 = 8'h2 == local_offset_1 ? phv_data_2 : _GEN_810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_812 = 8'h3 == local_offset_1 ? phv_data_3 : _GEN_811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_813 = 8'h4 == local_offset_1 ? phv_data_4 : _GEN_812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_814 = 8'h5 == local_offset_1 ? phv_data_5 : _GEN_813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_815 = 8'h6 == local_offset_1 ? phv_data_6 : _GEN_814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_816 = 8'h7 == local_offset_1 ? phv_data_7 : _GEN_815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_817 = 8'h8 == local_offset_1 ? phv_data_8 : _GEN_816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_818 = 8'h9 == local_offset_1 ? phv_data_9 : _GEN_817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_819 = 8'ha == local_offset_1 ? phv_data_10 : _GEN_818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_820 = 8'hb == local_offset_1 ? phv_data_11 : _GEN_819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_821 = 8'hc == local_offset_1 ? phv_data_12 : _GEN_820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_822 = 8'hd == local_offset_1 ? phv_data_13 : _GEN_821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_823 = 8'he == local_offset_1 ? phv_data_14 : _GEN_822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_824 = 8'hf == local_offset_1 ? phv_data_15 : _GEN_823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_825 = 8'h10 == local_offset_1 ? phv_data_16 : _GEN_824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_826 = 8'h11 == local_offset_1 ? phv_data_17 : _GEN_825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_827 = 8'h12 == local_offset_1 ? phv_data_18 : _GEN_826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_828 = 8'h13 == local_offset_1 ? phv_data_19 : _GEN_827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_829 = 8'h14 == local_offset_1 ? phv_data_20 : _GEN_828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_830 = 8'h15 == local_offset_1 ? phv_data_21 : _GEN_829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_831 = 8'h16 == local_offset_1 ? phv_data_22 : _GEN_830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_832 = 8'h17 == local_offset_1 ? phv_data_23 : _GEN_831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_833 = 8'h18 == local_offset_1 ? phv_data_24 : _GEN_832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_834 = 8'h19 == local_offset_1 ? phv_data_25 : _GEN_833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_835 = 8'h1a == local_offset_1 ? phv_data_26 : _GEN_834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_836 = 8'h1b == local_offset_1 ? phv_data_27 : _GEN_835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_837 = 8'h1c == local_offset_1 ? phv_data_28 : _GEN_836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_838 = 8'h1d == local_offset_1 ? phv_data_29 : _GEN_837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_839 = 8'h1e == local_offset_1 ? phv_data_30 : _GEN_838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_840 = 8'h1f == local_offset_1 ? phv_data_31 : _GEN_839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_841 = 8'h20 == local_offset_1 ? phv_data_32 : _GEN_840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_842 = 8'h21 == local_offset_1 ? phv_data_33 : _GEN_841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_843 = 8'h22 == local_offset_1 ? phv_data_34 : _GEN_842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_844 = 8'h23 == local_offset_1 ? phv_data_35 : _GEN_843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_845 = 8'h24 == local_offset_1 ? phv_data_36 : _GEN_844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_846 = 8'h25 == local_offset_1 ? phv_data_37 : _GEN_845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_847 = 8'h26 == local_offset_1 ? phv_data_38 : _GEN_846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_848 = 8'h27 == local_offset_1 ? phv_data_39 : _GEN_847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_849 = 8'h28 == local_offset_1 ? phv_data_40 : _GEN_848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_850 = 8'h29 == local_offset_1 ? phv_data_41 : _GEN_849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_851 = 8'h2a == local_offset_1 ? phv_data_42 : _GEN_850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_852 = 8'h2b == local_offset_1 ? phv_data_43 : _GEN_851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_853 = 8'h2c == local_offset_1 ? phv_data_44 : _GEN_852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_854 = 8'h2d == local_offset_1 ? phv_data_45 : _GEN_853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_855 = 8'h2e == local_offset_1 ? phv_data_46 : _GEN_854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_856 = 8'h2f == local_offset_1 ? phv_data_47 : _GEN_855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_857 = 8'h30 == local_offset_1 ? phv_data_48 : _GEN_856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_858 = 8'h31 == local_offset_1 ? phv_data_49 : _GEN_857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_859 = 8'h32 == local_offset_1 ? phv_data_50 : _GEN_858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_860 = 8'h33 == local_offset_1 ? phv_data_51 : _GEN_859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_861 = 8'h34 == local_offset_1 ? phv_data_52 : _GEN_860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_862 = 8'h35 == local_offset_1 ? phv_data_53 : _GEN_861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_863 = 8'h36 == local_offset_1 ? phv_data_54 : _GEN_862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_864 = 8'h37 == local_offset_1 ? phv_data_55 : _GEN_863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_865 = 8'h38 == local_offset_1 ? phv_data_56 : _GEN_864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_866 = 8'h39 == local_offset_1 ? phv_data_57 : _GEN_865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_867 = 8'h3a == local_offset_1 ? phv_data_58 : _GEN_866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_868 = 8'h3b == local_offset_1 ? phv_data_59 : _GEN_867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_869 = 8'h3c == local_offset_1 ? phv_data_60 : _GEN_868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_870 = 8'h3d == local_offset_1 ? phv_data_61 : _GEN_869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_871 = 8'h3e == local_offset_1 ? phv_data_62 : _GEN_870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_872 = 8'h3f == local_offset_1 ? phv_data_63 : _GEN_871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_873 = 8'h40 == local_offset_1 ? phv_data_64 : _GEN_872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_874 = 8'h41 == local_offset_1 ? phv_data_65 : _GEN_873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_875 = 8'h42 == local_offset_1 ? phv_data_66 : _GEN_874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_876 = 8'h43 == local_offset_1 ? phv_data_67 : _GEN_875; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_877 = 8'h44 == local_offset_1 ? phv_data_68 : _GEN_876; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_878 = 8'h45 == local_offset_1 ? phv_data_69 : _GEN_877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_879 = 8'h46 == local_offset_1 ? phv_data_70 : _GEN_878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_880 = 8'h47 == local_offset_1 ? phv_data_71 : _GEN_879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_881 = 8'h48 == local_offset_1 ? phv_data_72 : _GEN_880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_882 = 8'h49 == local_offset_1 ? phv_data_73 : _GEN_881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_883 = 8'h4a == local_offset_1 ? phv_data_74 : _GEN_882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_884 = 8'h4b == local_offset_1 ? phv_data_75 : _GEN_883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_885 = 8'h4c == local_offset_1 ? phv_data_76 : _GEN_884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_886 = 8'h4d == local_offset_1 ? phv_data_77 : _GEN_885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_887 = 8'h4e == local_offset_1 ? phv_data_78 : _GEN_886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_888 = 8'h4f == local_offset_1 ? phv_data_79 : _GEN_887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_889 = 8'h50 == local_offset_1 ? phv_data_80 : _GEN_888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_890 = 8'h51 == local_offset_1 ? phv_data_81 : _GEN_889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_891 = 8'h52 == local_offset_1 ? phv_data_82 : _GEN_890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_892 = 8'h53 == local_offset_1 ? phv_data_83 : _GEN_891; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_893 = 8'h54 == local_offset_1 ? phv_data_84 : _GEN_892; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_894 = 8'h55 == local_offset_1 ? phv_data_85 : _GEN_893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_895 = 8'h56 == local_offset_1 ? phv_data_86 : _GEN_894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_896 = 8'h57 == local_offset_1 ? phv_data_87 : _GEN_895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_897 = 8'h58 == local_offset_1 ? phv_data_88 : _GEN_896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_898 = 8'h59 == local_offset_1 ? phv_data_89 : _GEN_897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_899 = 8'h5a == local_offset_1 ? phv_data_90 : _GEN_898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_900 = 8'h5b == local_offset_1 ? phv_data_91 : _GEN_899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_901 = 8'h5c == local_offset_1 ? phv_data_92 : _GEN_900; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_902 = 8'h5d == local_offset_1 ? phv_data_93 : _GEN_901; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_903 = 8'h5e == local_offset_1 ? phv_data_94 : _GEN_902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_904 = 8'h5f == local_offset_1 ? phv_data_95 : _GEN_903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_905 = 8'h60 == local_offset_1 ? phv_data_96 : _GEN_904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_906 = 8'h61 == local_offset_1 ? phv_data_97 : _GEN_905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_907 = 8'h62 == local_offset_1 ? phv_data_98 : _GEN_906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_908 = 8'h63 == local_offset_1 ? phv_data_99 : _GEN_907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_909 = 8'h64 == local_offset_1 ? phv_data_100 : _GEN_908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_910 = 8'h65 == local_offset_1 ? phv_data_101 : _GEN_909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_911 = 8'h66 == local_offset_1 ? phv_data_102 : _GEN_910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_912 = 8'h67 == local_offset_1 ? phv_data_103 : _GEN_911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_913 = 8'h68 == local_offset_1 ? phv_data_104 : _GEN_912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_914 = 8'h69 == local_offset_1 ? phv_data_105 : _GEN_913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_915 = 8'h6a == local_offset_1 ? phv_data_106 : _GEN_914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_916 = 8'h6b == local_offset_1 ? phv_data_107 : _GEN_915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_917 = 8'h6c == local_offset_1 ? phv_data_108 : _GEN_916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_918 = 8'h6d == local_offset_1 ? phv_data_109 : _GEN_917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_919 = 8'h6e == local_offset_1 ? phv_data_110 : _GEN_918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_920 = 8'h6f == local_offset_1 ? phv_data_111 : _GEN_919; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_921 = 8'h70 == local_offset_1 ? phv_data_112 : _GEN_920; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_922 = 8'h71 == local_offset_1 ? phv_data_113 : _GEN_921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_923 = 8'h72 == local_offset_1 ? phv_data_114 : _GEN_922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_924 = 8'h73 == local_offset_1 ? phv_data_115 : _GEN_923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_925 = 8'h74 == local_offset_1 ? phv_data_116 : _GEN_924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_926 = 8'h75 == local_offset_1 ? phv_data_117 : _GEN_925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_927 = 8'h76 == local_offset_1 ? phv_data_118 : _GEN_926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_928 = 8'h77 == local_offset_1 ? phv_data_119 : _GEN_927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_929 = 8'h78 == local_offset_1 ? phv_data_120 : _GEN_928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_930 = 8'h79 == local_offset_1 ? phv_data_121 : _GEN_929; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_931 = 8'h7a == local_offset_1 ? phv_data_122 : _GEN_930; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_932 = 8'h7b == local_offset_1 ? phv_data_123 : _GEN_931; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_933 = 8'h7c == local_offset_1 ? phv_data_124 : _GEN_932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_934 = 8'h7d == local_offset_1 ? phv_data_125 : _GEN_933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_935 = 8'h7e == local_offset_1 ? phv_data_126 : _GEN_934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_936 = 8'h7f == local_offset_1 ? phv_data_127 : _GEN_935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_937 = 8'h80 == local_offset_1 ? phv_data_128 : _GEN_936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_938 = 8'h81 == local_offset_1 ? phv_data_129 : _GEN_937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_939 = 8'h82 == local_offset_1 ? phv_data_130 : _GEN_938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_940 = 8'h83 == local_offset_1 ? phv_data_131 : _GEN_939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_941 = 8'h84 == local_offset_1 ? phv_data_132 : _GEN_940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_942 = 8'h85 == local_offset_1 ? phv_data_133 : _GEN_941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_943 = 8'h86 == local_offset_1 ? phv_data_134 : _GEN_942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_944 = 8'h87 == local_offset_1 ? phv_data_135 : _GEN_943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_945 = 8'h88 == local_offset_1 ? phv_data_136 : _GEN_944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_946 = 8'h89 == local_offset_1 ? phv_data_137 : _GEN_945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_947 = 8'h8a == local_offset_1 ? phv_data_138 : _GEN_946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_948 = 8'h8b == local_offset_1 ? phv_data_139 : _GEN_947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_949 = 8'h8c == local_offset_1 ? phv_data_140 : _GEN_948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_950 = 8'h8d == local_offset_1 ? phv_data_141 : _GEN_949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_951 = 8'h8e == local_offset_1 ? phv_data_142 : _GEN_950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_952 = 8'h8f == local_offset_1 ? phv_data_143 : _GEN_951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_953 = 8'h90 == local_offset_1 ? phv_data_144 : _GEN_952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_954 = 8'h91 == local_offset_1 ? phv_data_145 : _GEN_953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_955 = 8'h92 == local_offset_1 ? phv_data_146 : _GEN_954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_956 = 8'h93 == local_offset_1 ? phv_data_147 : _GEN_955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_957 = 8'h94 == local_offset_1 ? phv_data_148 : _GEN_956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_958 = 8'h95 == local_offset_1 ? phv_data_149 : _GEN_957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_959 = 8'h96 == local_offset_1 ? phv_data_150 : _GEN_958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_960 = 8'h97 == local_offset_1 ? phv_data_151 : _GEN_959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_961 = 8'h98 == local_offset_1 ? phv_data_152 : _GEN_960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_962 = 8'h99 == local_offset_1 ? phv_data_153 : _GEN_961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_963 = 8'h9a == local_offset_1 ? phv_data_154 : _GEN_962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_964 = 8'h9b == local_offset_1 ? phv_data_155 : _GEN_963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_965 = 8'h9c == local_offset_1 ? phv_data_156 : _GEN_964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_966 = 8'h9d == local_offset_1 ? phv_data_157 : _GEN_965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_967 = 8'h9e == local_offset_1 ? phv_data_158 : _GEN_966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_968 = 8'h9f == local_offset_1 ? phv_data_159 : _GEN_967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_970 = 8'h1 == _match_key_qbytes_1_T ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_971 = 8'h2 == _match_key_qbytes_1_T ? phv_data_2 : _GEN_970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_972 = 8'h3 == _match_key_qbytes_1_T ? phv_data_3 : _GEN_971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_973 = 8'h4 == _match_key_qbytes_1_T ? phv_data_4 : _GEN_972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_974 = 8'h5 == _match_key_qbytes_1_T ? phv_data_5 : _GEN_973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_975 = 8'h6 == _match_key_qbytes_1_T ? phv_data_6 : _GEN_974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_976 = 8'h7 == _match_key_qbytes_1_T ? phv_data_7 : _GEN_975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_977 = 8'h8 == _match_key_qbytes_1_T ? phv_data_8 : _GEN_976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_978 = 8'h9 == _match_key_qbytes_1_T ? phv_data_9 : _GEN_977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_979 = 8'ha == _match_key_qbytes_1_T ? phv_data_10 : _GEN_978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_980 = 8'hb == _match_key_qbytes_1_T ? phv_data_11 : _GEN_979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_981 = 8'hc == _match_key_qbytes_1_T ? phv_data_12 : _GEN_980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_982 = 8'hd == _match_key_qbytes_1_T ? phv_data_13 : _GEN_981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_983 = 8'he == _match_key_qbytes_1_T ? phv_data_14 : _GEN_982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_984 = 8'hf == _match_key_qbytes_1_T ? phv_data_15 : _GEN_983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_985 = 8'h10 == _match_key_qbytes_1_T ? phv_data_16 : _GEN_984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_986 = 8'h11 == _match_key_qbytes_1_T ? phv_data_17 : _GEN_985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_987 = 8'h12 == _match_key_qbytes_1_T ? phv_data_18 : _GEN_986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_988 = 8'h13 == _match_key_qbytes_1_T ? phv_data_19 : _GEN_987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_989 = 8'h14 == _match_key_qbytes_1_T ? phv_data_20 : _GEN_988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_990 = 8'h15 == _match_key_qbytes_1_T ? phv_data_21 : _GEN_989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_991 = 8'h16 == _match_key_qbytes_1_T ? phv_data_22 : _GEN_990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_992 = 8'h17 == _match_key_qbytes_1_T ? phv_data_23 : _GEN_991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_993 = 8'h18 == _match_key_qbytes_1_T ? phv_data_24 : _GEN_992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_994 = 8'h19 == _match_key_qbytes_1_T ? phv_data_25 : _GEN_993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_995 = 8'h1a == _match_key_qbytes_1_T ? phv_data_26 : _GEN_994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_996 = 8'h1b == _match_key_qbytes_1_T ? phv_data_27 : _GEN_995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_997 = 8'h1c == _match_key_qbytes_1_T ? phv_data_28 : _GEN_996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_998 = 8'h1d == _match_key_qbytes_1_T ? phv_data_29 : _GEN_997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_999 = 8'h1e == _match_key_qbytes_1_T ? phv_data_30 : _GEN_998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1000 = 8'h1f == _match_key_qbytes_1_T ? phv_data_31 : _GEN_999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1001 = 8'h20 == _match_key_qbytes_1_T ? phv_data_32 : _GEN_1000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1002 = 8'h21 == _match_key_qbytes_1_T ? phv_data_33 : _GEN_1001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1003 = 8'h22 == _match_key_qbytes_1_T ? phv_data_34 : _GEN_1002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1004 = 8'h23 == _match_key_qbytes_1_T ? phv_data_35 : _GEN_1003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1005 = 8'h24 == _match_key_qbytes_1_T ? phv_data_36 : _GEN_1004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1006 = 8'h25 == _match_key_qbytes_1_T ? phv_data_37 : _GEN_1005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1007 = 8'h26 == _match_key_qbytes_1_T ? phv_data_38 : _GEN_1006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1008 = 8'h27 == _match_key_qbytes_1_T ? phv_data_39 : _GEN_1007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1009 = 8'h28 == _match_key_qbytes_1_T ? phv_data_40 : _GEN_1008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1010 = 8'h29 == _match_key_qbytes_1_T ? phv_data_41 : _GEN_1009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1011 = 8'h2a == _match_key_qbytes_1_T ? phv_data_42 : _GEN_1010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1012 = 8'h2b == _match_key_qbytes_1_T ? phv_data_43 : _GEN_1011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1013 = 8'h2c == _match_key_qbytes_1_T ? phv_data_44 : _GEN_1012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1014 = 8'h2d == _match_key_qbytes_1_T ? phv_data_45 : _GEN_1013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1015 = 8'h2e == _match_key_qbytes_1_T ? phv_data_46 : _GEN_1014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1016 = 8'h2f == _match_key_qbytes_1_T ? phv_data_47 : _GEN_1015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1017 = 8'h30 == _match_key_qbytes_1_T ? phv_data_48 : _GEN_1016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1018 = 8'h31 == _match_key_qbytes_1_T ? phv_data_49 : _GEN_1017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1019 = 8'h32 == _match_key_qbytes_1_T ? phv_data_50 : _GEN_1018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1020 = 8'h33 == _match_key_qbytes_1_T ? phv_data_51 : _GEN_1019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1021 = 8'h34 == _match_key_qbytes_1_T ? phv_data_52 : _GEN_1020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1022 = 8'h35 == _match_key_qbytes_1_T ? phv_data_53 : _GEN_1021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1023 = 8'h36 == _match_key_qbytes_1_T ? phv_data_54 : _GEN_1022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1024 = 8'h37 == _match_key_qbytes_1_T ? phv_data_55 : _GEN_1023; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1025 = 8'h38 == _match_key_qbytes_1_T ? phv_data_56 : _GEN_1024; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1026 = 8'h39 == _match_key_qbytes_1_T ? phv_data_57 : _GEN_1025; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1027 = 8'h3a == _match_key_qbytes_1_T ? phv_data_58 : _GEN_1026; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1028 = 8'h3b == _match_key_qbytes_1_T ? phv_data_59 : _GEN_1027; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1029 = 8'h3c == _match_key_qbytes_1_T ? phv_data_60 : _GEN_1028; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1030 = 8'h3d == _match_key_qbytes_1_T ? phv_data_61 : _GEN_1029; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1031 = 8'h3e == _match_key_qbytes_1_T ? phv_data_62 : _GEN_1030; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1032 = 8'h3f == _match_key_qbytes_1_T ? phv_data_63 : _GEN_1031; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1033 = 8'h40 == _match_key_qbytes_1_T ? phv_data_64 : _GEN_1032; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1034 = 8'h41 == _match_key_qbytes_1_T ? phv_data_65 : _GEN_1033; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1035 = 8'h42 == _match_key_qbytes_1_T ? phv_data_66 : _GEN_1034; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1036 = 8'h43 == _match_key_qbytes_1_T ? phv_data_67 : _GEN_1035; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1037 = 8'h44 == _match_key_qbytes_1_T ? phv_data_68 : _GEN_1036; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1038 = 8'h45 == _match_key_qbytes_1_T ? phv_data_69 : _GEN_1037; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1039 = 8'h46 == _match_key_qbytes_1_T ? phv_data_70 : _GEN_1038; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1040 = 8'h47 == _match_key_qbytes_1_T ? phv_data_71 : _GEN_1039; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1041 = 8'h48 == _match_key_qbytes_1_T ? phv_data_72 : _GEN_1040; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1042 = 8'h49 == _match_key_qbytes_1_T ? phv_data_73 : _GEN_1041; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1043 = 8'h4a == _match_key_qbytes_1_T ? phv_data_74 : _GEN_1042; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1044 = 8'h4b == _match_key_qbytes_1_T ? phv_data_75 : _GEN_1043; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1045 = 8'h4c == _match_key_qbytes_1_T ? phv_data_76 : _GEN_1044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1046 = 8'h4d == _match_key_qbytes_1_T ? phv_data_77 : _GEN_1045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1047 = 8'h4e == _match_key_qbytes_1_T ? phv_data_78 : _GEN_1046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1048 = 8'h4f == _match_key_qbytes_1_T ? phv_data_79 : _GEN_1047; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1049 = 8'h50 == _match_key_qbytes_1_T ? phv_data_80 : _GEN_1048; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1050 = 8'h51 == _match_key_qbytes_1_T ? phv_data_81 : _GEN_1049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1051 = 8'h52 == _match_key_qbytes_1_T ? phv_data_82 : _GEN_1050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1052 = 8'h53 == _match_key_qbytes_1_T ? phv_data_83 : _GEN_1051; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1053 = 8'h54 == _match_key_qbytes_1_T ? phv_data_84 : _GEN_1052; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1054 = 8'h55 == _match_key_qbytes_1_T ? phv_data_85 : _GEN_1053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1055 = 8'h56 == _match_key_qbytes_1_T ? phv_data_86 : _GEN_1054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1056 = 8'h57 == _match_key_qbytes_1_T ? phv_data_87 : _GEN_1055; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1057 = 8'h58 == _match_key_qbytes_1_T ? phv_data_88 : _GEN_1056; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1058 = 8'h59 == _match_key_qbytes_1_T ? phv_data_89 : _GEN_1057; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1059 = 8'h5a == _match_key_qbytes_1_T ? phv_data_90 : _GEN_1058; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1060 = 8'h5b == _match_key_qbytes_1_T ? phv_data_91 : _GEN_1059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1061 = 8'h5c == _match_key_qbytes_1_T ? phv_data_92 : _GEN_1060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1062 = 8'h5d == _match_key_qbytes_1_T ? phv_data_93 : _GEN_1061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1063 = 8'h5e == _match_key_qbytes_1_T ? phv_data_94 : _GEN_1062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1064 = 8'h5f == _match_key_qbytes_1_T ? phv_data_95 : _GEN_1063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1065 = 8'h60 == _match_key_qbytes_1_T ? phv_data_96 : _GEN_1064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1066 = 8'h61 == _match_key_qbytes_1_T ? phv_data_97 : _GEN_1065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1067 = 8'h62 == _match_key_qbytes_1_T ? phv_data_98 : _GEN_1066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1068 = 8'h63 == _match_key_qbytes_1_T ? phv_data_99 : _GEN_1067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1069 = 8'h64 == _match_key_qbytes_1_T ? phv_data_100 : _GEN_1068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1070 = 8'h65 == _match_key_qbytes_1_T ? phv_data_101 : _GEN_1069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1071 = 8'h66 == _match_key_qbytes_1_T ? phv_data_102 : _GEN_1070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1072 = 8'h67 == _match_key_qbytes_1_T ? phv_data_103 : _GEN_1071; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1073 = 8'h68 == _match_key_qbytes_1_T ? phv_data_104 : _GEN_1072; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1074 = 8'h69 == _match_key_qbytes_1_T ? phv_data_105 : _GEN_1073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1075 = 8'h6a == _match_key_qbytes_1_T ? phv_data_106 : _GEN_1074; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1076 = 8'h6b == _match_key_qbytes_1_T ? phv_data_107 : _GEN_1075; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1077 = 8'h6c == _match_key_qbytes_1_T ? phv_data_108 : _GEN_1076; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1078 = 8'h6d == _match_key_qbytes_1_T ? phv_data_109 : _GEN_1077; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1079 = 8'h6e == _match_key_qbytes_1_T ? phv_data_110 : _GEN_1078; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1080 = 8'h6f == _match_key_qbytes_1_T ? phv_data_111 : _GEN_1079; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1081 = 8'h70 == _match_key_qbytes_1_T ? phv_data_112 : _GEN_1080; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1082 = 8'h71 == _match_key_qbytes_1_T ? phv_data_113 : _GEN_1081; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1083 = 8'h72 == _match_key_qbytes_1_T ? phv_data_114 : _GEN_1082; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1084 = 8'h73 == _match_key_qbytes_1_T ? phv_data_115 : _GEN_1083; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1085 = 8'h74 == _match_key_qbytes_1_T ? phv_data_116 : _GEN_1084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1086 = 8'h75 == _match_key_qbytes_1_T ? phv_data_117 : _GEN_1085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1087 = 8'h76 == _match_key_qbytes_1_T ? phv_data_118 : _GEN_1086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1088 = 8'h77 == _match_key_qbytes_1_T ? phv_data_119 : _GEN_1087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1089 = 8'h78 == _match_key_qbytes_1_T ? phv_data_120 : _GEN_1088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1090 = 8'h79 == _match_key_qbytes_1_T ? phv_data_121 : _GEN_1089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1091 = 8'h7a == _match_key_qbytes_1_T ? phv_data_122 : _GEN_1090; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1092 = 8'h7b == _match_key_qbytes_1_T ? phv_data_123 : _GEN_1091; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1093 = 8'h7c == _match_key_qbytes_1_T ? phv_data_124 : _GEN_1092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1094 = 8'h7d == _match_key_qbytes_1_T ? phv_data_125 : _GEN_1093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1095 = 8'h7e == _match_key_qbytes_1_T ? phv_data_126 : _GEN_1094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1096 = 8'h7f == _match_key_qbytes_1_T ? phv_data_127 : _GEN_1095; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1097 = 8'h80 == _match_key_qbytes_1_T ? phv_data_128 : _GEN_1096; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1098 = 8'h81 == _match_key_qbytes_1_T ? phv_data_129 : _GEN_1097; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1099 = 8'h82 == _match_key_qbytes_1_T ? phv_data_130 : _GEN_1098; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1100 = 8'h83 == _match_key_qbytes_1_T ? phv_data_131 : _GEN_1099; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1101 = 8'h84 == _match_key_qbytes_1_T ? phv_data_132 : _GEN_1100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1102 = 8'h85 == _match_key_qbytes_1_T ? phv_data_133 : _GEN_1101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1103 = 8'h86 == _match_key_qbytes_1_T ? phv_data_134 : _GEN_1102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1104 = 8'h87 == _match_key_qbytes_1_T ? phv_data_135 : _GEN_1103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1105 = 8'h88 == _match_key_qbytes_1_T ? phv_data_136 : _GEN_1104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1106 = 8'h89 == _match_key_qbytes_1_T ? phv_data_137 : _GEN_1105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1107 = 8'h8a == _match_key_qbytes_1_T ? phv_data_138 : _GEN_1106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1108 = 8'h8b == _match_key_qbytes_1_T ? phv_data_139 : _GEN_1107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1109 = 8'h8c == _match_key_qbytes_1_T ? phv_data_140 : _GEN_1108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1110 = 8'h8d == _match_key_qbytes_1_T ? phv_data_141 : _GEN_1109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1111 = 8'h8e == _match_key_qbytes_1_T ? phv_data_142 : _GEN_1110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1112 = 8'h8f == _match_key_qbytes_1_T ? phv_data_143 : _GEN_1111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1113 = 8'h90 == _match_key_qbytes_1_T ? phv_data_144 : _GEN_1112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1114 = 8'h91 == _match_key_qbytes_1_T ? phv_data_145 : _GEN_1113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1115 = 8'h92 == _match_key_qbytes_1_T ? phv_data_146 : _GEN_1114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1116 = 8'h93 == _match_key_qbytes_1_T ? phv_data_147 : _GEN_1115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1117 = 8'h94 == _match_key_qbytes_1_T ? phv_data_148 : _GEN_1116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1118 = 8'h95 == _match_key_qbytes_1_T ? phv_data_149 : _GEN_1117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1119 = 8'h96 == _match_key_qbytes_1_T ? phv_data_150 : _GEN_1118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1120 = 8'h97 == _match_key_qbytes_1_T ? phv_data_151 : _GEN_1119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1121 = 8'h98 == _match_key_qbytes_1_T ? phv_data_152 : _GEN_1120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1122 = 8'h99 == _match_key_qbytes_1_T ? phv_data_153 : _GEN_1121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1123 = 8'h9a == _match_key_qbytes_1_T ? phv_data_154 : _GEN_1122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1124 = 8'h9b == _match_key_qbytes_1_T ? phv_data_155 : _GEN_1123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1125 = 8'h9c == _match_key_qbytes_1_T ? phv_data_156 : _GEN_1124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1126 = 8'h9d == _match_key_qbytes_1_T ? phv_data_157 : _GEN_1125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1127 = 8'h9e == _match_key_qbytes_1_T ? phv_data_158 : _GEN_1126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1128 = 8'h9f == _match_key_qbytes_1_T ? phv_data_159 : _GEN_1127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1130 = 8'h1 == _match_key_qbytes_1_T_1 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1131 = 8'h2 == _match_key_qbytes_1_T_1 ? phv_data_2 : _GEN_1130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1132 = 8'h3 == _match_key_qbytes_1_T_1 ? phv_data_3 : _GEN_1131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1133 = 8'h4 == _match_key_qbytes_1_T_1 ? phv_data_4 : _GEN_1132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1134 = 8'h5 == _match_key_qbytes_1_T_1 ? phv_data_5 : _GEN_1133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1135 = 8'h6 == _match_key_qbytes_1_T_1 ? phv_data_6 : _GEN_1134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1136 = 8'h7 == _match_key_qbytes_1_T_1 ? phv_data_7 : _GEN_1135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1137 = 8'h8 == _match_key_qbytes_1_T_1 ? phv_data_8 : _GEN_1136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1138 = 8'h9 == _match_key_qbytes_1_T_1 ? phv_data_9 : _GEN_1137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1139 = 8'ha == _match_key_qbytes_1_T_1 ? phv_data_10 : _GEN_1138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1140 = 8'hb == _match_key_qbytes_1_T_1 ? phv_data_11 : _GEN_1139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1141 = 8'hc == _match_key_qbytes_1_T_1 ? phv_data_12 : _GEN_1140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1142 = 8'hd == _match_key_qbytes_1_T_1 ? phv_data_13 : _GEN_1141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1143 = 8'he == _match_key_qbytes_1_T_1 ? phv_data_14 : _GEN_1142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1144 = 8'hf == _match_key_qbytes_1_T_1 ? phv_data_15 : _GEN_1143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1145 = 8'h10 == _match_key_qbytes_1_T_1 ? phv_data_16 : _GEN_1144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1146 = 8'h11 == _match_key_qbytes_1_T_1 ? phv_data_17 : _GEN_1145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1147 = 8'h12 == _match_key_qbytes_1_T_1 ? phv_data_18 : _GEN_1146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1148 = 8'h13 == _match_key_qbytes_1_T_1 ? phv_data_19 : _GEN_1147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1149 = 8'h14 == _match_key_qbytes_1_T_1 ? phv_data_20 : _GEN_1148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1150 = 8'h15 == _match_key_qbytes_1_T_1 ? phv_data_21 : _GEN_1149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1151 = 8'h16 == _match_key_qbytes_1_T_1 ? phv_data_22 : _GEN_1150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1152 = 8'h17 == _match_key_qbytes_1_T_1 ? phv_data_23 : _GEN_1151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1153 = 8'h18 == _match_key_qbytes_1_T_1 ? phv_data_24 : _GEN_1152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1154 = 8'h19 == _match_key_qbytes_1_T_1 ? phv_data_25 : _GEN_1153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1155 = 8'h1a == _match_key_qbytes_1_T_1 ? phv_data_26 : _GEN_1154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1156 = 8'h1b == _match_key_qbytes_1_T_1 ? phv_data_27 : _GEN_1155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1157 = 8'h1c == _match_key_qbytes_1_T_1 ? phv_data_28 : _GEN_1156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1158 = 8'h1d == _match_key_qbytes_1_T_1 ? phv_data_29 : _GEN_1157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1159 = 8'h1e == _match_key_qbytes_1_T_1 ? phv_data_30 : _GEN_1158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1160 = 8'h1f == _match_key_qbytes_1_T_1 ? phv_data_31 : _GEN_1159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1161 = 8'h20 == _match_key_qbytes_1_T_1 ? phv_data_32 : _GEN_1160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1162 = 8'h21 == _match_key_qbytes_1_T_1 ? phv_data_33 : _GEN_1161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1163 = 8'h22 == _match_key_qbytes_1_T_1 ? phv_data_34 : _GEN_1162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1164 = 8'h23 == _match_key_qbytes_1_T_1 ? phv_data_35 : _GEN_1163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1165 = 8'h24 == _match_key_qbytes_1_T_1 ? phv_data_36 : _GEN_1164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1166 = 8'h25 == _match_key_qbytes_1_T_1 ? phv_data_37 : _GEN_1165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1167 = 8'h26 == _match_key_qbytes_1_T_1 ? phv_data_38 : _GEN_1166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1168 = 8'h27 == _match_key_qbytes_1_T_1 ? phv_data_39 : _GEN_1167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1169 = 8'h28 == _match_key_qbytes_1_T_1 ? phv_data_40 : _GEN_1168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1170 = 8'h29 == _match_key_qbytes_1_T_1 ? phv_data_41 : _GEN_1169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1171 = 8'h2a == _match_key_qbytes_1_T_1 ? phv_data_42 : _GEN_1170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1172 = 8'h2b == _match_key_qbytes_1_T_1 ? phv_data_43 : _GEN_1171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1173 = 8'h2c == _match_key_qbytes_1_T_1 ? phv_data_44 : _GEN_1172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1174 = 8'h2d == _match_key_qbytes_1_T_1 ? phv_data_45 : _GEN_1173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1175 = 8'h2e == _match_key_qbytes_1_T_1 ? phv_data_46 : _GEN_1174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1176 = 8'h2f == _match_key_qbytes_1_T_1 ? phv_data_47 : _GEN_1175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1177 = 8'h30 == _match_key_qbytes_1_T_1 ? phv_data_48 : _GEN_1176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1178 = 8'h31 == _match_key_qbytes_1_T_1 ? phv_data_49 : _GEN_1177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1179 = 8'h32 == _match_key_qbytes_1_T_1 ? phv_data_50 : _GEN_1178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1180 = 8'h33 == _match_key_qbytes_1_T_1 ? phv_data_51 : _GEN_1179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1181 = 8'h34 == _match_key_qbytes_1_T_1 ? phv_data_52 : _GEN_1180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1182 = 8'h35 == _match_key_qbytes_1_T_1 ? phv_data_53 : _GEN_1181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1183 = 8'h36 == _match_key_qbytes_1_T_1 ? phv_data_54 : _GEN_1182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1184 = 8'h37 == _match_key_qbytes_1_T_1 ? phv_data_55 : _GEN_1183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1185 = 8'h38 == _match_key_qbytes_1_T_1 ? phv_data_56 : _GEN_1184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1186 = 8'h39 == _match_key_qbytes_1_T_1 ? phv_data_57 : _GEN_1185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1187 = 8'h3a == _match_key_qbytes_1_T_1 ? phv_data_58 : _GEN_1186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1188 = 8'h3b == _match_key_qbytes_1_T_1 ? phv_data_59 : _GEN_1187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1189 = 8'h3c == _match_key_qbytes_1_T_1 ? phv_data_60 : _GEN_1188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1190 = 8'h3d == _match_key_qbytes_1_T_1 ? phv_data_61 : _GEN_1189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1191 = 8'h3e == _match_key_qbytes_1_T_1 ? phv_data_62 : _GEN_1190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1192 = 8'h3f == _match_key_qbytes_1_T_1 ? phv_data_63 : _GEN_1191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1193 = 8'h40 == _match_key_qbytes_1_T_1 ? phv_data_64 : _GEN_1192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1194 = 8'h41 == _match_key_qbytes_1_T_1 ? phv_data_65 : _GEN_1193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1195 = 8'h42 == _match_key_qbytes_1_T_1 ? phv_data_66 : _GEN_1194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1196 = 8'h43 == _match_key_qbytes_1_T_1 ? phv_data_67 : _GEN_1195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1197 = 8'h44 == _match_key_qbytes_1_T_1 ? phv_data_68 : _GEN_1196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1198 = 8'h45 == _match_key_qbytes_1_T_1 ? phv_data_69 : _GEN_1197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1199 = 8'h46 == _match_key_qbytes_1_T_1 ? phv_data_70 : _GEN_1198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1200 = 8'h47 == _match_key_qbytes_1_T_1 ? phv_data_71 : _GEN_1199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1201 = 8'h48 == _match_key_qbytes_1_T_1 ? phv_data_72 : _GEN_1200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1202 = 8'h49 == _match_key_qbytes_1_T_1 ? phv_data_73 : _GEN_1201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1203 = 8'h4a == _match_key_qbytes_1_T_1 ? phv_data_74 : _GEN_1202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1204 = 8'h4b == _match_key_qbytes_1_T_1 ? phv_data_75 : _GEN_1203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1205 = 8'h4c == _match_key_qbytes_1_T_1 ? phv_data_76 : _GEN_1204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1206 = 8'h4d == _match_key_qbytes_1_T_1 ? phv_data_77 : _GEN_1205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1207 = 8'h4e == _match_key_qbytes_1_T_1 ? phv_data_78 : _GEN_1206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1208 = 8'h4f == _match_key_qbytes_1_T_1 ? phv_data_79 : _GEN_1207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1209 = 8'h50 == _match_key_qbytes_1_T_1 ? phv_data_80 : _GEN_1208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1210 = 8'h51 == _match_key_qbytes_1_T_1 ? phv_data_81 : _GEN_1209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1211 = 8'h52 == _match_key_qbytes_1_T_1 ? phv_data_82 : _GEN_1210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1212 = 8'h53 == _match_key_qbytes_1_T_1 ? phv_data_83 : _GEN_1211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1213 = 8'h54 == _match_key_qbytes_1_T_1 ? phv_data_84 : _GEN_1212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1214 = 8'h55 == _match_key_qbytes_1_T_1 ? phv_data_85 : _GEN_1213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1215 = 8'h56 == _match_key_qbytes_1_T_1 ? phv_data_86 : _GEN_1214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1216 = 8'h57 == _match_key_qbytes_1_T_1 ? phv_data_87 : _GEN_1215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1217 = 8'h58 == _match_key_qbytes_1_T_1 ? phv_data_88 : _GEN_1216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1218 = 8'h59 == _match_key_qbytes_1_T_1 ? phv_data_89 : _GEN_1217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1219 = 8'h5a == _match_key_qbytes_1_T_1 ? phv_data_90 : _GEN_1218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1220 = 8'h5b == _match_key_qbytes_1_T_1 ? phv_data_91 : _GEN_1219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1221 = 8'h5c == _match_key_qbytes_1_T_1 ? phv_data_92 : _GEN_1220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1222 = 8'h5d == _match_key_qbytes_1_T_1 ? phv_data_93 : _GEN_1221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1223 = 8'h5e == _match_key_qbytes_1_T_1 ? phv_data_94 : _GEN_1222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1224 = 8'h5f == _match_key_qbytes_1_T_1 ? phv_data_95 : _GEN_1223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1225 = 8'h60 == _match_key_qbytes_1_T_1 ? phv_data_96 : _GEN_1224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1226 = 8'h61 == _match_key_qbytes_1_T_1 ? phv_data_97 : _GEN_1225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1227 = 8'h62 == _match_key_qbytes_1_T_1 ? phv_data_98 : _GEN_1226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1228 = 8'h63 == _match_key_qbytes_1_T_1 ? phv_data_99 : _GEN_1227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1229 = 8'h64 == _match_key_qbytes_1_T_1 ? phv_data_100 : _GEN_1228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1230 = 8'h65 == _match_key_qbytes_1_T_1 ? phv_data_101 : _GEN_1229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1231 = 8'h66 == _match_key_qbytes_1_T_1 ? phv_data_102 : _GEN_1230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1232 = 8'h67 == _match_key_qbytes_1_T_1 ? phv_data_103 : _GEN_1231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1233 = 8'h68 == _match_key_qbytes_1_T_1 ? phv_data_104 : _GEN_1232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1234 = 8'h69 == _match_key_qbytes_1_T_1 ? phv_data_105 : _GEN_1233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1235 = 8'h6a == _match_key_qbytes_1_T_1 ? phv_data_106 : _GEN_1234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1236 = 8'h6b == _match_key_qbytes_1_T_1 ? phv_data_107 : _GEN_1235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1237 = 8'h6c == _match_key_qbytes_1_T_1 ? phv_data_108 : _GEN_1236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1238 = 8'h6d == _match_key_qbytes_1_T_1 ? phv_data_109 : _GEN_1237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1239 = 8'h6e == _match_key_qbytes_1_T_1 ? phv_data_110 : _GEN_1238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1240 = 8'h6f == _match_key_qbytes_1_T_1 ? phv_data_111 : _GEN_1239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1241 = 8'h70 == _match_key_qbytes_1_T_1 ? phv_data_112 : _GEN_1240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1242 = 8'h71 == _match_key_qbytes_1_T_1 ? phv_data_113 : _GEN_1241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1243 = 8'h72 == _match_key_qbytes_1_T_1 ? phv_data_114 : _GEN_1242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1244 = 8'h73 == _match_key_qbytes_1_T_1 ? phv_data_115 : _GEN_1243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1245 = 8'h74 == _match_key_qbytes_1_T_1 ? phv_data_116 : _GEN_1244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1246 = 8'h75 == _match_key_qbytes_1_T_1 ? phv_data_117 : _GEN_1245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1247 = 8'h76 == _match_key_qbytes_1_T_1 ? phv_data_118 : _GEN_1246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1248 = 8'h77 == _match_key_qbytes_1_T_1 ? phv_data_119 : _GEN_1247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1249 = 8'h78 == _match_key_qbytes_1_T_1 ? phv_data_120 : _GEN_1248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1250 = 8'h79 == _match_key_qbytes_1_T_1 ? phv_data_121 : _GEN_1249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1251 = 8'h7a == _match_key_qbytes_1_T_1 ? phv_data_122 : _GEN_1250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1252 = 8'h7b == _match_key_qbytes_1_T_1 ? phv_data_123 : _GEN_1251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1253 = 8'h7c == _match_key_qbytes_1_T_1 ? phv_data_124 : _GEN_1252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1254 = 8'h7d == _match_key_qbytes_1_T_1 ? phv_data_125 : _GEN_1253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1255 = 8'h7e == _match_key_qbytes_1_T_1 ? phv_data_126 : _GEN_1254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1256 = 8'h7f == _match_key_qbytes_1_T_1 ? phv_data_127 : _GEN_1255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1257 = 8'h80 == _match_key_qbytes_1_T_1 ? phv_data_128 : _GEN_1256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1258 = 8'h81 == _match_key_qbytes_1_T_1 ? phv_data_129 : _GEN_1257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1259 = 8'h82 == _match_key_qbytes_1_T_1 ? phv_data_130 : _GEN_1258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1260 = 8'h83 == _match_key_qbytes_1_T_1 ? phv_data_131 : _GEN_1259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1261 = 8'h84 == _match_key_qbytes_1_T_1 ? phv_data_132 : _GEN_1260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1262 = 8'h85 == _match_key_qbytes_1_T_1 ? phv_data_133 : _GEN_1261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1263 = 8'h86 == _match_key_qbytes_1_T_1 ? phv_data_134 : _GEN_1262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1264 = 8'h87 == _match_key_qbytes_1_T_1 ? phv_data_135 : _GEN_1263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1265 = 8'h88 == _match_key_qbytes_1_T_1 ? phv_data_136 : _GEN_1264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1266 = 8'h89 == _match_key_qbytes_1_T_1 ? phv_data_137 : _GEN_1265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1267 = 8'h8a == _match_key_qbytes_1_T_1 ? phv_data_138 : _GEN_1266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1268 = 8'h8b == _match_key_qbytes_1_T_1 ? phv_data_139 : _GEN_1267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1269 = 8'h8c == _match_key_qbytes_1_T_1 ? phv_data_140 : _GEN_1268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1270 = 8'h8d == _match_key_qbytes_1_T_1 ? phv_data_141 : _GEN_1269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1271 = 8'h8e == _match_key_qbytes_1_T_1 ? phv_data_142 : _GEN_1270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1272 = 8'h8f == _match_key_qbytes_1_T_1 ? phv_data_143 : _GEN_1271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1273 = 8'h90 == _match_key_qbytes_1_T_1 ? phv_data_144 : _GEN_1272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1274 = 8'h91 == _match_key_qbytes_1_T_1 ? phv_data_145 : _GEN_1273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1275 = 8'h92 == _match_key_qbytes_1_T_1 ? phv_data_146 : _GEN_1274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1276 = 8'h93 == _match_key_qbytes_1_T_1 ? phv_data_147 : _GEN_1275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1277 = 8'h94 == _match_key_qbytes_1_T_1 ? phv_data_148 : _GEN_1276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1278 = 8'h95 == _match_key_qbytes_1_T_1 ? phv_data_149 : _GEN_1277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1279 = 8'h96 == _match_key_qbytes_1_T_1 ? phv_data_150 : _GEN_1278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1280 = 8'h97 == _match_key_qbytes_1_T_1 ? phv_data_151 : _GEN_1279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1281 = 8'h98 == _match_key_qbytes_1_T_1 ? phv_data_152 : _GEN_1280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1282 = 8'h99 == _match_key_qbytes_1_T_1 ? phv_data_153 : _GEN_1281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1283 = 8'h9a == _match_key_qbytes_1_T_1 ? phv_data_154 : _GEN_1282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1284 = 8'h9b == _match_key_qbytes_1_T_1 ? phv_data_155 : _GEN_1283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1285 = 8'h9c == _match_key_qbytes_1_T_1 ? phv_data_156 : _GEN_1284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1286 = 8'h9d == _match_key_qbytes_1_T_1 ? phv_data_157 : _GEN_1285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1287 = 8'h9e == _match_key_qbytes_1_T_1 ? phv_data_158 : _GEN_1286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1288 = 8'h9f == _match_key_qbytes_1_T_1 ? phv_data_159 : _GEN_1287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [31:0] _match_key_qbytes_1_T_3 = {_GEN_1128,_GEN_1288,_GEN_808,_GEN_968}; // @[Cat.scala 30:58]
  wire [31:0] match_key_qbytes_1 = local_offset_1 < end_offset ? _match_key_qbytes_1_T_3 : 32'h0; // @[matcher.scala 88:54 matcher.scala 89:45 matcher.scala 97:45]
  wire [7:0] local_offset_2 = 8'h8 + read_key_offset; // @[matcher.scala 87:77]
  wire [5:0] match_key_qbytes_2_hi = local_offset_2[7:2]; // @[matcher.scala 91:54]
  wire [7:0] _match_key_qbytes_2_T = {match_key_qbytes_2_hi,2'h3}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_2_T_1 = {match_key_qbytes_2_hi,2'h2}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_2_T_2 = {match_key_qbytes_2_hi,2'h1}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_1291 = 8'h1 == _match_key_qbytes_2_T_2 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1292 = 8'h2 == _match_key_qbytes_2_T_2 ? phv_data_2 : _GEN_1291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1293 = 8'h3 == _match_key_qbytes_2_T_2 ? phv_data_3 : _GEN_1292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1294 = 8'h4 == _match_key_qbytes_2_T_2 ? phv_data_4 : _GEN_1293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1295 = 8'h5 == _match_key_qbytes_2_T_2 ? phv_data_5 : _GEN_1294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1296 = 8'h6 == _match_key_qbytes_2_T_2 ? phv_data_6 : _GEN_1295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1297 = 8'h7 == _match_key_qbytes_2_T_2 ? phv_data_7 : _GEN_1296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1298 = 8'h8 == _match_key_qbytes_2_T_2 ? phv_data_8 : _GEN_1297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1299 = 8'h9 == _match_key_qbytes_2_T_2 ? phv_data_9 : _GEN_1298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1300 = 8'ha == _match_key_qbytes_2_T_2 ? phv_data_10 : _GEN_1299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1301 = 8'hb == _match_key_qbytes_2_T_2 ? phv_data_11 : _GEN_1300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1302 = 8'hc == _match_key_qbytes_2_T_2 ? phv_data_12 : _GEN_1301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1303 = 8'hd == _match_key_qbytes_2_T_2 ? phv_data_13 : _GEN_1302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1304 = 8'he == _match_key_qbytes_2_T_2 ? phv_data_14 : _GEN_1303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1305 = 8'hf == _match_key_qbytes_2_T_2 ? phv_data_15 : _GEN_1304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1306 = 8'h10 == _match_key_qbytes_2_T_2 ? phv_data_16 : _GEN_1305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1307 = 8'h11 == _match_key_qbytes_2_T_2 ? phv_data_17 : _GEN_1306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1308 = 8'h12 == _match_key_qbytes_2_T_2 ? phv_data_18 : _GEN_1307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1309 = 8'h13 == _match_key_qbytes_2_T_2 ? phv_data_19 : _GEN_1308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1310 = 8'h14 == _match_key_qbytes_2_T_2 ? phv_data_20 : _GEN_1309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1311 = 8'h15 == _match_key_qbytes_2_T_2 ? phv_data_21 : _GEN_1310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1312 = 8'h16 == _match_key_qbytes_2_T_2 ? phv_data_22 : _GEN_1311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1313 = 8'h17 == _match_key_qbytes_2_T_2 ? phv_data_23 : _GEN_1312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1314 = 8'h18 == _match_key_qbytes_2_T_2 ? phv_data_24 : _GEN_1313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1315 = 8'h19 == _match_key_qbytes_2_T_2 ? phv_data_25 : _GEN_1314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1316 = 8'h1a == _match_key_qbytes_2_T_2 ? phv_data_26 : _GEN_1315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1317 = 8'h1b == _match_key_qbytes_2_T_2 ? phv_data_27 : _GEN_1316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1318 = 8'h1c == _match_key_qbytes_2_T_2 ? phv_data_28 : _GEN_1317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1319 = 8'h1d == _match_key_qbytes_2_T_2 ? phv_data_29 : _GEN_1318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1320 = 8'h1e == _match_key_qbytes_2_T_2 ? phv_data_30 : _GEN_1319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1321 = 8'h1f == _match_key_qbytes_2_T_2 ? phv_data_31 : _GEN_1320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1322 = 8'h20 == _match_key_qbytes_2_T_2 ? phv_data_32 : _GEN_1321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1323 = 8'h21 == _match_key_qbytes_2_T_2 ? phv_data_33 : _GEN_1322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1324 = 8'h22 == _match_key_qbytes_2_T_2 ? phv_data_34 : _GEN_1323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1325 = 8'h23 == _match_key_qbytes_2_T_2 ? phv_data_35 : _GEN_1324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1326 = 8'h24 == _match_key_qbytes_2_T_2 ? phv_data_36 : _GEN_1325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1327 = 8'h25 == _match_key_qbytes_2_T_2 ? phv_data_37 : _GEN_1326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1328 = 8'h26 == _match_key_qbytes_2_T_2 ? phv_data_38 : _GEN_1327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1329 = 8'h27 == _match_key_qbytes_2_T_2 ? phv_data_39 : _GEN_1328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1330 = 8'h28 == _match_key_qbytes_2_T_2 ? phv_data_40 : _GEN_1329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1331 = 8'h29 == _match_key_qbytes_2_T_2 ? phv_data_41 : _GEN_1330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1332 = 8'h2a == _match_key_qbytes_2_T_2 ? phv_data_42 : _GEN_1331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1333 = 8'h2b == _match_key_qbytes_2_T_2 ? phv_data_43 : _GEN_1332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1334 = 8'h2c == _match_key_qbytes_2_T_2 ? phv_data_44 : _GEN_1333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1335 = 8'h2d == _match_key_qbytes_2_T_2 ? phv_data_45 : _GEN_1334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1336 = 8'h2e == _match_key_qbytes_2_T_2 ? phv_data_46 : _GEN_1335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1337 = 8'h2f == _match_key_qbytes_2_T_2 ? phv_data_47 : _GEN_1336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1338 = 8'h30 == _match_key_qbytes_2_T_2 ? phv_data_48 : _GEN_1337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1339 = 8'h31 == _match_key_qbytes_2_T_2 ? phv_data_49 : _GEN_1338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1340 = 8'h32 == _match_key_qbytes_2_T_2 ? phv_data_50 : _GEN_1339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1341 = 8'h33 == _match_key_qbytes_2_T_2 ? phv_data_51 : _GEN_1340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1342 = 8'h34 == _match_key_qbytes_2_T_2 ? phv_data_52 : _GEN_1341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1343 = 8'h35 == _match_key_qbytes_2_T_2 ? phv_data_53 : _GEN_1342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1344 = 8'h36 == _match_key_qbytes_2_T_2 ? phv_data_54 : _GEN_1343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1345 = 8'h37 == _match_key_qbytes_2_T_2 ? phv_data_55 : _GEN_1344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1346 = 8'h38 == _match_key_qbytes_2_T_2 ? phv_data_56 : _GEN_1345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1347 = 8'h39 == _match_key_qbytes_2_T_2 ? phv_data_57 : _GEN_1346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1348 = 8'h3a == _match_key_qbytes_2_T_2 ? phv_data_58 : _GEN_1347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1349 = 8'h3b == _match_key_qbytes_2_T_2 ? phv_data_59 : _GEN_1348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1350 = 8'h3c == _match_key_qbytes_2_T_2 ? phv_data_60 : _GEN_1349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1351 = 8'h3d == _match_key_qbytes_2_T_2 ? phv_data_61 : _GEN_1350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1352 = 8'h3e == _match_key_qbytes_2_T_2 ? phv_data_62 : _GEN_1351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1353 = 8'h3f == _match_key_qbytes_2_T_2 ? phv_data_63 : _GEN_1352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1354 = 8'h40 == _match_key_qbytes_2_T_2 ? phv_data_64 : _GEN_1353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1355 = 8'h41 == _match_key_qbytes_2_T_2 ? phv_data_65 : _GEN_1354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1356 = 8'h42 == _match_key_qbytes_2_T_2 ? phv_data_66 : _GEN_1355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1357 = 8'h43 == _match_key_qbytes_2_T_2 ? phv_data_67 : _GEN_1356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1358 = 8'h44 == _match_key_qbytes_2_T_2 ? phv_data_68 : _GEN_1357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1359 = 8'h45 == _match_key_qbytes_2_T_2 ? phv_data_69 : _GEN_1358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1360 = 8'h46 == _match_key_qbytes_2_T_2 ? phv_data_70 : _GEN_1359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1361 = 8'h47 == _match_key_qbytes_2_T_2 ? phv_data_71 : _GEN_1360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1362 = 8'h48 == _match_key_qbytes_2_T_2 ? phv_data_72 : _GEN_1361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1363 = 8'h49 == _match_key_qbytes_2_T_2 ? phv_data_73 : _GEN_1362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1364 = 8'h4a == _match_key_qbytes_2_T_2 ? phv_data_74 : _GEN_1363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1365 = 8'h4b == _match_key_qbytes_2_T_2 ? phv_data_75 : _GEN_1364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1366 = 8'h4c == _match_key_qbytes_2_T_2 ? phv_data_76 : _GEN_1365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1367 = 8'h4d == _match_key_qbytes_2_T_2 ? phv_data_77 : _GEN_1366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1368 = 8'h4e == _match_key_qbytes_2_T_2 ? phv_data_78 : _GEN_1367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1369 = 8'h4f == _match_key_qbytes_2_T_2 ? phv_data_79 : _GEN_1368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1370 = 8'h50 == _match_key_qbytes_2_T_2 ? phv_data_80 : _GEN_1369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1371 = 8'h51 == _match_key_qbytes_2_T_2 ? phv_data_81 : _GEN_1370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1372 = 8'h52 == _match_key_qbytes_2_T_2 ? phv_data_82 : _GEN_1371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1373 = 8'h53 == _match_key_qbytes_2_T_2 ? phv_data_83 : _GEN_1372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1374 = 8'h54 == _match_key_qbytes_2_T_2 ? phv_data_84 : _GEN_1373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1375 = 8'h55 == _match_key_qbytes_2_T_2 ? phv_data_85 : _GEN_1374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1376 = 8'h56 == _match_key_qbytes_2_T_2 ? phv_data_86 : _GEN_1375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1377 = 8'h57 == _match_key_qbytes_2_T_2 ? phv_data_87 : _GEN_1376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1378 = 8'h58 == _match_key_qbytes_2_T_2 ? phv_data_88 : _GEN_1377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1379 = 8'h59 == _match_key_qbytes_2_T_2 ? phv_data_89 : _GEN_1378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1380 = 8'h5a == _match_key_qbytes_2_T_2 ? phv_data_90 : _GEN_1379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1381 = 8'h5b == _match_key_qbytes_2_T_2 ? phv_data_91 : _GEN_1380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1382 = 8'h5c == _match_key_qbytes_2_T_2 ? phv_data_92 : _GEN_1381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1383 = 8'h5d == _match_key_qbytes_2_T_2 ? phv_data_93 : _GEN_1382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1384 = 8'h5e == _match_key_qbytes_2_T_2 ? phv_data_94 : _GEN_1383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1385 = 8'h5f == _match_key_qbytes_2_T_2 ? phv_data_95 : _GEN_1384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1386 = 8'h60 == _match_key_qbytes_2_T_2 ? phv_data_96 : _GEN_1385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1387 = 8'h61 == _match_key_qbytes_2_T_2 ? phv_data_97 : _GEN_1386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1388 = 8'h62 == _match_key_qbytes_2_T_2 ? phv_data_98 : _GEN_1387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1389 = 8'h63 == _match_key_qbytes_2_T_2 ? phv_data_99 : _GEN_1388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1390 = 8'h64 == _match_key_qbytes_2_T_2 ? phv_data_100 : _GEN_1389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1391 = 8'h65 == _match_key_qbytes_2_T_2 ? phv_data_101 : _GEN_1390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1392 = 8'h66 == _match_key_qbytes_2_T_2 ? phv_data_102 : _GEN_1391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1393 = 8'h67 == _match_key_qbytes_2_T_2 ? phv_data_103 : _GEN_1392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1394 = 8'h68 == _match_key_qbytes_2_T_2 ? phv_data_104 : _GEN_1393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1395 = 8'h69 == _match_key_qbytes_2_T_2 ? phv_data_105 : _GEN_1394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1396 = 8'h6a == _match_key_qbytes_2_T_2 ? phv_data_106 : _GEN_1395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1397 = 8'h6b == _match_key_qbytes_2_T_2 ? phv_data_107 : _GEN_1396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1398 = 8'h6c == _match_key_qbytes_2_T_2 ? phv_data_108 : _GEN_1397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1399 = 8'h6d == _match_key_qbytes_2_T_2 ? phv_data_109 : _GEN_1398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1400 = 8'h6e == _match_key_qbytes_2_T_2 ? phv_data_110 : _GEN_1399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1401 = 8'h6f == _match_key_qbytes_2_T_2 ? phv_data_111 : _GEN_1400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1402 = 8'h70 == _match_key_qbytes_2_T_2 ? phv_data_112 : _GEN_1401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1403 = 8'h71 == _match_key_qbytes_2_T_2 ? phv_data_113 : _GEN_1402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1404 = 8'h72 == _match_key_qbytes_2_T_2 ? phv_data_114 : _GEN_1403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1405 = 8'h73 == _match_key_qbytes_2_T_2 ? phv_data_115 : _GEN_1404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1406 = 8'h74 == _match_key_qbytes_2_T_2 ? phv_data_116 : _GEN_1405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1407 = 8'h75 == _match_key_qbytes_2_T_2 ? phv_data_117 : _GEN_1406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1408 = 8'h76 == _match_key_qbytes_2_T_2 ? phv_data_118 : _GEN_1407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1409 = 8'h77 == _match_key_qbytes_2_T_2 ? phv_data_119 : _GEN_1408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1410 = 8'h78 == _match_key_qbytes_2_T_2 ? phv_data_120 : _GEN_1409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1411 = 8'h79 == _match_key_qbytes_2_T_2 ? phv_data_121 : _GEN_1410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1412 = 8'h7a == _match_key_qbytes_2_T_2 ? phv_data_122 : _GEN_1411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1413 = 8'h7b == _match_key_qbytes_2_T_2 ? phv_data_123 : _GEN_1412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1414 = 8'h7c == _match_key_qbytes_2_T_2 ? phv_data_124 : _GEN_1413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1415 = 8'h7d == _match_key_qbytes_2_T_2 ? phv_data_125 : _GEN_1414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1416 = 8'h7e == _match_key_qbytes_2_T_2 ? phv_data_126 : _GEN_1415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1417 = 8'h7f == _match_key_qbytes_2_T_2 ? phv_data_127 : _GEN_1416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1418 = 8'h80 == _match_key_qbytes_2_T_2 ? phv_data_128 : _GEN_1417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1419 = 8'h81 == _match_key_qbytes_2_T_2 ? phv_data_129 : _GEN_1418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1420 = 8'h82 == _match_key_qbytes_2_T_2 ? phv_data_130 : _GEN_1419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1421 = 8'h83 == _match_key_qbytes_2_T_2 ? phv_data_131 : _GEN_1420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1422 = 8'h84 == _match_key_qbytes_2_T_2 ? phv_data_132 : _GEN_1421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1423 = 8'h85 == _match_key_qbytes_2_T_2 ? phv_data_133 : _GEN_1422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1424 = 8'h86 == _match_key_qbytes_2_T_2 ? phv_data_134 : _GEN_1423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1425 = 8'h87 == _match_key_qbytes_2_T_2 ? phv_data_135 : _GEN_1424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1426 = 8'h88 == _match_key_qbytes_2_T_2 ? phv_data_136 : _GEN_1425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1427 = 8'h89 == _match_key_qbytes_2_T_2 ? phv_data_137 : _GEN_1426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1428 = 8'h8a == _match_key_qbytes_2_T_2 ? phv_data_138 : _GEN_1427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1429 = 8'h8b == _match_key_qbytes_2_T_2 ? phv_data_139 : _GEN_1428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1430 = 8'h8c == _match_key_qbytes_2_T_2 ? phv_data_140 : _GEN_1429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1431 = 8'h8d == _match_key_qbytes_2_T_2 ? phv_data_141 : _GEN_1430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1432 = 8'h8e == _match_key_qbytes_2_T_2 ? phv_data_142 : _GEN_1431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1433 = 8'h8f == _match_key_qbytes_2_T_2 ? phv_data_143 : _GEN_1432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1434 = 8'h90 == _match_key_qbytes_2_T_2 ? phv_data_144 : _GEN_1433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1435 = 8'h91 == _match_key_qbytes_2_T_2 ? phv_data_145 : _GEN_1434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1436 = 8'h92 == _match_key_qbytes_2_T_2 ? phv_data_146 : _GEN_1435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1437 = 8'h93 == _match_key_qbytes_2_T_2 ? phv_data_147 : _GEN_1436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1438 = 8'h94 == _match_key_qbytes_2_T_2 ? phv_data_148 : _GEN_1437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1439 = 8'h95 == _match_key_qbytes_2_T_2 ? phv_data_149 : _GEN_1438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1440 = 8'h96 == _match_key_qbytes_2_T_2 ? phv_data_150 : _GEN_1439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1441 = 8'h97 == _match_key_qbytes_2_T_2 ? phv_data_151 : _GEN_1440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1442 = 8'h98 == _match_key_qbytes_2_T_2 ? phv_data_152 : _GEN_1441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1443 = 8'h99 == _match_key_qbytes_2_T_2 ? phv_data_153 : _GEN_1442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1444 = 8'h9a == _match_key_qbytes_2_T_2 ? phv_data_154 : _GEN_1443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1445 = 8'h9b == _match_key_qbytes_2_T_2 ? phv_data_155 : _GEN_1444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1446 = 8'h9c == _match_key_qbytes_2_T_2 ? phv_data_156 : _GEN_1445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1447 = 8'h9d == _match_key_qbytes_2_T_2 ? phv_data_157 : _GEN_1446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1448 = 8'h9e == _match_key_qbytes_2_T_2 ? phv_data_158 : _GEN_1447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1449 = 8'h9f == _match_key_qbytes_2_T_2 ? phv_data_159 : _GEN_1448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1451 = 8'h1 == local_offset_2 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1452 = 8'h2 == local_offset_2 ? phv_data_2 : _GEN_1451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1453 = 8'h3 == local_offset_2 ? phv_data_3 : _GEN_1452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1454 = 8'h4 == local_offset_2 ? phv_data_4 : _GEN_1453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1455 = 8'h5 == local_offset_2 ? phv_data_5 : _GEN_1454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1456 = 8'h6 == local_offset_2 ? phv_data_6 : _GEN_1455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1457 = 8'h7 == local_offset_2 ? phv_data_7 : _GEN_1456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1458 = 8'h8 == local_offset_2 ? phv_data_8 : _GEN_1457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1459 = 8'h9 == local_offset_2 ? phv_data_9 : _GEN_1458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1460 = 8'ha == local_offset_2 ? phv_data_10 : _GEN_1459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1461 = 8'hb == local_offset_2 ? phv_data_11 : _GEN_1460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1462 = 8'hc == local_offset_2 ? phv_data_12 : _GEN_1461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1463 = 8'hd == local_offset_2 ? phv_data_13 : _GEN_1462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1464 = 8'he == local_offset_2 ? phv_data_14 : _GEN_1463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1465 = 8'hf == local_offset_2 ? phv_data_15 : _GEN_1464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1466 = 8'h10 == local_offset_2 ? phv_data_16 : _GEN_1465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1467 = 8'h11 == local_offset_2 ? phv_data_17 : _GEN_1466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1468 = 8'h12 == local_offset_2 ? phv_data_18 : _GEN_1467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1469 = 8'h13 == local_offset_2 ? phv_data_19 : _GEN_1468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1470 = 8'h14 == local_offset_2 ? phv_data_20 : _GEN_1469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1471 = 8'h15 == local_offset_2 ? phv_data_21 : _GEN_1470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1472 = 8'h16 == local_offset_2 ? phv_data_22 : _GEN_1471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1473 = 8'h17 == local_offset_2 ? phv_data_23 : _GEN_1472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1474 = 8'h18 == local_offset_2 ? phv_data_24 : _GEN_1473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1475 = 8'h19 == local_offset_2 ? phv_data_25 : _GEN_1474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1476 = 8'h1a == local_offset_2 ? phv_data_26 : _GEN_1475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1477 = 8'h1b == local_offset_2 ? phv_data_27 : _GEN_1476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1478 = 8'h1c == local_offset_2 ? phv_data_28 : _GEN_1477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1479 = 8'h1d == local_offset_2 ? phv_data_29 : _GEN_1478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1480 = 8'h1e == local_offset_2 ? phv_data_30 : _GEN_1479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1481 = 8'h1f == local_offset_2 ? phv_data_31 : _GEN_1480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1482 = 8'h20 == local_offset_2 ? phv_data_32 : _GEN_1481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1483 = 8'h21 == local_offset_2 ? phv_data_33 : _GEN_1482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1484 = 8'h22 == local_offset_2 ? phv_data_34 : _GEN_1483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1485 = 8'h23 == local_offset_2 ? phv_data_35 : _GEN_1484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1486 = 8'h24 == local_offset_2 ? phv_data_36 : _GEN_1485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1487 = 8'h25 == local_offset_2 ? phv_data_37 : _GEN_1486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1488 = 8'h26 == local_offset_2 ? phv_data_38 : _GEN_1487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1489 = 8'h27 == local_offset_2 ? phv_data_39 : _GEN_1488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1490 = 8'h28 == local_offset_2 ? phv_data_40 : _GEN_1489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1491 = 8'h29 == local_offset_2 ? phv_data_41 : _GEN_1490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1492 = 8'h2a == local_offset_2 ? phv_data_42 : _GEN_1491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1493 = 8'h2b == local_offset_2 ? phv_data_43 : _GEN_1492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1494 = 8'h2c == local_offset_2 ? phv_data_44 : _GEN_1493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1495 = 8'h2d == local_offset_2 ? phv_data_45 : _GEN_1494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1496 = 8'h2e == local_offset_2 ? phv_data_46 : _GEN_1495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1497 = 8'h2f == local_offset_2 ? phv_data_47 : _GEN_1496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1498 = 8'h30 == local_offset_2 ? phv_data_48 : _GEN_1497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1499 = 8'h31 == local_offset_2 ? phv_data_49 : _GEN_1498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1500 = 8'h32 == local_offset_2 ? phv_data_50 : _GEN_1499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1501 = 8'h33 == local_offset_2 ? phv_data_51 : _GEN_1500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1502 = 8'h34 == local_offset_2 ? phv_data_52 : _GEN_1501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1503 = 8'h35 == local_offset_2 ? phv_data_53 : _GEN_1502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1504 = 8'h36 == local_offset_2 ? phv_data_54 : _GEN_1503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1505 = 8'h37 == local_offset_2 ? phv_data_55 : _GEN_1504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1506 = 8'h38 == local_offset_2 ? phv_data_56 : _GEN_1505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1507 = 8'h39 == local_offset_2 ? phv_data_57 : _GEN_1506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1508 = 8'h3a == local_offset_2 ? phv_data_58 : _GEN_1507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1509 = 8'h3b == local_offset_2 ? phv_data_59 : _GEN_1508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1510 = 8'h3c == local_offset_2 ? phv_data_60 : _GEN_1509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1511 = 8'h3d == local_offset_2 ? phv_data_61 : _GEN_1510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1512 = 8'h3e == local_offset_2 ? phv_data_62 : _GEN_1511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1513 = 8'h3f == local_offset_2 ? phv_data_63 : _GEN_1512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1514 = 8'h40 == local_offset_2 ? phv_data_64 : _GEN_1513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1515 = 8'h41 == local_offset_2 ? phv_data_65 : _GEN_1514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1516 = 8'h42 == local_offset_2 ? phv_data_66 : _GEN_1515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1517 = 8'h43 == local_offset_2 ? phv_data_67 : _GEN_1516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1518 = 8'h44 == local_offset_2 ? phv_data_68 : _GEN_1517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1519 = 8'h45 == local_offset_2 ? phv_data_69 : _GEN_1518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1520 = 8'h46 == local_offset_2 ? phv_data_70 : _GEN_1519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1521 = 8'h47 == local_offset_2 ? phv_data_71 : _GEN_1520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1522 = 8'h48 == local_offset_2 ? phv_data_72 : _GEN_1521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1523 = 8'h49 == local_offset_2 ? phv_data_73 : _GEN_1522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1524 = 8'h4a == local_offset_2 ? phv_data_74 : _GEN_1523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1525 = 8'h4b == local_offset_2 ? phv_data_75 : _GEN_1524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1526 = 8'h4c == local_offset_2 ? phv_data_76 : _GEN_1525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1527 = 8'h4d == local_offset_2 ? phv_data_77 : _GEN_1526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1528 = 8'h4e == local_offset_2 ? phv_data_78 : _GEN_1527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1529 = 8'h4f == local_offset_2 ? phv_data_79 : _GEN_1528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1530 = 8'h50 == local_offset_2 ? phv_data_80 : _GEN_1529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1531 = 8'h51 == local_offset_2 ? phv_data_81 : _GEN_1530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1532 = 8'h52 == local_offset_2 ? phv_data_82 : _GEN_1531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1533 = 8'h53 == local_offset_2 ? phv_data_83 : _GEN_1532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1534 = 8'h54 == local_offset_2 ? phv_data_84 : _GEN_1533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1535 = 8'h55 == local_offset_2 ? phv_data_85 : _GEN_1534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1536 = 8'h56 == local_offset_2 ? phv_data_86 : _GEN_1535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1537 = 8'h57 == local_offset_2 ? phv_data_87 : _GEN_1536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1538 = 8'h58 == local_offset_2 ? phv_data_88 : _GEN_1537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1539 = 8'h59 == local_offset_2 ? phv_data_89 : _GEN_1538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1540 = 8'h5a == local_offset_2 ? phv_data_90 : _GEN_1539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1541 = 8'h5b == local_offset_2 ? phv_data_91 : _GEN_1540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1542 = 8'h5c == local_offset_2 ? phv_data_92 : _GEN_1541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1543 = 8'h5d == local_offset_2 ? phv_data_93 : _GEN_1542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1544 = 8'h5e == local_offset_2 ? phv_data_94 : _GEN_1543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1545 = 8'h5f == local_offset_2 ? phv_data_95 : _GEN_1544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1546 = 8'h60 == local_offset_2 ? phv_data_96 : _GEN_1545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1547 = 8'h61 == local_offset_2 ? phv_data_97 : _GEN_1546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1548 = 8'h62 == local_offset_2 ? phv_data_98 : _GEN_1547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1549 = 8'h63 == local_offset_2 ? phv_data_99 : _GEN_1548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1550 = 8'h64 == local_offset_2 ? phv_data_100 : _GEN_1549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1551 = 8'h65 == local_offset_2 ? phv_data_101 : _GEN_1550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1552 = 8'h66 == local_offset_2 ? phv_data_102 : _GEN_1551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1553 = 8'h67 == local_offset_2 ? phv_data_103 : _GEN_1552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1554 = 8'h68 == local_offset_2 ? phv_data_104 : _GEN_1553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1555 = 8'h69 == local_offset_2 ? phv_data_105 : _GEN_1554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1556 = 8'h6a == local_offset_2 ? phv_data_106 : _GEN_1555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1557 = 8'h6b == local_offset_2 ? phv_data_107 : _GEN_1556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1558 = 8'h6c == local_offset_2 ? phv_data_108 : _GEN_1557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1559 = 8'h6d == local_offset_2 ? phv_data_109 : _GEN_1558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1560 = 8'h6e == local_offset_2 ? phv_data_110 : _GEN_1559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1561 = 8'h6f == local_offset_2 ? phv_data_111 : _GEN_1560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1562 = 8'h70 == local_offset_2 ? phv_data_112 : _GEN_1561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1563 = 8'h71 == local_offset_2 ? phv_data_113 : _GEN_1562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1564 = 8'h72 == local_offset_2 ? phv_data_114 : _GEN_1563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1565 = 8'h73 == local_offset_2 ? phv_data_115 : _GEN_1564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1566 = 8'h74 == local_offset_2 ? phv_data_116 : _GEN_1565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1567 = 8'h75 == local_offset_2 ? phv_data_117 : _GEN_1566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1568 = 8'h76 == local_offset_2 ? phv_data_118 : _GEN_1567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1569 = 8'h77 == local_offset_2 ? phv_data_119 : _GEN_1568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1570 = 8'h78 == local_offset_2 ? phv_data_120 : _GEN_1569; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1571 = 8'h79 == local_offset_2 ? phv_data_121 : _GEN_1570; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1572 = 8'h7a == local_offset_2 ? phv_data_122 : _GEN_1571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1573 = 8'h7b == local_offset_2 ? phv_data_123 : _GEN_1572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1574 = 8'h7c == local_offset_2 ? phv_data_124 : _GEN_1573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1575 = 8'h7d == local_offset_2 ? phv_data_125 : _GEN_1574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1576 = 8'h7e == local_offset_2 ? phv_data_126 : _GEN_1575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1577 = 8'h7f == local_offset_2 ? phv_data_127 : _GEN_1576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1578 = 8'h80 == local_offset_2 ? phv_data_128 : _GEN_1577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1579 = 8'h81 == local_offset_2 ? phv_data_129 : _GEN_1578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1580 = 8'h82 == local_offset_2 ? phv_data_130 : _GEN_1579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1581 = 8'h83 == local_offset_2 ? phv_data_131 : _GEN_1580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1582 = 8'h84 == local_offset_2 ? phv_data_132 : _GEN_1581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1583 = 8'h85 == local_offset_2 ? phv_data_133 : _GEN_1582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1584 = 8'h86 == local_offset_2 ? phv_data_134 : _GEN_1583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1585 = 8'h87 == local_offset_2 ? phv_data_135 : _GEN_1584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1586 = 8'h88 == local_offset_2 ? phv_data_136 : _GEN_1585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1587 = 8'h89 == local_offset_2 ? phv_data_137 : _GEN_1586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1588 = 8'h8a == local_offset_2 ? phv_data_138 : _GEN_1587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1589 = 8'h8b == local_offset_2 ? phv_data_139 : _GEN_1588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1590 = 8'h8c == local_offset_2 ? phv_data_140 : _GEN_1589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1591 = 8'h8d == local_offset_2 ? phv_data_141 : _GEN_1590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1592 = 8'h8e == local_offset_2 ? phv_data_142 : _GEN_1591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1593 = 8'h8f == local_offset_2 ? phv_data_143 : _GEN_1592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1594 = 8'h90 == local_offset_2 ? phv_data_144 : _GEN_1593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1595 = 8'h91 == local_offset_2 ? phv_data_145 : _GEN_1594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1596 = 8'h92 == local_offset_2 ? phv_data_146 : _GEN_1595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1597 = 8'h93 == local_offset_2 ? phv_data_147 : _GEN_1596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1598 = 8'h94 == local_offset_2 ? phv_data_148 : _GEN_1597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1599 = 8'h95 == local_offset_2 ? phv_data_149 : _GEN_1598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1600 = 8'h96 == local_offset_2 ? phv_data_150 : _GEN_1599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1601 = 8'h97 == local_offset_2 ? phv_data_151 : _GEN_1600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1602 = 8'h98 == local_offset_2 ? phv_data_152 : _GEN_1601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1603 = 8'h99 == local_offset_2 ? phv_data_153 : _GEN_1602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1604 = 8'h9a == local_offset_2 ? phv_data_154 : _GEN_1603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1605 = 8'h9b == local_offset_2 ? phv_data_155 : _GEN_1604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1606 = 8'h9c == local_offset_2 ? phv_data_156 : _GEN_1605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1607 = 8'h9d == local_offset_2 ? phv_data_157 : _GEN_1606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1608 = 8'h9e == local_offset_2 ? phv_data_158 : _GEN_1607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1609 = 8'h9f == local_offset_2 ? phv_data_159 : _GEN_1608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1611 = 8'h1 == _match_key_qbytes_2_T ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1612 = 8'h2 == _match_key_qbytes_2_T ? phv_data_2 : _GEN_1611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1613 = 8'h3 == _match_key_qbytes_2_T ? phv_data_3 : _GEN_1612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1614 = 8'h4 == _match_key_qbytes_2_T ? phv_data_4 : _GEN_1613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1615 = 8'h5 == _match_key_qbytes_2_T ? phv_data_5 : _GEN_1614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1616 = 8'h6 == _match_key_qbytes_2_T ? phv_data_6 : _GEN_1615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1617 = 8'h7 == _match_key_qbytes_2_T ? phv_data_7 : _GEN_1616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1618 = 8'h8 == _match_key_qbytes_2_T ? phv_data_8 : _GEN_1617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1619 = 8'h9 == _match_key_qbytes_2_T ? phv_data_9 : _GEN_1618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1620 = 8'ha == _match_key_qbytes_2_T ? phv_data_10 : _GEN_1619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1621 = 8'hb == _match_key_qbytes_2_T ? phv_data_11 : _GEN_1620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1622 = 8'hc == _match_key_qbytes_2_T ? phv_data_12 : _GEN_1621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1623 = 8'hd == _match_key_qbytes_2_T ? phv_data_13 : _GEN_1622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1624 = 8'he == _match_key_qbytes_2_T ? phv_data_14 : _GEN_1623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1625 = 8'hf == _match_key_qbytes_2_T ? phv_data_15 : _GEN_1624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1626 = 8'h10 == _match_key_qbytes_2_T ? phv_data_16 : _GEN_1625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1627 = 8'h11 == _match_key_qbytes_2_T ? phv_data_17 : _GEN_1626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1628 = 8'h12 == _match_key_qbytes_2_T ? phv_data_18 : _GEN_1627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1629 = 8'h13 == _match_key_qbytes_2_T ? phv_data_19 : _GEN_1628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1630 = 8'h14 == _match_key_qbytes_2_T ? phv_data_20 : _GEN_1629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1631 = 8'h15 == _match_key_qbytes_2_T ? phv_data_21 : _GEN_1630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1632 = 8'h16 == _match_key_qbytes_2_T ? phv_data_22 : _GEN_1631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1633 = 8'h17 == _match_key_qbytes_2_T ? phv_data_23 : _GEN_1632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1634 = 8'h18 == _match_key_qbytes_2_T ? phv_data_24 : _GEN_1633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1635 = 8'h19 == _match_key_qbytes_2_T ? phv_data_25 : _GEN_1634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1636 = 8'h1a == _match_key_qbytes_2_T ? phv_data_26 : _GEN_1635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1637 = 8'h1b == _match_key_qbytes_2_T ? phv_data_27 : _GEN_1636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1638 = 8'h1c == _match_key_qbytes_2_T ? phv_data_28 : _GEN_1637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1639 = 8'h1d == _match_key_qbytes_2_T ? phv_data_29 : _GEN_1638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1640 = 8'h1e == _match_key_qbytes_2_T ? phv_data_30 : _GEN_1639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1641 = 8'h1f == _match_key_qbytes_2_T ? phv_data_31 : _GEN_1640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1642 = 8'h20 == _match_key_qbytes_2_T ? phv_data_32 : _GEN_1641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1643 = 8'h21 == _match_key_qbytes_2_T ? phv_data_33 : _GEN_1642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1644 = 8'h22 == _match_key_qbytes_2_T ? phv_data_34 : _GEN_1643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1645 = 8'h23 == _match_key_qbytes_2_T ? phv_data_35 : _GEN_1644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1646 = 8'h24 == _match_key_qbytes_2_T ? phv_data_36 : _GEN_1645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1647 = 8'h25 == _match_key_qbytes_2_T ? phv_data_37 : _GEN_1646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1648 = 8'h26 == _match_key_qbytes_2_T ? phv_data_38 : _GEN_1647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1649 = 8'h27 == _match_key_qbytes_2_T ? phv_data_39 : _GEN_1648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1650 = 8'h28 == _match_key_qbytes_2_T ? phv_data_40 : _GEN_1649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1651 = 8'h29 == _match_key_qbytes_2_T ? phv_data_41 : _GEN_1650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1652 = 8'h2a == _match_key_qbytes_2_T ? phv_data_42 : _GEN_1651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1653 = 8'h2b == _match_key_qbytes_2_T ? phv_data_43 : _GEN_1652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1654 = 8'h2c == _match_key_qbytes_2_T ? phv_data_44 : _GEN_1653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1655 = 8'h2d == _match_key_qbytes_2_T ? phv_data_45 : _GEN_1654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1656 = 8'h2e == _match_key_qbytes_2_T ? phv_data_46 : _GEN_1655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1657 = 8'h2f == _match_key_qbytes_2_T ? phv_data_47 : _GEN_1656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1658 = 8'h30 == _match_key_qbytes_2_T ? phv_data_48 : _GEN_1657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1659 = 8'h31 == _match_key_qbytes_2_T ? phv_data_49 : _GEN_1658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1660 = 8'h32 == _match_key_qbytes_2_T ? phv_data_50 : _GEN_1659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1661 = 8'h33 == _match_key_qbytes_2_T ? phv_data_51 : _GEN_1660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1662 = 8'h34 == _match_key_qbytes_2_T ? phv_data_52 : _GEN_1661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1663 = 8'h35 == _match_key_qbytes_2_T ? phv_data_53 : _GEN_1662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1664 = 8'h36 == _match_key_qbytes_2_T ? phv_data_54 : _GEN_1663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1665 = 8'h37 == _match_key_qbytes_2_T ? phv_data_55 : _GEN_1664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1666 = 8'h38 == _match_key_qbytes_2_T ? phv_data_56 : _GEN_1665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1667 = 8'h39 == _match_key_qbytes_2_T ? phv_data_57 : _GEN_1666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1668 = 8'h3a == _match_key_qbytes_2_T ? phv_data_58 : _GEN_1667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1669 = 8'h3b == _match_key_qbytes_2_T ? phv_data_59 : _GEN_1668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1670 = 8'h3c == _match_key_qbytes_2_T ? phv_data_60 : _GEN_1669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1671 = 8'h3d == _match_key_qbytes_2_T ? phv_data_61 : _GEN_1670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1672 = 8'h3e == _match_key_qbytes_2_T ? phv_data_62 : _GEN_1671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1673 = 8'h3f == _match_key_qbytes_2_T ? phv_data_63 : _GEN_1672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1674 = 8'h40 == _match_key_qbytes_2_T ? phv_data_64 : _GEN_1673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1675 = 8'h41 == _match_key_qbytes_2_T ? phv_data_65 : _GEN_1674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1676 = 8'h42 == _match_key_qbytes_2_T ? phv_data_66 : _GEN_1675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1677 = 8'h43 == _match_key_qbytes_2_T ? phv_data_67 : _GEN_1676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1678 = 8'h44 == _match_key_qbytes_2_T ? phv_data_68 : _GEN_1677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1679 = 8'h45 == _match_key_qbytes_2_T ? phv_data_69 : _GEN_1678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1680 = 8'h46 == _match_key_qbytes_2_T ? phv_data_70 : _GEN_1679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1681 = 8'h47 == _match_key_qbytes_2_T ? phv_data_71 : _GEN_1680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1682 = 8'h48 == _match_key_qbytes_2_T ? phv_data_72 : _GEN_1681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1683 = 8'h49 == _match_key_qbytes_2_T ? phv_data_73 : _GEN_1682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1684 = 8'h4a == _match_key_qbytes_2_T ? phv_data_74 : _GEN_1683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1685 = 8'h4b == _match_key_qbytes_2_T ? phv_data_75 : _GEN_1684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1686 = 8'h4c == _match_key_qbytes_2_T ? phv_data_76 : _GEN_1685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1687 = 8'h4d == _match_key_qbytes_2_T ? phv_data_77 : _GEN_1686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1688 = 8'h4e == _match_key_qbytes_2_T ? phv_data_78 : _GEN_1687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1689 = 8'h4f == _match_key_qbytes_2_T ? phv_data_79 : _GEN_1688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1690 = 8'h50 == _match_key_qbytes_2_T ? phv_data_80 : _GEN_1689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1691 = 8'h51 == _match_key_qbytes_2_T ? phv_data_81 : _GEN_1690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1692 = 8'h52 == _match_key_qbytes_2_T ? phv_data_82 : _GEN_1691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1693 = 8'h53 == _match_key_qbytes_2_T ? phv_data_83 : _GEN_1692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1694 = 8'h54 == _match_key_qbytes_2_T ? phv_data_84 : _GEN_1693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1695 = 8'h55 == _match_key_qbytes_2_T ? phv_data_85 : _GEN_1694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1696 = 8'h56 == _match_key_qbytes_2_T ? phv_data_86 : _GEN_1695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1697 = 8'h57 == _match_key_qbytes_2_T ? phv_data_87 : _GEN_1696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1698 = 8'h58 == _match_key_qbytes_2_T ? phv_data_88 : _GEN_1697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1699 = 8'h59 == _match_key_qbytes_2_T ? phv_data_89 : _GEN_1698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1700 = 8'h5a == _match_key_qbytes_2_T ? phv_data_90 : _GEN_1699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1701 = 8'h5b == _match_key_qbytes_2_T ? phv_data_91 : _GEN_1700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1702 = 8'h5c == _match_key_qbytes_2_T ? phv_data_92 : _GEN_1701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1703 = 8'h5d == _match_key_qbytes_2_T ? phv_data_93 : _GEN_1702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1704 = 8'h5e == _match_key_qbytes_2_T ? phv_data_94 : _GEN_1703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1705 = 8'h5f == _match_key_qbytes_2_T ? phv_data_95 : _GEN_1704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1706 = 8'h60 == _match_key_qbytes_2_T ? phv_data_96 : _GEN_1705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1707 = 8'h61 == _match_key_qbytes_2_T ? phv_data_97 : _GEN_1706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1708 = 8'h62 == _match_key_qbytes_2_T ? phv_data_98 : _GEN_1707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1709 = 8'h63 == _match_key_qbytes_2_T ? phv_data_99 : _GEN_1708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1710 = 8'h64 == _match_key_qbytes_2_T ? phv_data_100 : _GEN_1709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1711 = 8'h65 == _match_key_qbytes_2_T ? phv_data_101 : _GEN_1710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1712 = 8'h66 == _match_key_qbytes_2_T ? phv_data_102 : _GEN_1711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1713 = 8'h67 == _match_key_qbytes_2_T ? phv_data_103 : _GEN_1712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1714 = 8'h68 == _match_key_qbytes_2_T ? phv_data_104 : _GEN_1713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1715 = 8'h69 == _match_key_qbytes_2_T ? phv_data_105 : _GEN_1714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1716 = 8'h6a == _match_key_qbytes_2_T ? phv_data_106 : _GEN_1715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1717 = 8'h6b == _match_key_qbytes_2_T ? phv_data_107 : _GEN_1716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1718 = 8'h6c == _match_key_qbytes_2_T ? phv_data_108 : _GEN_1717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1719 = 8'h6d == _match_key_qbytes_2_T ? phv_data_109 : _GEN_1718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1720 = 8'h6e == _match_key_qbytes_2_T ? phv_data_110 : _GEN_1719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1721 = 8'h6f == _match_key_qbytes_2_T ? phv_data_111 : _GEN_1720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1722 = 8'h70 == _match_key_qbytes_2_T ? phv_data_112 : _GEN_1721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1723 = 8'h71 == _match_key_qbytes_2_T ? phv_data_113 : _GEN_1722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1724 = 8'h72 == _match_key_qbytes_2_T ? phv_data_114 : _GEN_1723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1725 = 8'h73 == _match_key_qbytes_2_T ? phv_data_115 : _GEN_1724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1726 = 8'h74 == _match_key_qbytes_2_T ? phv_data_116 : _GEN_1725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1727 = 8'h75 == _match_key_qbytes_2_T ? phv_data_117 : _GEN_1726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1728 = 8'h76 == _match_key_qbytes_2_T ? phv_data_118 : _GEN_1727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1729 = 8'h77 == _match_key_qbytes_2_T ? phv_data_119 : _GEN_1728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1730 = 8'h78 == _match_key_qbytes_2_T ? phv_data_120 : _GEN_1729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1731 = 8'h79 == _match_key_qbytes_2_T ? phv_data_121 : _GEN_1730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1732 = 8'h7a == _match_key_qbytes_2_T ? phv_data_122 : _GEN_1731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1733 = 8'h7b == _match_key_qbytes_2_T ? phv_data_123 : _GEN_1732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1734 = 8'h7c == _match_key_qbytes_2_T ? phv_data_124 : _GEN_1733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1735 = 8'h7d == _match_key_qbytes_2_T ? phv_data_125 : _GEN_1734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1736 = 8'h7e == _match_key_qbytes_2_T ? phv_data_126 : _GEN_1735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1737 = 8'h7f == _match_key_qbytes_2_T ? phv_data_127 : _GEN_1736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1738 = 8'h80 == _match_key_qbytes_2_T ? phv_data_128 : _GEN_1737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1739 = 8'h81 == _match_key_qbytes_2_T ? phv_data_129 : _GEN_1738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1740 = 8'h82 == _match_key_qbytes_2_T ? phv_data_130 : _GEN_1739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1741 = 8'h83 == _match_key_qbytes_2_T ? phv_data_131 : _GEN_1740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1742 = 8'h84 == _match_key_qbytes_2_T ? phv_data_132 : _GEN_1741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1743 = 8'h85 == _match_key_qbytes_2_T ? phv_data_133 : _GEN_1742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1744 = 8'h86 == _match_key_qbytes_2_T ? phv_data_134 : _GEN_1743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1745 = 8'h87 == _match_key_qbytes_2_T ? phv_data_135 : _GEN_1744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1746 = 8'h88 == _match_key_qbytes_2_T ? phv_data_136 : _GEN_1745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1747 = 8'h89 == _match_key_qbytes_2_T ? phv_data_137 : _GEN_1746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1748 = 8'h8a == _match_key_qbytes_2_T ? phv_data_138 : _GEN_1747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1749 = 8'h8b == _match_key_qbytes_2_T ? phv_data_139 : _GEN_1748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1750 = 8'h8c == _match_key_qbytes_2_T ? phv_data_140 : _GEN_1749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1751 = 8'h8d == _match_key_qbytes_2_T ? phv_data_141 : _GEN_1750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1752 = 8'h8e == _match_key_qbytes_2_T ? phv_data_142 : _GEN_1751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1753 = 8'h8f == _match_key_qbytes_2_T ? phv_data_143 : _GEN_1752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1754 = 8'h90 == _match_key_qbytes_2_T ? phv_data_144 : _GEN_1753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1755 = 8'h91 == _match_key_qbytes_2_T ? phv_data_145 : _GEN_1754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1756 = 8'h92 == _match_key_qbytes_2_T ? phv_data_146 : _GEN_1755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1757 = 8'h93 == _match_key_qbytes_2_T ? phv_data_147 : _GEN_1756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1758 = 8'h94 == _match_key_qbytes_2_T ? phv_data_148 : _GEN_1757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1759 = 8'h95 == _match_key_qbytes_2_T ? phv_data_149 : _GEN_1758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1760 = 8'h96 == _match_key_qbytes_2_T ? phv_data_150 : _GEN_1759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1761 = 8'h97 == _match_key_qbytes_2_T ? phv_data_151 : _GEN_1760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1762 = 8'h98 == _match_key_qbytes_2_T ? phv_data_152 : _GEN_1761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1763 = 8'h99 == _match_key_qbytes_2_T ? phv_data_153 : _GEN_1762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1764 = 8'h9a == _match_key_qbytes_2_T ? phv_data_154 : _GEN_1763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1765 = 8'h9b == _match_key_qbytes_2_T ? phv_data_155 : _GEN_1764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1766 = 8'h9c == _match_key_qbytes_2_T ? phv_data_156 : _GEN_1765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1767 = 8'h9d == _match_key_qbytes_2_T ? phv_data_157 : _GEN_1766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1768 = 8'h9e == _match_key_qbytes_2_T ? phv_data_158 : _GEN_1767; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1769 = 8'h9f == _match_key_qbytes_2_T ? phv_data_159 : _GEN_1768; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1771 = 8'h1 == _match_key_qbytes_2_T_1 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1772 = 8'h2 == _match_key_qbytes_2_T_1 ? phv_data_2 : _GEN_1771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1773 = 8'h3 == _match_key_qbytes_2_T_1 ? phv_data_3 : _GEN_1772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1774 = 8'h4 == _match_key_qbytes_2_T_1 ? phv_data_4 : _GEN_1773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1775 = 8'h5 == _match_key_qbytes_2_T_1 ? phv_data_5 : _GEN_1774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1776 = 8'h6 == _match_key_qbytes_2_T_1 ? phv_data_6 : _GEN_1775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1777 = 8'h7 == _match_key_qbytes_2_T_1 ? phv_data_7 : _GEN_1776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1778 = 8'h8 == _match_key_qbytes_2_T_1 ? phv_data_8 : _GEN_1777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1779 = 8'h9 == _match_key_qbytes_2_T_1 ? phv_data_9 : _GEN_1778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1780 = 8'ha == _match_key_qbytes_2_T_1 ? phv_data_10 : _GEN_1779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1781 = 8'hb == _match_key_qbytes_2_T_1 ? phv_data_11 : _GEN_1780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1782 = 8'hc == _match_key_qbytes_2_T_1 ? phv_data_12 : _GEN_1781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1783 = 8'hd == _match_key_qbytes_2_T_1 ? phv_data_13 : _GEN_1782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1784 = 8'he == _match_key_qbytes_2_T_1 ? phv_data_14 : _GEN_1783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1785 = 8'hf == _match_key_qbytes_2_T_1 ? phv_data_15 : _GEN_1784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1786 = 8'h10 == _match_key_qbytes_2_T_1 ? phv_data_16 : _GEN_1785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1787 = 8'h11 == _match_key_qbytes_2_T_1 ? phv_data_17 : _GEN_1786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1788 = 8'h12 == _match_key_qbytes_2_T_1 ? phv_data_18 : _GEN_1787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1789 = 8'h13 == _match_key_qbytes_2_T_1 ? phv_data_19 : _GEN_1788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1790 = 8'h14 == _match_key_qbytes_2_T_1 ? phv_data_20 : _GEN_1789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1791 = 8'h15 == _match_key_qbytes_2_T_1 ? phv_data_21 : _GEN_1790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1792 = 8'h16 == _match_key_qbytes_2_T_1 ? phv_data_22 : _GEN_1791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1793 = 8'h17 == _match_key_qbytes_2_T_1 ? phv_data_23 : _GEN_1792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1794 = 8'h18 == _match_key_qbytes_2_T_1 ? phv_data_24 : _GEN_1793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1795 = 8'h19 == _match_key_qbytes_2_T_1 ? phv_data_25 : _GEN_1794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1796 = 8'h1a == _match_key_qbytes_2_T_1 ? phv_data_26 : _GEN_1795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1797 = 8'h1b == _match_key_qbytes_2_T_1 ? phv_data_27 : _GEN_1796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1798 = 8'h1c == _match_key_qbytes_2_T_1 ? phv_data_28 : _GEN_1797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1799 = 8'h1d == _match_key_qbytes_2_T_1 ? phv_data_29 : _GEN_1798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1800 = 8'h1e == _match_key_qbytes_2_T_1 ? phv_data_30 : _GEN_1799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1801 = 8'h1f == _match_key_qbytes_2_T_1 ? phv_data_31 : _GEN_1800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1802 = 8'h20 == _match_key_qbytes_2_T_1 ? phv_data_32 : _GEN_1801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1803 = 8'h21 == _match_key_qbytes_2_T_1 ? phv_data_33 : _GEN_1802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1804 = 8'h22 == _match_key_qbytes_2_T_1 ? phv_data_34 : _GEN_1803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1805 = 8'h23 == _match_key_qbytes_2_T_1 ? phv_data_35 : _GEN_1804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1806 = 8'h24 == _match_key_qbytes_2_T_1 ? phv_data_36 : _GEN_1805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1807 = 8'h25 == _match_key_qbytes_2_T_1 ? phv_data_37 : _GEN_1806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1808 = 8'h26 == _match_key_qbytes_2_T_1 ? phv_data_38 : _GEN_1807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1809 = 8'h27 == _match_key_qbytes_2_T_1 ? phv_data_39 : _GEN_1808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1810 = 8'h28 == _match_key_qbytes_2_T_1 ? phv_data_40 : _GEN_1809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1811 = 8'h29 == _match_key_qbytes_2_T_1 ? phv_data_41 : _GEN_1810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1812 = 8'h2a == _match_key_qbytes_2_T_1 ? phv_data_42 : _GEN_1811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1813 = 8'h2b == _match_key_qbytes_2_T_1 ? phv_data_43 : _GEN_1812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1814 = 8'h2c == _match_key_qbytes_2_T_1 ? phv_data_44 : _GEN_1813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1815 = 8'h2d == _match_key_qbytes_2_T_1 ? phv_data_45 : _GEN_1814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1816 = 8'h2e == _match_key_qbytes_2_T_1 ? phv_data_46 : _GEN_1815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1817 = 8'h2f == _match_key_qbytes_2_T_1 ? phv_data_47 : _GEN_1816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1818 = 8'h30 == _match_key_qbytes_2_T_1 ? phv_data_48 : _GEN_1817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1819 = 8'h31 == _match_key_qbytes_2_T_1 ? phv_data_49 : _GEN_1818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1820 = 8'h32 == _match_key_qbytes_2_T_1 ? phv_data_50 : _GEN_1819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1821 = 8'h33 == _match_key_qbytes_2_T_1 ? phv_data_51 : _GEN_1820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1822 = 8'h34 == _match_key_qbytes_2_T_1 ? phv_data_52 : _GEN_1821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1823 = 8'h35 == _match_key_qbytes_2_T_1 ? phv_data_53 : _GEN_1822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1824 = 8'h36 == _match_key_qbytes_2_T_1 ? phv_data_54 : _GEN_1823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1825 = 8'h37 == _match_key_qbytes_2_T_1 ? phv_data_55 : _GEN_1824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1826 = 8'h38 == _match_key_qbytes_2_T_1 ? phv_data_56 : _GEN_1825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1827 = 8'h39 == _match_key_qbytes_2_T_1 ? phv_data_57 : _GEN_1826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1828 = 8'h3a == _match_key_qbytes_2_T_1 ? phv_data_58 : _GEN_1827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1829 = 8'h3b == _match_key_qbytes_2_T_1 ? phv_data_59 : _GEN_1828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1830 = 8'h3c == _match_key_qbytes_2_T_1 ? phv_data_60 : _GEN_1829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1831 = 8'h3d == _match_key_qbytes_2_T_1 ? phv_data_61 : _GEN_1830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1832 = 8'h3e == _match_key_qbytes_2_T_1 ? phv_data_62 : _GEN_1831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1833 = 8'h3f == _match_key_qbytes_2_T_1 ? phv_data_63 : _GEN_1832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1834 = 8'h40 == _match_key_qbytes_2_T_1 ? phv_data_64 : _GEN_1833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1835 = 8'h41 == _match_key_qbytes_2_T_1 ? phv_data_65 : _GEN_1834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1836 = 8'h42 == _match_key_qbytes_2_T_1 ? phv_data_66 : _GEN_1835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1837 = 8'h43 == _match_key_qbytes_2_T_1 ? phv_data_67 : _GEN_1836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1838 = 8'h44 == _match_key_qbytes_2_T_1 ? phv_data_68 : _GEN_1837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1839 = 8'h45 == _match_key_qbytes_2_T_1 ? phv_data_69 : _GEN_1838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1840 = 8'h46 == _match_key_qbytes_2_T_1 ? phv_data_70 : _GEN_1839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1841 = 8'h47 == _match_key_qbytes_2_T_1 ? phv_data_71 : _GEN_1840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1842 = 8'h48 == _match_key_qbytes_2_T_1 ? phv_data_72 : _GEN_1841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1843 = 8'h49 == _match_key_qbytes_2_T_1 ? phv_data_73 : _GEN_1842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1844 = 8'h4a == _match_key_qbytes_2_T_1 ? phv_data_74 : _GEN_1843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1845 = 8'h4b == _match_key_qbytes_2_T_1 ? phv_data_75 : _GEN_1844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1846 = 8'h4c == _match_key_qbytes_2_T_1 ? phv_data_76 : _GEN_1845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1847 = 8'h4d == _match_key_qbytes_2_T_1 ? phv_data_77 : _GEN_1846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1848 = 8'h4e == _match_key_qbytes_2_T_1 ? phv_data_78 : _GEN_1847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1849 = 8'h4f == _match_key_qbytes_2_T_1 ? phv_data_79 : _GEN_1848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1850 = 8'h50 == _match_key_qbytes_2_T_1 ? phv_data_80 : _GEN_1849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1851 = 8'h51 == _match_key_qbytes_2_T_1 ? phv_data_81 : _GEN_1850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1852 = 8'h52 == _match_key_qbytes_2_T_1 ? phv_data_82 : _GEN_1851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1853 = 8'h53 == _match_key_qbytes_2_T_1 ? phv_data_83 : _GEN_1852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1854 = 8'h54 == _match_key_qbytes_2_T_1 ? phv_data_84 : _GEN_1853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1855 = 8'h55 == _match_key_qbytes_2_T_1 ? phv_data_85 : _GEN_1854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1856 = 8'h56 == _match_key_qbytes_2_T_1 ? phv_data_86 : _GEN_1855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1857 = 8'h57 == _match_key_qbytes_2_T_1 ? phv_data_87 : _GEN_1856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1858 = 8'h58 == _match_key_qbytes_2_T_1 ? phv_data_88 : _GEN_1857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1859 = 8'h59 == _match_key_qbytes_2_T_1 ? phv_data_89 : _GEN_1858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1860 = 8'h5a == _match_key_qbytes_2_T_1 ? phv_data_90 : _GEN_1859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1861 = 8'h5b == _match_key_qbytes_2_T_1 ? phv_data_91 : _GEN_1860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1862 = 8'h5c == _match_key_qbytes_2_T_1 ? phv_data_92 : _GEN_1861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1863 = 8'h5d == _match_key_qbytes_2_T_1 ? phv_data_93 : _GEN_1862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1864 = 8'h5e == _match_key_qbytes_2_T_1 ? phv_data_94 : _GEN_1863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1865 = 8'h5f == _match_key_qbytes_2_T_1 ? phv_data_95 : _GEN_1864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1866 = 8'h60 == _match_key_qbytes_2_T_1 ? phv_data_96 : _GEN_1865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1867 = 8'h61 == _match_key_qbytes_2_T_1 ? phv_data_97 : _GEN_1866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1868 = 8'h62 == _match_key_qbytes_2_T_1 ? phv_data_98 : _GEN_1867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1869 = 8'h63 == _match_key_qbytes_2_T_1 ? phv_data_99 : _GEN_1868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1870 = 8'h64 == _match_key_qbytes_2_T_1 ? phv_data_100 : _GEN_1869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1871 = 8'h65 == _match_key_qbytes_2_T_1 ? phv_data_101 : _GEN_1870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1872 = 8'h66 == _match_key_qbytes_2_T_1 ? phv_data_102 : _GEN_1871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1873 = 8'h67 == _match_key_qbytes_2_T_1 ? phv_data_103 : _GEN_1872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1874 = 8'h68 == _match_key_qbytes_2_T_1 ? phv_data_104 : _GEN_1873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1875 = 8'h69 == _match_key_qbytes_2_T_1 ? phv_data_105 : _GEN_1874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1876 = 8'h6a == _match_key_qbytes_2_T_1 ? phv_data_106 : _GEN_1875; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1877 = 8'h6b == _match_key_qbytes_2_T_1 ? phv_data_107 : _GEN_1876; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1878 = 8'h6c == _match_key_qbytes_2_T_1 ? phv_data_108 : _GEN_1877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1879 = 8'h6d == _match_key_qbytes_2_T_1 ? phv_data_109 : _GEN_1878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1880 = 8'h6e == _match_key_qbytes_2_T_1 ? phv_data_110 : _GEN_1879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1881 = 8'h6f == _match_key_qbytes_2_T_1 ? phv_data_111 : _GEN_1880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1882 = 8'h70 == _match_key_qbytes_2_T_1 ? phv_data_112 : _GEN_1881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1883 = 8'h71 == _match_key_qbytes_2_T_1 ? phv_data_113 : _GEN_1882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1884 = 8'h72 == _match_key_qbytes_2_T_1 ? phv_data_114 : _GEN_1883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1885 = 8'h73 == _match_key_qbytes_2_T_1 ? phv_data_115 : _GEN_1884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1886 = 8'h74 == _match_key_qbytes_2_T_1 ? phv_data_116 : _GEN_1885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1887 = 8'h75 == _match_key_qbytes_2_T_1 ? phv_data_117 : _GEN_1886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1888 = 8'h76 == _match_key_qbytes_2_T_1 ? phv_data_118 : _GEN_1887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1889 = 8'h77 == _match_key_qbytes_2_T_1 ? phv_data_119 : _GEN_1888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1890 = 8'h78 == _match_key_qbytes_2_T_1 ? phv_data_120 : _GEN_1889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1891 = 8'h79 == _match_key_qbytes_2_T_1 ? phv_data_121 : _GEN_1890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1892 = 8'h7a == _match_key_qbytes_2_T_1 ? phv_data_122 : _GEN_1891; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1893 = 8'h7b == _match_key_qbytes_2_T_1 ? phv_data_123 : _GEN_1892; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1894 = 8'h7c == _match_key_qbytes_2_T_1 ? phv_data_124 : _GEN_1893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1895 = 8'h7d == _match_key_qbytes_2_T_1 ? phv_data_125 : _GEN_1894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1896 = 8'h7e == _match_key_qbytes_2_T_1 ? phv_data_126 : _GEN_1895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1897 = 8'h7f == _match_key_qbytes_2_T_1 ? phv_data_127 : _GEN_1896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1898 = 8'h80 == _match_key_qbytes_2_T_1 ? phv_data_128 : _GEN_1897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1899 = 8'h81 == _match_key_qbytes_2_T_1 ? phv_data_129 : _GEN_1898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1900 = 8'h82 == _match_key_qbytes_2_T_1 ? phv_data_130 : _GEN_1899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1901 = 8'h83 == _match_key_qbytes_2_T_1 ? phv_data_131 : _GEN_1900; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1902 = 8'h84 == _match_key_qbytes_2_T_1 ? phv_data_132 : _GEN_1901; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1903 = 8'h85 == _match_key_qbytes_2_T_1 ? phv_data_133 : _GEN_1902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1904 = 8'h86 == _match_key_qbytes_2_T_1 ? phv_data_134 : _GEN_1903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1905 = 8'h87 == _match_key_qbytes_2_T_1 ? phv_data_135 : _GEN_1904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1906 = 8'h88 == _match_key_qbytes_2_T_1 ? phv_data_136 : _GEN_1905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1907 = 8'h89 == _match_key_qbytes_2_T_1 ? phv_data_137 : _GEN_1906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1908 = 8'h8a == _match_key_qbytes_2_T_1 ? phv_data_138 : _GEN_1907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1909 = 8'h8b == _match_key_qbytes_2_T_1 ? phv_data_139 : _GEN_1908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1910 = 8'h8c == _match_key_qbytes_2_T_1 ? phv_data_140 : _GEN_1909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1911 = 8'h8d == _match_key_qbytes_2_T_1 ? phv_data_141 : _GEN_1910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1912 = 8'h8e == _match_key_qbytes_2_T_1 ? phv_data_142 : _GEN_1911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1913 = 8'h8f == _match_key_qbytes_2_T_1 ? phv_data_143 : _GEN_1912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1914 = 8'h90 == _match_key_qbytes_2_T_1 ? phv_data_144 : _GEN_1913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1915 = 8'h91 == _match_key_qbytes_2_T_1 ? phv_data_145 : _GEN_1914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1916 = 8'h92 == _match_key_qbytes_2_T_1 ? phv_data_146 : _GEN_1915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1917 = 8'h93 == _match_key_qbytes_2_T_1 ? phv_data_147 : _GEN_1916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1918 = 8'h94 == _match_key_qbytes_2_T_1 ? phv_data_148 : _GEN_1917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1919 = 8'h95 == _match_key_qbytes_2_T_1 ? phv_data_149 : _GEN_1918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1920 = 8'h96 == _match_key_qbytes_2_T_1 ? phv_data_150 : _GEN_1919; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1921 = 8'h97 == _match_key_qbytes_2_T_1 ? phv_data_151 : _GEN_1920; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1922 = 8'h98 == _match_key_qbytes_2_T_1 ? phv_data_152 : _GEN_1921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1923 = 8'h99 == _match_key_qbytes_2_T_1 ? phv_data_153 : _GEN_1922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1924 = 8'h9a == _match_key_qbytes_2_T_1 ? phv_data_154 : _GEN_1923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1925 = 8'h9b == _match_key_qbytes_2_T_1 ? phv_data_155 : _GEN_1924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1926 = 8'h9c == _match_key_qbytes_2_T_1 ? phv_data_156 : _GEN_1925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1927 = 8'h9d == _match_key_qbytes_2_T_1 ? phv_data_157 : _GEN_1926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1928 = 8'h9e == _match_key_qbytes_2_T_1 ? phv_data_158 : _GEN_1927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1929 = 8'h9f == _match_key_qbytes_2_T_1 ? phv_data_159 : _GEN_1928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [31:0] _match_key_qbytes_2_T_3 = {_GEN_1769,_GEN_1929,_GEN_1449,_GEN_1609}; // @[Cat.scala 30:58]
  wire [31:0] match_key_qbytes_2 = local_offset_2 < end_offset ? _match_key_qbytes_2_T_3 : 32'h0; // @[matcher.scala 88:54 matcher.scala 89:45 matcher.scala 97:45]
  wire [7:0] local_offset_3 = 8'hc + read_key_offset; // @[matcher.scala 87:77]
  wire [5:0] match_key_qbytes_3_hi = local_offset_3[7:2]; // @[matcher.scala 91:54]
  wire [7:0] _match_key_qbytes_3_T = {match_key_qbytes_3_hi,2'h3}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_3_T_1 = {match_key_qbytes_3_hi,2'h2}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_3_T_2 = {match_key_qbytes_3_hi,2'h1}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_1932 = 8'h1 == _match_key_qbytes_3_T_2 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1933 = 8'h2 == _match_key_qbytes_3_T_2 ? phv_data_2 : _GEN_1932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1934 = 8'h3 == _match_key_qbytes_3_T_2 ? phv_data_3 : _GEN_1933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1935 = 8'h4 == _match_key_qbytes_3_T_2 ? phv_data_4 : _GEN_1934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1936 = 8'h5 == _match_key_qbytes_3_T_2 ? phv_data_5 : _GEN_1935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1937 = 8'h6 == _match_key_qbytes_3_T_2 ? phv_data_6 : _GEN_1936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1938 = 8'h7 == _match_key_qbytes_3_T_2 ? phv_data_7 : _GEN_1937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1939 = 8'h8 == _match_key_qbytes_3_T_2 ? phv_data_8 : _GEN_1938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1940 = 8'h9 == _match_key_qbytes_3_T_2 ? phv_data_9 : _GEN_1939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1941 = 8'ha == _match_key_qbytes_3_T_2 ? phv_data_10 : _GEN_1940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1942 = 8'hb == _match_key_qbytes_3_T_2 ? phv_data_11 : _GEN_1941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1943 = 8'hc == _match_key_qbytes_3_T_2 ? phv_data_12 : _GEN_1942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1944 = 8'hd == _match_key_qbytes_3_T_2 ? phv_data_13 : _GEN_1943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1945 = 8'he == _match_key_qbytes_3_T_2 ? phv_data_14 : _GEN_1944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1946 = 8'hf == _match_key_qbytes_3_T_2 ? phv_data_15 : _GEN_1945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1947 = 8'h10 == _match_key_qbytes_3_T_2 ? phv_data_16 : _GEN_1946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1948 = 8'h11 == _match_key_qbytes_3_T_2 ? phv_data_17 : _GEN_1947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1949 = 8'h12 == _match_key_qbytes_3_T_2 ? phv_data_18 : _GEN_1948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1950 = 8'h13 == _match_key_qbytes_3_T_2 ? phv_data_19 : _GEN_1949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1951 = 8'h14 == _match_key_qbytes_3_T_2 ? phv_data_20 : _GEN_1950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1952 = 8'h15 == _match_key_qbytes_3_T_2 ? phv_data_21 : _GEN_1951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1953 = 8'h16 == _match_key_qbytes_3_T_2 ? phv_data_22 : _GEN_1952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1954 = 8'h17 == _match_key_qbytes_3_T_2 ? phv_data_23 : _GEN_1953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1955 = 8'h18 == _match_key_qbytes_3_T_2 ? phv_data_24 : _GEN_1954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1956 = 8'h19 == _match_key_qbytes_3_T_2 ? phv_data_25 : _GEN_1955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1957 = 8'h1a == _match_key_qbytes_3_T_2 ? phv_data_26 : _GEN_1956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1958 = 8'h1b == _match_key_qbytes_3_T_2 ? phv_data_27 : _GEN_1957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1959 = 8'h1c == _match_key_qbytes_3_T_2 ? phv_data_28 : _GEN_1958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1960 = 8'h1d == _match_key_qbytes_3_T_2 ? phv_data_29 : _GEN_1959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1961 = 8'h1e == _match_key_qbytes_3_T_2 ? phv_data_30 : _GEN_1960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1962 = 8'h1f == _match_key_qbytes_3_T_2 ? phv_data_31 : _GEN_1961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1963 = 8'h20 == _match_key_qbytes_3_T_2 ? phv_data_32 : _GEN_1962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1964 = 8'h21 == _match_key_qbytes_3_T_2 ? phv_data_33 : _GEN_1963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1965 = 8'h22 == _match_key_qbytes_3_T_2 ? phv_data_34 : _GEN_1964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1966 = 8'h23 == _match_key_qbytes_3_T_2 ? phv_data_35 : _GEN_1965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1967 = 8'h24 == _match_key_qbytes_3_T_2 ? phv_data_36 : _GEN_1966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1968 = 8'h25 == _match_key_qbytes_3_T_2 ? phv_data_37 : _GEN_1967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1969 = 8'h26 == _match_key_qbytes_3_T_2 ? phv_data_38 : _GEN_1968; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1970 = 8'h27 == _match_key_qbytes_3_T_2 ? phv_data_39 : _GEN_1969; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1971 = 8'h28 == _match_key_qbytes_3_T_2 ? phv_data_40 : _GEN_1970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1972 = 8'h29 == _match_key_qbytes_3_T_2 ? phv_data_41 : _GEN_1971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1973 = 8'h2a == _match_key_qbytes_3_T_2 ? phv_data_42 : _GEN_1972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1974 = 8'h2b == _match_key_qbytes_3_T_2 ? phv_data_43 : _GEN_1973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1975 = 8'h2c == _match_key_qbytes_3_T_2 ? phv_data_44 : _GEN_1974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1976 = 8'h2d == _match_key_qbytes_3_T_2 ? phv_data_45 : _GEN_1975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1977 = 8'h2e == _match_key_qbytes_3_T_2 ? phv_data_46 : _GEN_1976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1978 = 8'h2f == _match_key_qbytes_3_T_2 ? phv_data_47 : _GEN_1977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1979 = 8'h30 == _match_key_qbytes_3_T_2 ? phv_data_48 : _GEN_1978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1980 = 8'h31 == _match_key_qbytes_3_T_2 ? phv_data_49 : _GEN_1979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1981 = 8'h32 == _match_key_qbytes_3_T_2 ? phv_data_50 : _GEN_1980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1982 = 8'h33 == _match_key_qbytes_3_T_2 ? phv_data_51 : _GEN_1981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1983 = 8'h34 == _match_key_qbytes_3_T_2 ? phv_data_52 : _GEN_1982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1984 = 8'h35 == _match_key_qbytes_3_T_2 ? phv_data_53 : _GEN_1983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1985 = 8'h36 == _match_key_qbytes_3_T_2 ? phv_data_54 : _GEN_1984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1986 = 8'h37 == _match_key_qbytes_3_T_2 ? phv_data_55 : _GEN_1985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1987 = 8'h38 == _match_key_qbytes_3_T_2 ? phv_data_56 : _GEN_1986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1988 = 8'h39 == _match_key_qbytes_3_T_2 ? phv_data_57 : _GEN_1987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1989 = 8'h3a == _match_key_qbytes_3_T_2 ? phv_data_58 : _GEN_1988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1990 = 8'h3b == _match_key_qbytes_3_T_2 ? phv_data_59 : _GEN_1989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1991 = 8'h3c == _match_key_qbytes_3_T_2 ? phv_data_60 : _GEN_1990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1992 = 8'h3d == _match_key_qbytes_3_T_2 ? phv_data_61 : _GEN_1991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1993 = 8'h3e == _match_key_qbytes_3_T_2 ? phv_data_62 : _GEN_1992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1994 = 8'h3f == _match_key_qbytes_3_T_2 ? phv_data_63 : _GEN_1993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1995 = 8'h40 == _match_key_qbytes_3_T_2 ? phv_data_64 : _GEN_1994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1996 = 8'h41 == _match_key_qbytes_3_T_2 ? phv_data_65 : _GEN_1995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1997 = 8'h42 == _match_key_qbytes_3_T_2 ? phv_data_66 : _GEN_1996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1998 = 8'h43 == _match_key_qbytes_3_T_2 ? phv_data_67 : _GEN_1997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1999 = 8'h44 == _match_key_qbytes_3_T_2 ? phv_data_68 : _GEN_1998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2000 = 8'h45 == _match_key_qbytes_3_T_2 ? phv_data_69 : _GEN_1999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2001 = 8'h46 == _match_key_qbytes_3_T_2 ? phv_data_70 : _GEN_2000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2002 = 8'h47 == _match_key_qbytes_3_T_2 ? phv_data_71 : _GEN_2001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2003 = 8'h48 == _match_key_qbytes_3_T_2 ? phv_data_72 : _GEN_2002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2004 = 8'h49 == _match_key_qbytes_3_T_2 ? phv_data_73 : _GEN_2003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2005 = 8'h4a == _match_key_qbytes_3_T_2 ? phv_data_74 : _GEN_2004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2006 = 8'h4b == _match_key_qbytes_3_T_2 ? phv_data_75 : _GEN_2005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2007 = 8'h4c == _match_key_qbytes_3_T_2 ? phv_data_76 : _GEN_2006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2008 = 8'h4d == _match_key_qbytes_3_T_2 ? phv_data_77 : _GEN_2007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2009 = 8'h4e == _match_key_qbytes_3_T_2 ? phv_data_78 : _GEN_2008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2010 = 8'h4f == _match_key_qbytes_3_T_2 ? phv_data_79 : _GEN_2009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2011 = 8'h50 == _match_key_qbytes_3_T_2 ? phv_data_80 : _GEN_2010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2012 = 8'h51 == _match_key_qbytes_3_T_2 ? phv_data_81 : _GEN_2011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2013 = 8'h52 == _match_key_qbytes_3_T_2 ? phv_data_82 : _GEN_2012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2014 = 8'h53 == _match_key_qbytes_3_T_2 ? phv_data_83 : _GEN_2013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2015 = 8'h54 == _match_key_qbytes_3_T_2 ? phv_data_84 : _GEN_2014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2016 = 8'h55 == _match_key_qbytes_3_T_2 ? phv_data_85 : _GEN_2015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2017 = 8'h56 == _match_key_qbytes_3_T_2 ? phv_data_86 : _GEN_2016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2018 = 8'h57 == _match_key_qbytes_3_T_2 ? phv_data_87 : _GEN_2017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2019 = 8'h58 == _match_key_qbytes_3_T_2 ? phv_data_88 : _GEN_2018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2020 = 8'h59 == _match_key_qbytes_3_T_2 ? phv_data_89 : _GEN_2019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2021 = 8'h5a == _match_key_qbytes_3_T_2 ? phv_data_90 : _GEN_2020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2022 = 8'h5b == _match_key_qbytes_3_T_2 ? phv_data_91 : _GEN_2021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2023 = 8'h5c == _match_key_qbytes_3_T_2 ? phv_data_92 : _GEN_2022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2024 = 8'h5d == _match_key_qbytes_3_T_2 ? phv_data_93 : _GEN_2023; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2025 = 8'h5e == _match_key_qbytes_3_T_2 ? phv_data_94 : _GEN_2024; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2026 = 8'h5f == _match_key_qbytes_3_T_2 ? phv_data_95 : _GEN_2025; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2027 = 8'h60 == _match_key_qbytes_3_T_2 ? phv_data_96 : _GEN_2026; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2028 = 8'h61 == _match_key_qbytes_3_T_2 ? phv_data_97 : _GEN_2027; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2029 = 8'h62 == _match_key_qbytes_3_T_2 ? phv_data_98 : _GEN_2028; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2030 = 8'h63 == _match_key_qbytes_3_T_2 ? phv_data_99 : _GEN_2029; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2031 = 8'h64 == _match_key_qbytes_3_T_2 ? phv_data_100 : _GEN_2030; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2032 = 8'h65 == _match_key_qbytes_3_T_2 ? phv_data_101 : _GEN_2031; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2033 = 8'h66 == _match_key_qbytes_3_T_2 ? phv_data_102 : _GEN_2032; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2034 = 8'h67 == _match_key_qbytes_3_T_2 ? phv_data_103 : _GEN_2033; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2035 = 8'h68 == _match_key_qbytes_3_T_2 ? phv_data_104 : _GEN_2034; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2036 = 8'h69 == _match_key_qbytes_3_T_2 ? phv_data_105 : _GEN_2035; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2037 = 8'h6a == _match_key_qbytes_3_T_2 ? phv_data_106 : _GEN_2036; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2038 = 8'h6b == _match_key_qbytes_3_T_2 ? phv_data_107 : _GEN_2037; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2039 = 8'h6c == _match_key_qbytes_3_T_2 ? phv_data_108 : _GEN_2038; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2040 = 8'h6d == _match_key_qbytes_3_T_2 ? phv_data_109 : _GEN_2039; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2041 = 8'h6e == _match_key_qbytes_3_T_2 ? phv_data_110 : _GEN_2040; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2042 = 8'h6f == _match_key_qbytes_3_T_2 ? phv_data_111 : _GEN_2041; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2043 = 8'h70 == _match_key_qbytes_3_T_2 ? phv_data_112 : _GEN_2042; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2044 = 8'h71 == _match_key_qbytes_3_T_2 ? phv_data_113 : _GEN_2043; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2045 = 8'h72 == _match_key_qbytes_3_T_2 ? phv_data_114 : _GEN_2044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2046 = 8'h73 == _match_key_qbytes_3_T_2 ? phv_data_115 : _GEN_2045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2047 = 8'h74 == _match_key_qbytes_3_T_2 ? phv_data_116 : _GEN_2046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2048 = 8'h75 == _match_key_qbytes_3_T_2 ? phv_data_117 : _GEN_2047; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2049 = 8'h76 == _match_key_qbytes_3_T_2 ? phv_data_118 : _GEN_2048; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2050 = 8'h77 == _match_key_qbytes_3_T_2 ? phv_data_119 : _GEN_2049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2051 = 8'h78 == _match_key_qbytes_3_T_2 ? phv_data_120 : _GEN_2050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2052 = 8'h79 == _match_key_qbytes_3_T_2 ? phv_data_121 : _GEN_2051; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2053 = 8'h7a == _match_key_qbytes_3_T_2 ? phv_data_122 : _GEN_2052; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2054 = 8'h7b == _match_key_qbytes_3_T_2 ? phv_data_123 : _GEN_2053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2055 = 8'h7c == _match_key_qbytes_3_T_2 ? phv_data_124 : _GEN_2054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2056 = 8'h7d == _match_key_qbytes_3_T_2 ? phv_data_125 : _GEN_2055; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2057 = 8'h7e == _match_key_qbytes_3_T_2 ? phv_data_126 : _GEN_2056; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2058 = 8'h7f == _match_key_qbytes_3_T_2 ? phv_data_127 : _GEN_2057; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2059 = 8'h80 == _match_key_qbytes_3_T_2 ? phv_data_128 : _GEN_2058; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2060 = 8'h81 == _match_key_qbytes_3_T_2 ? phv_data_129 : _GEN_2059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2061 = 8'h82 == _match_key_qbytes_3_T_2 ? phv_data_130 : _GEN_2060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2062 = 8'h83 == _match_key_qbytes_3_T_2 ? phv_data_131 : _GEN_2061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2063 = 8'h84 == _match_key_qbytes_3_T_2 ? phv_data_132 : _GEN_2062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2064 = 8'h85 == _match_key_qbytes_3_T_2 ? phv_data_133 : _GEN_2063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2065 = 8'h86 == _match_key_qbytes_3_T_2 ? phv_data_134 : _GEN_2064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2066 = 8'h87 == _match_key_qbytes_3_T_2 ? phv_data_135 : _GEN_2065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2067 = 8'h88 == _match_key_qbytes_3_T_2 ? phv_data_136 : _GEN_2066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2068 = 8'h89 == _match_key_qbytes_3_T_2 ? phv_data_137 : _GEN_2067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2069 = 8'h8a == _match_key_qbytes_3_T_2 ? phv_data_138 : _GEN_2068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2070 = 8'h8b == _match_key_qbytes_3_T_2 ? phv_data_139 : _GEN_2069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2071 = 8'h8c == _match_key_qbytes_3_T_2 ? phv_data_140 : _GEN_2070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2072 = 8'h8d == _match_key_qbytes_3_T_2 ? phv_data_141 : _GEN_2071; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2073 = 8'h8e == _match_key_qbytes_3_T_2 ? phv_data_142 : _GEN_2072; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2074 = 8'h8f == _match_key_qbytes_3_T_2 ? phv_data_143 : _GEN_2073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2075 = 8'h90 == _match_key_qbytes_3_T_2 ? phv_data_144 : _GEN_2074; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2076 = 8'h91 == _match_key_qbytes_3_T_2 ? phv_data_145 : _GEN_2075; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2077 = 8'h92 == _match_key_qbytes_3_T_2 ? phv_data_146 : _GEN_2076; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2078 = 8'h93 == _match_key_qbytes_3_T_2 ? phv_data_147 : _GEN_2077; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2079 = 8'h94 == _match_key_qbytes_3_T_2 ? phv_data_148 : _GEN_2078; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2080 = 8'h95 == _match_key_qbytes_3_T_2 ? phv_data_149 : _GEN_2079; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2081 = 8'h96 == _match_key_qbytes_3_T_2 ? phv_data_150 : _GEN_2080; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2082 = 8'h97 == _match_key_qbytes_3_T_2 ? phv_data_151 : _GEN_2081; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2083 = 8'h98 == _match_key_qbytes_3_T_2 ? phv_data_152 : _GEN_2082; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2084 = 8'h99 == _match_key_qbytes_3_T_2 ? phv_data_153 : _GEN_2083; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2085 = 8'h9a == _match_key_qbytes_3_T_2 ? phv_data_154 : _GEN_2084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2086 = 8'h9b == _match_key_qbytes_3_T_2 ? phv_data_155 : _GEN_2085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2087 = 8'h9c == _match_key_qbytes_3_T_2 ? phv_data_156 : _GEN_2086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2088 = 8'h9d == _match_key_qbytes_3_T_2 ? phv_data_157 : _GEN_2087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2089 = 8'h9e == _match_key_qbytes_3_T_2 ? phv_data_158 : _GEN_2088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2090 = 8'h9f == _match_key_qbytes_3_T_2 ? phv_data_159 : _GEN_2089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2092 = 8'h1 == local_offset_3 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2093 = 8'h2 == local_offset_3 ? phv_data_2 : _GEN_2092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2094 = 8'h3 == local_offset_3 ? phv_data_3 : _GEN_2093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2095 = 8'h4 == local_offset_3 ? phv_data_4 : _GEN_2094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2096 = 8'h5 == local_offset_3 ? phv_data_5 : _GEN_2095; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2097 = 8'h6 == local_offset_3 ? phv_data_6 : _GEN_2096; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2098 = 8'h7 == local_offset_3 ? phv_data_7 : _GEN_2097; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2099 = 8'h8 == local_offset_3 ? phv_data_8 : _GEN_2098; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2100 = 8'h9 == local_offset_3 ? phv_data_9 : _GEN_2099; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2101 = 8'ha == local_offset_3 ? phv_data_10 : _GEN_2100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2102 = 8'hb == local_offset_3 ? phv_data_11 : _GEN_2101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2103 = 8'hc == local_offset_3 ? phv_data_12 : _GEN_2102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2104 = 8'hd == local_offset_3 ? phv_data_13 : _GEN_2103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2105 = 8'he == local_offset_3 ? phv_data_14 : _GEN_2104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2106 = 8'hf == local_offset_3 ? phv_data_15 : _GEN_2105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2107 = 8'h10 == local_offset_3 ? phv_data_16 : _GEN_2106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2108 = 8'h11 == local_offset_3 ? phv_data_17 : _GEN_2107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2109 = 8'h12 == local_offset_3 ? phv_data_18 : _GEN_2108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2110 = 8'h13 == local_offset_3 ? phv_data_19 : _GEN_2109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2111 = 8'h14 == local_offset_3 ? phv_data_20 : _GEN_2110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2112 = 8'h15 == local_offset_3 ? phv_data_21 : _GEN_2111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2113 = 8'h16 == local_offset_3 ? phv_data_22 : _GEN_2112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2114 = 8'h17 == local_offset_3 ? phv_data_23 : _GEN_2113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2115 = 8'h18 == local_offset_3 ? phv_data_24 : _GEN_2114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2116 = 8'h19 == local_offset_3 ? phv_data_25 : _GEN_2115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2117 = 8'h1a == local_offset_3 ? phv_data_26 : _GEN_2116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2118 = 8'h1b == local_offset_3 ? phv_data_27 : _GEN_2117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2119 = 8'h1c == local_offset_3 ? phv_data_28 : _GEN_2118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2120 = 8'h1d == local_offset_3 ? phv_data_29 : _GEN_2119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2121 = 8'h1e == local_offset_3 ? phv_data_30 : _GEN_2120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2122 = 8'h1f == local_offset_3 ? phv_data_31 : _GEN_2121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2123 = 8'h20 == local_offset_3 ? phv_data_32 : _GEN_2122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2124 = 8'h21 == local_offset_3 ? phv_data_33 : _GEN_2123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2125 = 8'h22 == local_offset_3 ? phv_data_34 : _GEN_2124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2126 = 8'h23 == local_offset_3 ? phv_data_35 : _GEN_2125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2127 = 8'h24 == local_offset_3 ? phv_data_36 : _GEN_2126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2128 = 8'h25 == local_offset_3 ? phv_data_37 : _GEN_2127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2129 = 8'h26 == local_offset_3 ? phv_data_38 : _GEN_2128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2130 = 8'h27 == local_offset_3 ? phv_data_39 : _GEN_2129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2131 = 8'h28 == local_offset_3 ? phv_data_40 : _GEN_2130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2132 = 8'h29 == local_offset_3 ? phv_data_41 : _GEN_2131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2133 = 8'h2a == local_offset_3 ? phv_data_42 : _GEN_2132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2134 = 8'h2b == local_offset_3 ? phv_data_43 : _GEN_2133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2135 = 8'h2c == local_offset_3 ? phv_data_44 : _GEN_2134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2136 = 8'h2d == local_offset_3 ? phv_data_45 : _GEN_2135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2137 = 8'h2e == local_offset_3 ? phv_data_46 : _GEN_2136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2138 = 8'h2f == local_offset_3 ? phv_data_47 : _GEN_2137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2139 = 8'h30 == local_offset_3 ? phv_data_48 : _GEN_2138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2140 = 8'h31 == local_offset_3 ? phv_data_49 : _GEN_2139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2141 = 8'h32 == local_offset_3 ? phv_data_50 : _GEN_2140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2142 = 8'h33 == local_offset_3 ? phv_data_51 : _GEN_2141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2143 = 8'h34 == local_offset_3 ? phv_data_52 : _GEN_2142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2144 = 8'h35 == local_offset_3 ? phv_data_53 : _GEN_2143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2145 = 8'h36 == local_offset_3 ? phv_data_54 : _GEN_2144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2146 = 8'h37 == local_offset_3 ? phv_data_55 : _GEN_2145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2147 = 8'h38 == local_offset_3 ? phv_data_56 : _GEN_2146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2148 = 8'h39 == local_offset_3 ? phv_data_57 : _GEN_2147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2149 = 8'h3a == local_offset_3 ? phv_data_58 : _GEN_2148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2150 = 8'h3b == local_offset_3 ? phv_data_59 : _GEN_2149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2151 = 8'h3c == local_offset_3 ? phv_data_60 : _GEN_2150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2152 = 8'h3d == local_offset_3 ? phv_data_61 : _GEN_2151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2153 = 8'h3e == local_offset_3 ? phv_data_62 : _GEN_2152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2154 = 8'h3f == local_offset_3 ? phv_data_63 : _GEN_2153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2155 = 8'h40 == local_offset_3 ? phv_data_64 : _GEN_2154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2156 = 8'h41 == local_offset_3 ? phv_data_65 : _GEN_2155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2157 = 8'h42 == local_offset_3 ? phv_data_66 : _GEN_2156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2158 = 8'h43 == local_offset_3 ? phv_data_67 : _GEN_2157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2159 = 8'h44 == local_offset_3 ? phv_data_68 : _GEN_2158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2160 = 8'h45 == local_offset_3 ? phv_data_69 : _GEN_2159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2161 = 8'h46 == local_offset_3 ? phv_data_70 : _GEN_2160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2162 = 8'h47 == local_offset_3 ? phv_data_71 : _GEN_2161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2163 = 8'h48 == local_offset_3 ? phv_data_72 : _GEN_2162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2164 = 8'h49 == local_offset_3 ? phv_data_73 : _GEN_2163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2165 = 8'h4a == local_offset_3 ? phv_data_74 : _GEN_2164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2166 = 8'h4b == local_offset_3 ? phv_data_75 : _GEN_2165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2167 = 8'h4c == local_offset_3 ? phv_data_76 : _GEN_2166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2168 = 8'h4d == local_offset_3 ? phv_data_77 : _GEN_2167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2169 = 8'h4e == local_offset_3 ? phv_data_78 : _GEN_2168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2170 = 8'h4f == local_offset_3 ? phv_data_79 : _GEN_2169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2171 = 8'h50 == local_offset_3 ? phv_data_80 : _GEN_2170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2172 = 8'h51 == local_offset_3 ? phv_data_81 : _GEN_2171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2173 = 8'h52 == local_offset_3 ? phv_data_82 : _GEN_2172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2174 = 8'h53 == local_offset_3 ? phv_data_83 : _GEN_2173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2175 = 8'h54 == local_offset_3 ? phv_data_84 : _GEN_2174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2176 = 8'h55 == local_offset_3 ? phv_data_85 : _GEN_2175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2177 = 8'h56 == local_offset_3 ? phv_data_86 : _GEN_2176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2178 = 8'h57 == local_offset_3 ? phv_data_87 : _GEN_2177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2179 = 8'h58 == local_offset_3 ? phv_data_88 : _GEN_2178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2180 = 8'h59 == local_offset_3 ? phv_data_89 : _GEN_2179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2181 = 8'h5a == local_offset_3 ? phv_data_90 : _GEN_2180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2182 = 8'h5b == local_offset_3 ? phv_data_91 : _GEN_2181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2183 = 8'h5c == local_offset_3 ? phv_data_92 : _GEN_2182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2184 = 8'h5d == local_offset_3 ? phv_data_93 : _GEN_2183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2185 = 8'h5e == local_offset_3 ? phv_data_94 : _GEN_2184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2186 = 8'h5f == local_offset_3 ? phv_data_95 : _GEN_2185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2187 = 8'h60 == local_offset_3 ? phv_data_96 : _GEN_2186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2188 = 8'h61 == local_offset_3 ? phv_data_97 : _GEN_2187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2189 = 8'h62 == local_offset_3 ? phv_data_98 : _GEN_2188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2190 = 8'h63 == local_offset_3 ? phv_data_99 : _GEN_2189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2191 = 8'h64 == local_offset_3 ? phv_data_100 : _GEN_2190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2192 = 8'h65 == local_offset_3 ? phv_data_101 : _GEN_2191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2193 = 8'h66 == local_offset_3 ? phv_data_102 : _GEN_2192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2194 = 8'h67 == local_offset_3 ? phv_data_103 : _GEN_2193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2195 = 8'h68 == local_offset_3 ? phv_data_104 : _GEN_2194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2196 = 8'h69 == local_offset_3 ? phv_data_105 : _GEN_2195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2197 = 8'h6a == local_offset_3 ? phv_data_106 : _GEN_2196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2198 = 8'h6b == local_offset_3 ? phv_data_107 : _GEN_2197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2199 = 8'h6c == local_offset_3 ? phv_data_108 : _GEN_2198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2200 = 8'h6d == local_offset_3 ? phv_data_109 : _GEN_2199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2201 = 8'h6e == local_offset_3 ? phv_data_110 : _GEN_2200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2202 = 8'h6f == local_offset_3 ? phv_data_111 : _GEN_2201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2203 = 8'h70 == local_offset_3 ? phv_data_112 : _GEN_2202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2204 = 8'h71 == local_offset_3 ? phv_data_113 : _GEN_2203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2205 = 8'h72 == local_offset_3 ? phv_data_114 : _GEN_2204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2206 = 8'h73 == local_offset_3 ? phv_data_115 : _GEN_2205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2207 = 8'h74 == local_offset_3 ? phv_data_116 : _GEN_2206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2208 = 8'h75 == local_offset_3 ? phv_data_117 : _GEN_2207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2209 = 8'h76 == local_offset_3 ? phv_data_118 : _GEN_2208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2210 = 8'h77 == local_offset_3 ? phv_data_119 : _GEN_2209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2211 = 8'h78 == local_offset_3 ? phv_data_120 : _GEN_2210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2212 = 8'h79 == local_offset_3 ? phv_data_121 : _GEN_2211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2213 = 8'h7a == local_offset_3 ? phv_data_122 : _GEN_2212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2214 = 8'h7b == local_offset_3 ? phv_data_123 : _GEN_2213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2215 = 8'h7c == local_offset_3 ? phv_data_124 : _GEN_2214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2216 = 8'h7d == local_offset_3 ? phv_data_125 : _GEN_2215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2217 = 8'h7e == local_offset_3 ? phv_data_126 : _GEN_2216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2218 = 8'h7f == local_offset_3 ? phv_data_127 : _GEN_2217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2219 = 8'h80 == local_offset_3 ? phv_data_128 : _GEN_2218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2220 = 8'h81 == local_offset_3 ? phv_data_129 : _GEN_2219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2221 = 8'h82 == local_offset_3 ? phv_data_130 : _GEN_2220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2222 = 8'h83 == local_offset_3 ? phv_data_131 : _GEN_2221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2223 = 8'h84 == local_offset_3 ? phv_data_132 : _GEN_2222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2224 = 8'h85 == local_offset_3 ? phv_data_133 : _GEN_2223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2225 = 8'h86 == local_offset_3 ? phv_data_134 : _GEN_2224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2226 = 8'h87 == local_offset_3 ? phv_data_135 : _GEN_2225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2227 = 8'h88 == local_offset_3 ? phv_data_136 : _GEN_2226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2228 = 8'h89 == local_offset_3 ? phv_data_137 : _GEN_2227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2229 = 8'h8a == local_offset_3 ? phv_data_138 : _GEN_2228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2230 = 8'h8b == local_offset_3 ? phv_data_139 : _GEN_2229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2231 = 8'h8c == local_offset_3 ? phv_data_140 : _GEN_2230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2232 = 8'h8d == local_offset_3 ? phv_data_141 : _GEN_2231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2233 = 8'h8e == local_offset_3 ? phv_data_142 : _GEN_2232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2234 = 8'h8f == local_offset_3 ? phv_data_143 : _GEN_2233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2235 = 8'h90 == local_offset_3 ? phv_data_144 : _GEN_2234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2236 = 8'h91 == local_offset_3 ? phv_data_145 : _GEN_2235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2237 = 8'h92 == local_offset_3 ? phv_data_146 : _GEN_2236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2238 = 8'h93 == local_offset_3 ? phv_data_147 : _GEN_2237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2239 = 8'h94 == local_offset_3 ? phv_data_148 : _GEN_2238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2240 = 8'h95 == local_offset_3 ? phv_data_149 : _GEN_2239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2241 = 8'h96 == local_offset_3 ? phv_data_150 : _GEN_2240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2242 = 8'h97 == local_offset_3 ? phv_data_151 : _GEN_2241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2243 = 8'h98 == local_offset_3 ? phv_data_152 : _GEN_2242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2244 = 8'h99 == local_offset_3 ? phv_data_153 : _GEN_2243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2245 = 8'h9a == local_offset_3 ? phv_data_154 : _GEN_2244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2246 = 8'h9b == local_offset_3 ? phv_data_155 : _GEN_2245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2247 = 8'h9c == local_offset_3 ? phv_data_156 : _GEN_2246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2248 = 8'h9d == local_offset_3 ? phv_data_157 : _GEN_2247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2249 = 8'h9e == local_offset_3 ? phv_data_158 : _GEN_2248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2250 = 8'h9f == local_offset_3 ? phv_data_159 : _GEN_2249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2252 = 8'h1 == _match_key_qbytes_3_T ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2253 = 8'h2 == _match_key_qbytes_3_T ? phv_data_2 : _GEN_2252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2254 = 8'h3 == _match_key_qbytes_3_T ? phv_data_3 : _GEN_2253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2255 = 8'h4 == _match_key_qbytes_3_T ? phv_data_4 : _GEN_2254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2256 = 8'h5 == _match_key_qbytes_3_T ? phv_data_5 : _GEN_2255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2257 = 8'h6 == _match_key_qbytes_3_T ? phv_data_6 : _GEN_2256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2258 = 8'h7 == _match_key_qbytes_3_T ? phv_data_7 : _GEN_2257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2259 = 8'h8 == _match_key_qbytes_3_T ? phv_data_8 : _GEN_2258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2260 = 8'h9 == _match_key_qbytes_3_T ? phv_data_9 : _GEN_2259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2261 = 8'ha == _match_key_qbytes_3_T ? phv_data_10 : _GEN_2260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2262 = 8'hb == _match_key_qbytes_3_T ? phv_data_11 : _GEN_2261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2263 = 8'hc == _match_key_qbytes_3_T ? phv_data_12 : _GEN_2262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2264 = 8'hd == _match_key_qbytes_3_T ? phv_data_13 : _GEN_2263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2265 = 8'he == _match_key_qbytes_3_T ? phv_data_14 : _GEN_2264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2266 = 8'hf == _match_key_qbytes_3_T ? phv_data_15 : _GEN_2265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2267 = 8'h10 == _match_key_qbytes_3_T ? phv_data_16 : _GEN_2266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2268 = 8'h11 == _match_key_qbytes_3_T ? phv_data_17 : _GEN_2267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2269 = 8'h12 == _match_key_qbytes_3_T ? phv_data_18 : _GEN_2268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2270 = 8'h13 == _match_key_qbytes_3_T ? phv_data_19 : _GEN_2269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2271 = 8'h14 == _match_key_qbytes_3_T ? phv_data_20 : _GEN_2270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2272 = 8'h15 == _match_key_qbytes_3_T ? phv_data_21 : _GEN_2271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2273 = 8'h16 == _match_key_qbytes_3_T ? phv_data_22 : _GEN_2272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2274 = 8'h17 == _match_key_qbytes_3_T ? phv_data_23 : _GEN_2273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2275 = 8'h18 == _match_key_qbytes_3_T ? phv_data_24 : _GEN_2274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2276 = 8'h19 == _match_key_qbytes_3_T ? phv_data_25 : _GEN_2275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2277 = 8'h1a == _match_key_qbytes_3_T ? phv_data_26 : _GEN_2276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2278 = 8'h1b == _match_key_qbytes_3_T ? phv_data_27 : _GEN_2277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2279 = 8'h1c == _match_key_qbytes_3_T ? phv_data_28 : _GEN_2278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2280 = 8'h1d == _match_key_qbytes_3_T ? phv_data_29 : _GEN_2279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2281 = 8'h1e == _match_key_qbytes_3_T ? phv_data_30 : _GEN_2280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2282 = 8'h1f == _match_key_qbytes_3_T ? phv_data_31 : _GEN_2281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2283 = 8'h20 == _match_key_qbytes_3_T ? phv_data_32 : _GEN_2282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2284 = 8'h21 == _match_key_qbytes_3_T ? phv_data_33 : _GEN_2283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2285 = 8'h22 == _match_key_qbytes_3_T ? phv_data_34 : _GEN_2284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2286 = 8'h23 == _match_key_qbytes_3_T ? phv_data_35 : _GEN_2285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2287 = 8'h24 == _match_key_qbytes_3_T ? phv_data_36 : _GEN_2286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2288 = 8'h25 == _match_key_qbytes_3_T ? phv_data_37 : _GEN_2287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2289 = 8'h26 == _match_key_qbytes_3_T ? phv_data_38 : _GEN_2288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2290 = 8'h27 == _match_key_qbytes_3_T ? phv_data_39 : _GEN_2289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2291 = 8'h28 == _match_key_qbytes_3_T ? phv_data_40 : _GEN_2290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2292 = 8'h29 == _match_key_qbytes_3_T ? phv_data_41 : _GEN_2291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2293 = 8'h2a == _match_key_qbytes_3_T ? phv_data_42 : _GEN_2292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2294 = 8'h2b == _match_key_qbytes_3_T ? phv_data_43 : _GEN_2293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2295 = 8'h2c == _match_key_qbytes_3_T ? phv_data_44 : _GEN_2294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2296 = 8'h2d == _match_key_qbytes_3_T ? phv_data_45 : _GEN_2295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2297 = 8'h2e == _match_key_qbytes_3_T ? phv_data_46 : _GEN_2296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2298 = 8'h2f == _match_key_qbytes_3_T ? phv_data_47 : _GEN_2297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2299 = 8'h30 == _match_key_qbytes_3_T ? phv_data_48 : _GEN_2298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2300 = 8'h31 == _match_key_qbytes_3_T ? phv_data_49 : _GEN_2299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2301 = 8'h32 == _match_key_qbytes_3_T ? phv_data_50 : _GEN_2300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2302 = 8'h33 == _match_key_qbytes_3_T ? phv_data_51 : _GEN_2301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2303 = 8'h34 == _match_key_qbytes_3_T ? phv_data_52 : _GEN_2302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2304 = 8'h35 == _match_key_qbytes_3_T ? phv_data_53 : _GEN_2303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2305 = 8'h36 == _match_key_qbytes_3_T ? phv_data_54 : _GEN_2304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2306 = 8'h37 == _match_key_qbytes_3_T ? phv_data_55 : _GEN_2305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2307 = 8'h38 == _match_key_qbytes_3_T ? phv_data_56 : _GEN_2306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2308 = 8'h39 == _match_key_qbytes_3_T ? phv_data_57 : _GEN_2307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2309 = 8'h3a == _match_key_qbytes_3_T ? phv_data_58 : _GEN_2308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2310 = 8'h3b == _match_key_qbytes_3_T ? phv_data_59 : _GEN_2309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2311 = 8'h3c == _match_key_qbytes_3_T ? phv_data_60 : _GEN_2310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2312 = 8'h3d == _match_key_qbytes_3_T ? phv_data_61 : _GEN_2311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2313 = 8'h3e == _match_key_qbytes_3_T ? phv_data_62 : _GEN_2312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2314 = 8'h3f == _match_key_qbytes_3_T ? phv_data_63 : _GEN_2313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2315 = 8'h40 == _match_key_qbytes_3_T ? phv_data_64 : _GEN_2314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2316 = 8'h41 == _match_key_qbytes_3_T ? phv_data_65 : _GEN_2315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2317 = 8'h42 == _match_key_qbytes_3_T ? phv_data_66 : _GEN_2316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2318 = 8'h43 == _match_key_qbytes_3_T ? phv_data_67 : _GEN_2317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2319 = 8'h44 == _match_key_qbytes_3_T ? phv_data_68 : _GEN_2318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2320 = 8'h45 == _match_key_qbytes_3_T ? phv_data_69 : _GEN_2319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2321 = 8'h46 == _match_key_qbytes_3_T ? phv_data_70 : _GEN_2320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2322 = 8'h47 == _match_key_qbytes_3_T ? phv_data_71 : _GEN_2321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2323 = 8'h48 == _match_key_qbytes_3_T ? phv_data_72 : _GEN_2322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2324 = 8'h49 == _match_key_qbytes_3_T ? phv_data_73 : _GEN_2323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2325 = 8'h4a == _match_key_qbytes_3_T ? phv_data_74 : _GEN_2324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2326 = 8'h4b == _match_key_qbytes_3_T ? phv_data_75 : _GEN_2325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2327 = 8'h4c == _match_key_qbytes_3_T ? phv_data_76 : _GEN_2326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2328 = 8'h4d == _match_key_qbytes_3_T ? phv_data_77 : _GEN_2327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2329 = 8'h4e == _match_key_qbytes_3_T ? phv_data_78 : _GEN_2328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2330 = 8'h4f == _match_key_qbytes_3_T ? phv_data_79 : _GEN_2329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2331 = 8'h50 == _match_key_qbytes_3_T ? phv_data_80 : _GEN_2330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2332 = 8'h51 == _match_key_qbytes_3_T ? phv_data_81 : _GEN_2331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2333 = 8'h52 == _match_key_qbytes_3_T ? phv_data_82 : _GEN_2332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2334 = 8'h53 == _match_key_qbytes_3_T ? phv_data_83 : _GEN_2333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2335 = 8'h54 == _match_key_qbytes_3_T ? phv_data_84 : _GEN_2334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2336 = 8'h55 == _match_key_qbytes_3_T ? phv_data_85 : _GEN_2335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2337 = 8'h56 == _match_key_qbytes_3_T ? phv_data_86 : _GEN_2336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2338 = 8'h57 == _match_key_qbytes_3_T ? phv_data_87 : _GEN_2337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2339 = 8'h58 == _match_key_qbytes_3_T ? phv_data_88 : _GEN_2338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2340 = 8'h59 == _match_key_qbytes_3_T ? phv_data_89 : _GEN_2339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2341 = 8'h5a == _match_key_qbytes_3_T ? phv_data_90 : _GEN_2340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2342 = 8'h5b == _match_key_qbytes_3_T ? phv_data_91 : _GEN_2341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2343 = 8'h5c == _match_key_qbytes_3_T ? phv_data_92 : _GEN_2342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2344 = 8'h5d == _match_key_qbytes_3_T ? phv_data_93 : _GEN_2343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2345 = 8'h5e == _match_key_qbytes_3_T ? phv_data_94 : _GEN_2344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2346 = 8'h5f == _match_key_qbytes_3_T ? phv_data_95 : _GEN_2345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2347 = 8'h60 == _match_key_qbytes_3_T ? phv_data_96 : _GEN_2346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2348 = 8'h61 == _match_key_qbytes_3_T ? phv_data_97 : _GEN_2347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2349 = 8'h62 == _match_key_qbytes_3_T ? phv_data_98 : _GEN_2348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2350 = 8'h63 == _match_key_qbytes_3_T ? phv_data_99 : _GEN_2349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2351 = 8'h64 == _match_key_qbytes_3_T ? phv_data_100 : _GEN_2350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2352 = 8'h65 == _match_key_qbytes_3_T ? phv_data_101 : _GEN_2351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2353 = 8'h66 == _match_key_qbytes_3_T ? phv_data_102 : _GEN_2352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2354 = 8'h67 == _match_key_qbytes_3_T ? phv_data_103 : _GEN_2353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2355 = 8'h68 == _match_key_qbytes_3_T ? phv_data_104 : _GEN_2354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2356 = 8'h69 == _match_key_qbytes_3_T ? phv_data_105 : _GEN_2355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2357 = 8'h6a == _match_key_qbytes_3_T ? phv_data_106 : _GEN_2356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2358 = 8'h6b == _match_key_qbytes_3_T ? phv_data_107 : _GEN_2357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2359 = 8'h6c == _match_key_qbytes_3_T ? phv_data_108 : _GEN_2358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2360 = 8'h6d == _match_key_qbytes_3_T ? phv_data_109 : _GEN_2359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2361 = 8'h6e == _match_key_qbytes_3_T ? phv_data_110 : _GEN_2360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2362 = 8'h6f == _match_key_qbytes_3_T ? phv_data_111 : _GEN_2361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2363 = 8'h70 == _match_key_qbytes_3_T ? phv_data_112 : _GEN_2362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2364 = 8'h71 == _match_key_qbytes_3_T ? phv_data_113 : _GEN_2363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2365 = 8'h72 == _match_key_qbytes_3_T ? phv_data_114 : _GEN_2364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2366 = 8'h73 == _match_key_qbytes_3_T ? phv_data_115 : _GEN_2365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2367 = 8'h74 == _match_key_qbytes_3_T ? phv_data_116 : _GEN_2366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2368 = 8'h75 == _match_key_qbytes_3_T ? phv_data_117 : _GEN_2367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2369 = 8'h76 == _match_key_qbytes_3_T ? phv_data_118 : _GEN_2368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2370 = 8'h77 == _match_key_qbytes_3_T ? phv_data_119 : _GEN_2369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2371 = 8'h78 == _match_key_qbytes_3_T ? phv_data_120 : _GEN_2370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2372 = 8'h79 == _match_key_qbytes_3_T ? phv_data_121 : _GEN_2371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2373 = 8'h7a == _match_key_qbytes_3_T ? phv_data_122 : _GEN_2372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2374 = 8'h7b == _match_key_qbytes_3_T ? phv_data_123 : _GEN_2373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2375 = 8'h7c == _match_key_qbytes_3_T ? phv_data_124 : _GEN_2374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2376 = 8'h7d == _match_key_qbytes_3_T ? phv_data_125 : _GEN_2375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2377 = 8'h7e == _match_key_qbytes_3_T ? phv_data_126 : _GEN_2376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2378 = 8'h7f == _match_key_qbytes_3_T ? phv_data_127 : _GEN_2377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2379 = 8'h80 == _match_key_qbytes_3_T ? phv_data_128 : _GEN_2378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2380 = 8'h81 == _match_key_qbytes_3_T ? phv_data_129 : _GEN_2379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2381 = 8'h82 == _match_key_qbytes_3_T ? phv_data_130 : _GEN_2380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2382 = 8'h83 == _match_key_qbytes_3_T ? phv_data_131 : _GEN_2381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2383 = 8'h84 == _match_key_qbytes_3_T ? phv_data_132 : _GEN_2382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2384 = 8'h85 == _match_key_qbytes_3_T ? phv_data_133 : _GEN_2383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2385 = 8'h86 == _match_key_qbytes_3_T ? phv_data_134 : _GEN_2384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2386 = 8'h87 == _match_key_qbytes_3_T ? phv_data_135 : _GEN_2385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2387 = 8'h88 == _match_key_qbytes_3_T ? phv_data_136 : _GEN_2386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2388 = 8'h89 == _match_key_qbytes_3_T ? phv_data_137 : _GEN_2387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2389 = 8'h8a == _match_key_qbytes_3_T ? phv_data_138 : _GEN_2388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2390 = 8'h8b == _match_key_qbytes_3_T ? phv_data_139 : _GEN_2389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2391 = 8'h8c == _match_key_qbytes_3_T ? phv_data_140 : _GEN_2390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2392 = 8'h8d == _match_key_qbytes_3_T ? phv_data_141 : _GEN_2391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2393 = 8'h8e == _match_key_qbytes_3_T ? phv_data_142 : _GEN_2392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2394 = 8'h8f == _match_key_qbytes_3_T ? phv_data_143 : _GEN_2393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2395 = 8'h90 == _match_key_qbytes_3_T ? phv_data_144 : _GEN_2394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2396 = 8'h91 == _match_key_qbytes_3_T ? phv_data_145 : _GEN_2395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2397 = 8'h92 == _match_key_qbytes_3_T ? phv_data_146 : _GEN_2396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2398 = 8'h93 == _match_key_qbytes_3_T ? phv_data_147 : _GEN_2397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2399 = 8'h94 == _match_key_qbytes_3_T ? phv_data_148 : _GEN_2398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2400 = 8'h95 == _match_key_qbytes_3_T ? phv_data_149 : _GEN_2399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2401 = 8'h96 == _match_key_qbytes_3_T ? phv_data_150 : _GEN_2400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2402 = 8'h97 == _match_key_qbytes_3_T ? phv_data_151 : _GEN_2401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2403 = 8'h98 == _match_key_qbytes_3_T ? phv_data_152 : _GEN_2402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2404 = 8'h99 == _match_key_qbytes_3_T ? phv_data_153 : _GEN_2403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2405 = 8'h9a == _match_key_qbytes_3_T ? phv_data_154 : _GEN_2404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2406 = 8'h9b == _match_key_qbytes_3_T ? phv_data_155 : _GEN_2405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2407 = 8'h9c == _match_key_qbytes_3_T ? phv_data_156 : _GEN_2406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2408 = 8'h9d == _match_key_qbytes_3_T ? phv_data_157 : _GEN_2407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2409 = 8'h9e == _match_key_qbytes_3_T ? phv_data_158 : _GEN_2408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2410 = 8'h9f == _match_key_qbytes_3_T ? phv_data_159 : _GEN_2409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2412 = 8'h1 == _match_key_qbytes_3_T_1 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2413 = 8'h2 == _match_key_qbytes_3_T_1 ? phv_data_2 : _GEN_2412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2414 = 8'h3 == _match_key_qbytes_3_T_1 ? phv_data_3 : _GEN_2413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2415 = 8'h4 == _match_key_qbytes_3_T_1 ? phv_data_4 : _GEN_2414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2416 = 8'h5 == _match_key_qbytes_3_T_1 ? phv_data_5 : _GEN_2415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2417 = 8'h6 == _match_key_qbytes_3_T_1 ? phv_data_6 : _GEN_2416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2418 = 8'h7 == _match_key_qbytes_3_T_1 ? phv_data_7 : _GEN_2417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2419 = 8'h8 == _match_key_qbytes_3_T_1 ? phv_data_8 : _GEN_2418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2420 = 8'h9 == _match_key_qbytes_3_T_1 ? phv_data_9 : _GEN_2419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2421 = 8'ha == _match_key_qbytes_3_T_1 ? phv_data_10 : _GEN_2420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2422 = 8'hb == _match_key_qbytes_3_T_1 ? phv_data_11 : _GEN_2421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2423 = 8'hc == _match_key_qbytes_3_T_1 ? phv_data_12 : _GEN_2422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2424 = 8'hd == _match_key_qbytes_3_T_1 ? phv_data_13 : _GEN_2423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2425 = 8'he == _match_key_qbytes_3_T_1 ? phv_data_14 : _GEN_2424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2426 = 8'hf == _match_key_qbytes_3_T_1 ? phv_data_15 : _GEN_2425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2427 = 8'h10 == _match_key_qbytes_3_T_1 ? phv_data_16 : _GEN_2426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2428 = 8'h11 == _match_key_qbytes_3_T_1 ? phv_data_17 : _GEN_2427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2429 = 8'h12 == _match_key_qbytes_3_T_1 ? phv_data_18 : _GEN_2428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2430 = 8'h13 == _match_key_qbytes_3_T_1 ? phv_data_19 : _GEN_2429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2431 = 8'h14 == _match_key_qbytes_3_T_1 ? phv_data_20 : _GEN_2430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2432 = 8'h15 == _match_key_qbytes_3_T_1 ? phv_data_21 : _GEN_2431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2433 = 8'h16 == _match_key_qbytes_3_T_1 ? phv_data_22 : _GEN_2432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2434 = 8'h17 == _match_key_qbytes_3_T_1 ? phv_data_23 : _GEN_2433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2435 = 8'h18 == _match_key_qbytes_3_T_1 ? phv_data_24 : _GEN_2434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2436 = 8'h19 == _match_key_qbytes_3_T_1 ? phv_data_25 : _GEN_2435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2437 = 8'h1a == _match_key_qbytes_3_T_1 ? phv_data_26 : _GEN_2436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2438 = 8'h1b == _match_key_qbytes_3_T_1 ? phv_data_27 : _GEN_2437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2439 = 8'h1c == _match_key_qbytes_3_T_1 ? phv_data_28 : _GEN_2438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2440 = 8'h1d == _match_key_qbytes_3_T_1 ? phv_data_29 : _GEN_2439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2441 = 8'h1e == _match_key_qbytes_3_T_1 ? phv_data_30 : _GEN_2440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2442 = 8'h1f == _match_key_qbytes_3_T_1 ? phv_data_31 : _GEN_2441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2443 = 8'h20 == _match_key_qbytes_3_T_1 ? phv_data_32 : _GEN_2442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2444 = 8'h21 == _match_key_qbytes_3_T_1 ? phv_data_33 : _GEN_2443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2445 = 8'h22 == _match_key_qbytes_3_T_1 ? phv_data_34 : _GEN_2444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2446 = 8'h23 == _match_key_qbytes_3_T_1 ? phv_data_35 : _GEN_2445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2447 = 8'h24 == _match_key_qbytes_3_T_1 ? phv_data_36 : _GEN_2446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2448 = 8'h25 == _match_key_qbytes_3_T_1 ? phv_data_37 : _GEN_2447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2449 = 8'h26 == _match_key_qbytes_3_T_1 ? phv_data_38 : _GEN_2448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2450 = 8'h27 == _match_key_qbytes_3_T_1 ? phv_data_39 : _GEN_2449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2451 = 8'h28 == _match_key_qbytes_3_T_1 ? phv_data_40 : _GEN_2450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2452 = 8'h29 == _match_key_qbytes_3_T_1 ? phv_data_41 : _GEN_2451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2453 = 8'h2a == _match_key_qbytes_3_T_1 ? phv_data_42 : _GEN_2452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2454 = 8'h2b == _match_key_qbytes_3_T_1 ? phv_data_43 : _GEN_2453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2455 = 8'h2c == _match_key_qbytes_3_T_1 ? phv_data_44 : _GEN_2454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2456 = 8'h2d == _match_key_qbytes_3_T_1 ? phv_data_45 : _GEN_2455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2457 = 8'h2e == _match_key_qbytes_3_T_1 ? phv_data_46 : _GEN_2456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2458 = 8'h2f == _match_key_qbytes_3_T_1 ? phv_data_47 : _GEN_2457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2459 = 8'h30 == _match_key_qbytes_3_T_1 ? phv_data_48 : _GEN_2458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2460 = 8'h31 == _match_key_qbytes_3_T_1 ? phv_data_49 : _GEN_2459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2461 = 8'h32 == _match_key_qbytes_3_T_1 ? phv_data_50 : _GEN_2460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2462 = 8'h33 == _match_key_qbytes_3_T_1 ? phv_data_51 : _GEN_2461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2463 = 8'h34 == _match_key_qbytes_3_T_1 ? phv_data_52 : _GEN_2462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2464 = 8'h35 == _match_key_qbytes_3_T_1 ? phv_data_53 : _GEN_2463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2465 = 8'h36 == _match_key_qbytes_3_T_1 ? phv_data_54 : _GEN_2464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2466 = 8'h37 == _match_key_qbytes_3_T_1 ? phv_data_55 : _GEN_2465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2467 = 8'h38 == _match_key_qbytes_3_T_1 ? phv_data_56 : _GEN_2466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2468 = 8'h39 == _match_key_qbytes_3_T_1 ? phv_data_57 : _GEN_2467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2469 = 8'h3a == _match_key_qbytes_3_T_1 ? phv_data_58 : _GEN_2468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2470 = 8'h3b == _match_key_qbytes_3_T_1 ? phv_data_59 : _GEN_2469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2471 = 8'h3c == _match_key_qbytes_3_T_1 ? phv_data_60 : _GEN_2470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2472 = 8'h3d == _match_key_qbytes_3_T_1 ? phv_data_61 : _GEN_2471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2473 = 8'h3e == _match_key_qbytes_3_T_1 ? phv_data_62 : _GEN_2472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2474 = 8'h3f == _match_key_qbytes_3_T_1 ? phv_data_63 : _GEN_2473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2475 = 8'h40 == _match_key_qbytes_3_T_1 ? phv_data_64 : _GEN_2474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2476 = 8'h41 == _match_key_qbytes_3_T_1 ? phv_data_65 : _GEN_2475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2477 = 8'h42 == _match_key_qbytes_3_T_1 ? phv_data_66 : _GEN_2476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2478 = 8'h43 == _match_key_qbytes_3_T_1 ? phv_data_67 : _GEN_2477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2479 = 8'h44 == _match_key_qbytes_3_T_1 ? phv_data_68 : _GEN_2478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2480 = 8'h45 == _match_key_qbytes_3_T_1 ? phv_data_69 : _GEN_2479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2481 = 8'h46 == _match_key_qbytes_3_T_1 ? phv_data_70 : _GEN_2480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2482 = 8'h47 == _match_key_qbytes_3_T_1 ? phv_data_71 : _GEN_2481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2483 = 8'h48 == _match_key_qbytes_3_T_1 ? phv_data_72 : _GEN_2482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2484 = 8'h49 == _match_key_qbytes_3_T_1 ? phv_data_73 : _GEN_2483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2485 = 8'h4a == _match_key_qbytes_3_T_1 ? phv_data_74 : _GEN_2484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2486 = 8'h4b == _match_key_qbytes_3_T_1 ? phv_data_75 : _GEN_2485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2487 = 8'h4c == _match_key_qbytes_3_T_1 ? phv_data_76 : _GEN_2486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2488 = 8'h4d == _match_key_qbytes_3_T_1 ? phv_data_77 : _GEN_2487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2489 = 8'h4e == _match_key_qbytes_3_T_1 ? phv_data_78 : _GEN_2488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2490 = 8'h4f == _match_key_qbytes_3_T_1 ? phv_data_79 : _GEN_2489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2491 = 8'h50 == _match_key_qbytes_3_T_1 ? phv_data_80 : _GEN_2490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2492 = 8'h51 == _match_key_qbytes_3_T_1 ? phv_data_81 : _GEN_2491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2493 = 8'h52 == _match_key_qbytes_3_T_1 ? phv_data_82 : _GEN_2492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2494 = 8'h53 == _match_key_qbytes_3_T_1 ? phv_data_83 : _GEN_2493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2495 = 8'h54 == _match_key_qbytes_3_T_1 ? phv_data_84 : _GEN_2494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2496 = 8'h55 == _match_key_qbytes_3_T_1 ? phv_data_85 : _GEN_2495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2497 = 8'h56 == _match_key_qbytes_3_T_1 ? phv_data_86 : _GEN_2496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2498 = 8'h57 == _match_key_qbytes_3_T_1 ? phv_data_87 : _GEN_2497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2499 = 8'h58 == _match_key_qbytes_3_T_1 ? phv_data_88 : _GEN_2498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2500 = 8'h59 == _match_key_qbytes_3_T_1 ? phv_data_89 : _GEN_2499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2501 = 8'h5a == _match_key_qbytes_3_T_1 ? phv_data_90 : _GEN_2500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2502 = 8'h5b == _match_key_qbytes_3_T_1 ? phv_data_91 : _GEN_2501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2503 = 8'h5c == _match_key_qbytes_3_T_1 ? phv_data_92 : _GEN_2502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2504 = 8'h5d == _match_key_qbytes_3_T_1 ? phv_data_93 : _GEN_2503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2505 = 8'h5e == _match_key_qbytes_3_T_1 ? phv_data_94 : _GEN_2504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2506 = 8'h5f == _match_key_qbytes_3_T_1 ? phv_data_95 : _GEN_2505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2507 = 8'h60 == _match_key_qbytes_3_T_1 ? phv_data_96 : _GEN_2506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2508 = 8'h61 == _match_key_qbytes_3_T_1 ? phv_data_97 : _GEN_2507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2509 = 8'h62 == _match_key_qbytes_3_T_1 ? phv_data_98 : _GEN_2508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2510 = 8'h63 == _match_key_qbytes_3_T_1 ? phv_data_99 : _GEN_2509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2511 = 8'h64 == _match_key_qbytes_3_T_1 ? phv_data_100 : _GEN_2510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2512 = 8'h65 == _match_key_qbytes_3_T_1 ? phv_data_101 : _GEN_2511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2513 = 8'h66 == _match_key_qbytes_3_T_1 ? phv_data_102 : _GEN_2512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2514 = 8'h67 == _match_key_qbytes_3_T_1 ? phv_data_103 : _GEN_2513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2515 = 8'h68 == _match_key_qbytes_3_T_1 ? phv_data_104 : _GEN_2514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2516 = 8'h69 == _match_key_qbytes_3_T_1 ? phv_data_105 : _GEN_2515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2517 = 8'h6a == _match_key_qbytes_3_T_1 ? phv_data_106 : _GEN_2516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2518 = 8'h6b == _match_key_qbytes_3_T_1 ? phv_data_107 : _GEN_2517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2519 = 8'h6c == _match_key_qbytes_3_T_1 ? phv_data_108 : _GEN_2518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2520 = 8'h6d == _match_key_qbytes_3_T_1 ? phv_data_109 : _GEN_2519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2521 = 8'h6e == _match_key_qbytes_3_T_1 ? phv_data_110 : _GEN_2520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2522 = 8'h6f == _match_key_qbytes_3_T_1 ? phv_data_111 : _GEN_2521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2523 = 8'h70 == _match_key_qbytes_3_T_1 ? phv_data_112 : _GEN_2522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2524 = 8'h71 == _match_key_qbytes_3_T_1 ? phv_data_113 : _GEN_2523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2525 = 8'h72 == _match_key_qbytes_3_T_1 ? phv_data_114 : _GEN_2524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2526 = 8'h73 == _match_key_qbytes_3_T_1 ? phv_data_115 : _GEN_2525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2527 = 8'h74 == _match_key_qbytes_3_T_1 ? phv_data_116 : _GEN_2526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2528 = 8'h75 == _match_key_qbytes_3_T_1 ? phv_data_117 : _GEN_2527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2529 = 8'h76 == _match_key_qbytes_3_T_1 ? phv_data_118 : _GEN_2528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2530 = 8'h77 == _match_key_qbytes_3_T_1 ? phv_data_119 : _GEN_2529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2531 = 8'h78 == _match_key_qbytes_3_T_1 ? phv_data_120 : _GEN_2530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2532 = 8'h79 == _match_key_qbytes_3_T_1 ? phv_data_121 : _GEN_2531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2533 = 8'h7a == _match_key_qbytes_3_T_1 ? phv_data_122 : _GEN_2532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2534 = 8'h7b == _match_key_qbytes_3_T_1 ? phv_data_123 : _GEN_2533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2535 = 8'h7c == _match_key_qbytes_3_T_1 ? phv_data_124 : _GEN_2534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2536 = 8'h7d == _match_key_qbytes_3_T_1 ? phv_data_125 : _GEN_2535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2537 = 8'h7e == _match_key_qbytes_3_T_1 ? phv_data_126 : _GEN_2536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2538 = 8'h7f == _match_key_qbytes_3_T_1 ? phv_data_127 : _GEN_2537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2539 = 8'h80 == _match_key_qbytes_3_T_1 ? phv_data_128 : _GEN_2538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2540 = 8'h81 == _match_key_qbytes_3_T_1 ? phv_data_129 : _GEN_2539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2541 = 8'h82 == _match_key_qbytes_3_T_1 ? phv_data_130 : _GEN_2540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2542 = 8'h83 == _match_key_qbytes_3_T_1 ? phv_data_131 : _GEN_2541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2543 = 8'h84 == _match_key_qbytes_3_T_1 ? phv_data_132 : _GEN_2542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2544 = 8'h85 == _match_key_qbytes_3_T_1 ? phv_data_133 : _GEN_2543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2545 = 8'h86 == _match_key_qbytes_3_T_1 ? phv_data_134 : _GEN_2544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2546 = 8'h87 == _match_key_qbytes_3_T_1 ? phv_data_135 : _GEN_2545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2547 = 8'h88 == _match_key_qbytes_3_T_1 ? phv_data_136 : _GEN_2546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2548 = 8'h89 == _match_key_qbytes_3_T_1 ? phv_data_137 : _GEN_2547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2549 = 8'h8a == _match_key_qbytes_3_T_1 ? phv_data_138 : _GEN_2548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2550 = 8'h8b == _match_key_qbytes_3_T_1 ? phv_data_139 : _GEN_2549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2551 = 8'h8c == _match_key_qbytes_3_T_1 ? phv_data_140 : _GEN_2550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2552 = 8'h8d == _match_key_qbytes_3_T_1 ? phv_data_141 : _GEN_2551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2553 = 8'h8e == _match_key_qbytes_3_T_1 ? phv_data_142 : _GEN_2552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2554 = 8'h8f == _match_key_qbytes_3_T_1 ? phv_data_143 : _GEN_2553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2555 = 8'h90 == _match_key_qbytes_3_T_1 ? phv_data_144 : _GEN_2554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2556 = 8'h91 == _match_key_qbytes_3_T_1 ? phv_data_145 : _GEN_2555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2557 = 8'h92 == _match_key_qbytes_3_T_1 ? phv_data_146 : _GEN_2556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2558 = 8'h93 == _match_key_qbytes_3_T_1 ? phv_data_147 : _GEN_2557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2559 = 8'h94 == _match_key_qbytes_3_T_1 ? phv_data_148 : _GEN_2558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2560 = 8'h95 == _match_key_qbytes_3_T_1 ? phv_data_149 : _GEN_2559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2561 = 8'h96 == _match_key_qbytes_3_T_1 ? phv_data_150 : _GEN_2560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2562 = 8'h97 == _match_key_qbytes_3_T_1 ? phv_data_151 : _GEN_2561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2563 = 8'h98 == _match_key_qbytes_3_T_1 ? phv_data_152 : _GEN_2562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2564 = 8'h99 == _match_key_qbytes_3_T_1 ? phv_data_153 : _GEN_2563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2565 = 8'h9a == _match_key_qbytes_3_T_1 ? phv_data_154 : _GEN_2564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2566 = 8'h9b == _match_key_qbytes_3_T_1 ? phv_data_155 : _GEN_2565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2567 = 8'h9c == _match_key_qbytes_3_T_1 ? phv_data_156 : _GEN_2566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2568 = 8'h9d == _match_key_qbytes_3_T_1 ? phv_data_157 : _GEN_2567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2569 = 8'h9e == _match_key_qbytes_3_T_1 ? phv_data_158 : _GEN_2568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2570 = 8'h9f == _match_key_qbytes_3_T_1 ? phv_data_159 : _GEN_2569; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [31:0] _match_key_qbytes_3_T_3 = {_GEN_2410,_GEN_2570,_GEN_2090,_GEN_2250}; // @[Cat.scala 30:58]
  wire [31:0] match_key_qbytes_3 = local_offset_3 < end_offset ? _match_key_qbytes_3_T_3 : 32'h0; // @[matcher.scala 88:54 matcher.scala 89:45 matcher.scala 97:45]
  wire [7:0] local_offset_4 = 8'h10 + read_key_offset; // @[matcher.scala 87:77]
  wire [5:0] match_key_qbytes_4_hi = local_offset_4[7:2]; // @[matcher.scala 91:54]
  wire [7:0] _match_key_qbytes_4_T = {match_key_qbytes_4_hi,2'h3}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_4_T_1 = {match_key_qbytes_4_hi,2'h2}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_4_T_2 = {match_key_qbytes_4_hi,2'h1}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_2573 = 8'h1 == _match_key_qbytes_4_T_2 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2574 = 8'h2 == _match_key_qbytes_4_T_2 ? phv_data_2 : _GEN_2573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2575 = 8'h3 == _match_key_qbytes_4_T_2 ? phv_data_3 : _GEN_2574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2576 = 8'h4 == _match_key_qbytes_4_T_2 ? phv_data_4 : _GEN_2575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2577 = 8'h5 == _match_key_qbytes_4_T_2 ? phv_data_5 : _GEN_2576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2578 = 8'h6 == _match_key_qbytes_4_T_2 ? phv_data_6 : _GEN_2577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2579 = 8'h7 == _match_key_qbytes_4_T_2 ? phv_data_7 : _GEN_2578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2580 = 8'h8 == _match_key_qbytes_4_T_2 ? phv_data_8 : _GEN_2579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2581 = 8'h9 == _match_key_qbytes_4_T_2 ? phv_data_9 : _GEN_2580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2582 = 8'ha == _match_key_qbytes_4_T_2 ? phv_data_10 : _GEN_2581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2583 = 8'hb == _match_key_qbytes_4_T_2 ? phv_data_11 : _GEN_2582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2584 = 8'hc == _match_key_qbytes_4_T_2 ? phv_data_12 : _GEN_2583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2585 = 8'hd == _match_key_qbytes_4_T_2 ? phv_data_13 : _GEN_2584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2586 = 8'he == _match_key_qbytes_4_T_2 ? phv_data_14 : _GEN_2585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2587 = 8'hf == _match_key_qbytes_4_T_2 ? phv_data_15 : _GEN_2586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2588 = 8'h10 == _match_key_qbytes_4_T_2 ? phv_data_16 : _GEN_2587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2589 = 8'h11 == _match_key_qbytes_4_T_2 ? phv_data_17 : _GEN_2588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2590 = 8'h12 == _match_key_qbytes_4_T_2 ? phv_data_18 : _GEN_2589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2591 = 8'h13 == _match_key_qbytes_4_T_2 ? phv_data_19 : _GEN_2590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2592 = 8'h14 == _match_key_qbytes_4_T_2 ? phv_data_20 : _GEN_2591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2593 = 8'h15 == _match_key_qbytes_4_T_2 ? phv_data_21 : _GEN_2592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2594 = 8'h16 == _match_key_qbytes_4_T_2 ? phv_data_22 : _GEN_2593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2595 = 8'h17 == _match_key_qbytes_4_T_2 ? phv_data_23 : _GEN_2594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2596 = 8'h18 == _match_key_qbytes_4_T_2 ? phv_data_24 : _GEN_2595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2597 = 8'h19 == _match_key_qbytes_4_T_2 ? phv_data_25 : _GEN_2596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2598 = 8'h1a == _match_key_qbytes_4_T_2 ? phv_data_26 : _GEN_2597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2599 = 8'h1b == _match_key_qbytes_4_T_2 ? phv_data_27 : _GEN_2598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2600 = 8'h1c == _match_key_qbytes_4_T_2 ? phv_data_28 : _GEN_2599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2601 = 8'h1d == _match_key_qbytes_4_T_2 ? phv_data_29 : _GEN_2600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2602 = 8'h1e == _match_key_qbytes_4_T_2 ? phv_data_30 : _GEN_2601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2603 = 8'h1f == _match_key_qbytes_4_T_2 ? phv_data_31 : _GEN_2602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2604 = 8'h20 == _match_key_qbytes_4_T_2 ? phv_data_32 : _GEN_2603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2605 = 8'h21 == _match_key_qbytes_4_T_2 ? phv_data_33 : _GEN_2604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2606 = 8'h22 == _match_key_qbytes_4_T_2 ? phv_data_34 : _GEN_2605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2607 = 8'h23 == _match_key_qbytes_4_T_2 ? phv_data_35 : _GEN_2606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2608 = 8'h24 == _match_key_qbytes_4_T_2 ? phv_data_36 : _GEN_2607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2609 = 8'h25 == _match_key_qbytes_4_T_2 ? phv_data_37 : _GEN_2608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2610 = 8'h26 == _match_key_qbytes_4_T_2 ? phv_data_38 : _GEN_2609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2611 = 8'h27 == _match_key_qbytes_4_T_2 ? phv_data_39 : _GEN_2610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2612 = 8'h28 == _match_key_qbytes_4_T_2 ? phv_data_40 : _GEN_2611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2613 = 8'h29 == _match_key_qbytes_4_T_2 ? phv_data_41 : _GEN_2612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2614 = 8'h2a == _match_key_qbytes_4_T_2 ? phv_data_42 : _GEN_2613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2615 = 8'h2b == _match_key_qbytes_4_T_2 ? phv_data_43 : _GEN_2614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2616 = 8'h2c == _match_key_qbytes_4_T_2 ? phv_data_44 : _GEN_2615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2617 = 8'h2d == _match_key_qbytes_4_T_2 ? phv_data_45 : _GEN_2616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2618 = 8'h2e == _match_key_qbytes_4_T_2 ? phv_data_46 : _GEN_2617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2619 = 8'h2f == _match_key_qbytes_4_T_2 ? phv_data_47 : _GEN_2618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2620 = 8'h30 == _match_key_qbytes_4_T_2 ? phv_data_48 : _GEN_2619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2621 = 8'h31 == _match_key_qbytes_4_T_2 ? phv_data_49 : _GEN_2620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2622 = 8'h32 == _match_key_qbytes_4_T_2 ? phv_data_50 : _GEN_2621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2623 = 8'h33 == _match_key_qbytes_4_T_2 ? phv_data_51 : _GEN_2622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2624 = 8'h34 == _match_key_qbytes_4_T_2 ? phv_data_52 : _GEN_2623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2625 = 8'h35 == _match_key_qbytes_4_T_2 ? phv_data_53 : _GEN_2624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2626 = 8'h36 == _match_key_qbytes_4_T_2 ? phv_data_54 : _GEN_2625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2627 = 8'h37 == _match_key_qbytes_4_T_2 ? phv_data_55 : _GEN_2626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2628 = 8'h38 == _match_key_qbytes_4_T_2 ? phv_data_56 : _GEN_2627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2629 = 8'h39 == _match_key_qbytes_4_T_2 ? phv_data_57 : _GEN_2628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2630 = 8'h3a == _match_key_qbytes_4_T_2 ? phv_data_58 : _GEN_2629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2631 = 8'h3b == _match_key_qbytes_4_T_2 ? phv_data_59 : _GEN_2630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2632 = 8'h3c == _match_key_qbytes_4_T_2 ? phv_data_60 : _GEN_2631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2633 = 8'h3d == _match_key_qbytes_4_T_2 ? phv_data_61 : _GEN_2632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2634 = 8'h3e == _match_key_qbytes_4_T_2 ? phv_data_62 : _GEN_2633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2635 = 8'h3f == _match_key_qbytes_4_T_2 ? phv_data_63 : _GEN_2634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2636 = 8'h40 == _match_key_qbytes_4_T_2 ? phv_data_64 : _GEN_2635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2637 = 8'h41 == _match_key_qbytes_4_T_2 ? phv_data_65 : _GEN_2636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2638 = 8'h42 == _match_key_qbytes_4_T_2 ? phv_data_66 : _GEN_2637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2639 = 8'h43 == _match_key_qbytes_4_T_2 ? phv_data_67 : _GEN_2638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2640 = 8'h44 == _match_key_qbytes_4_T_2 ? phv_data_68 : _GEN_2639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2641 = 8'h45 == _match_key_qbytes_4_T_2 ? phv_data_69 : _GEN_2640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2642 = 8'h46 == _match_key_qbytes_4_T_2 ? phv_data_70 : _GEN_2641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2643 = 8'h47 == _match_key_qbytes_4_T_2 ? phv_data_71 : _GEN_2642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2644 = 8'h48 == _match_key_qbytes_4_T_2 ? phv_data_72 : _GEN_2643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2645 = 8'h49 == _match_key_qbytes_4_T_2 ? phv_data_73 : _GEN_2644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2646 = 8'h4a == _match_key_qbytes_4_T_2 ? phv_data_74 : _GEN_2645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2647 = 8'h4b == _match_key_qbytes_4_T_2 ? phv_data_75 : _GEN_2646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2648 = 8'h4c == _match_key_qbytes_4_T_2 ? phv_data_76 : _GEN_2647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2649 = 8'h4d == _match_key_qbytes_4_T_2 ? phv_data_77 : _GEN_2648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2650 = 8'h4e == _match_key_qbytes_4_T_2 ? phv_data_78 : _GEN_2649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2651 = 8'h4f == _match_key_qbytes_4_T_2 ? phv_data_79 : _GEN_2650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2652 = 8'h50 == _match_key_qbytes_4_T_2 ? phv_data_80 : _GEN_2651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2653 = 8'h51 == _match_key_qbytes_4_T_2 ? phv_data_81 : _GEN_2652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2654 = 8'h52 == _match_key_qbytes_4_T_2 ? phv_data_82 : _GEN_2653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2655 = 8'h53 == _match_key_qbytes_4_T_2 ? phv_data_83 : _GEN_2654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2656 = 8'h54 == _match_key_qbytes_4_T_2 ? phv_data_84 : _GEN_2655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2657 = 8'h55 == _match_key_qbytes_4_T_2 ? phv_data_85 : _GEN_2656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2658 = 8'h56 == _match_key_qbytes_4_T_2 ? phv_data_86 : _GEN_2657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2659 = 8'h57 == _match_key_qbytes_4_T_2 ? phv_data_87 : _GEN_2658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2660 = 8'h58 == _match_key_qbytes_4_T_2 ? phv_data_88 : _GEN_2659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2661 = 8'h59 == _match_key_qbytes_4_T_2 ? phv_data_89 : _GEN_2660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2662 = 8'h5a == _match_key_qbytes_4_T_2 ? phv_data_90 : _GEN_2661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2663 = 8'h5b == _match_key_qbytes_4_T_2 ? phv_data_91 : _GEN_2662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2664 = 8'h5c == _match_key_qbytes_4_T_2 ? phv_data_92 : _GEN_2663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2665 = 8'h5d == _match_key_qbytes_4_T_2 ? phv_data_93 : _GEN_2664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2666 = 8'h5e == _match_key_qbytes_4_T_2 ? phv_data_94 : _GEN_2665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2667 = 8'h5f == _match_key_qbytes_4_T_2 ? phv_data_95 : _GEN_2666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2668 = 8'h60 == _match_key_qbytes_4_T_2 ? phv_data_96 : _GEN_2667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2669 = 8'h61 == _match_key_qbytes_4_T_2 ? phv_data_97 : _GEN_2668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2670 = 8'h62 == _match_key_qbytes_4_T_2 ? phv_data_98 : _GEN_2669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2671 = 8'h63 == _match_key_qbytes_4_T_2 ? phv_data_99 : _GEN_2670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2672 = 8'h64 == _match_key_qbytes_4_T_2 ? phv_data_100 : _GEN_2671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2673 = 8'h65 == _match_key_qbytes_4_T_2 ? phv_data_101 : _GEN_2672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2674 = 8'h66 == _match_key_qbytes_4_T_2 ? phv_data_102 : _GEN_2673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2675 = 8'h67 == _match_key_qbytes_4_T_2 ? phv_data_103 : _GEN_2674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2676 = 8'h68 == _match_key_qbytes_4_T_2 ? phv_data_104 : _GEN_2675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2677 = 8'h69 == _match_key_qbytes_4_T_2 ? phv_data_105 : _GEN_2676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2678 = 8'h6a == _match_key_qbytes_4_T_2 ? phv_data_106 : _GEN_2677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2679 = 8'h6b == _match_key_qbytes_4_T_2 ? phv_data_107 : _GEN_2678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2680 = 8'h6c == _match_key_qbytes_4_T_2 ? phv_data_108 : _GEN_2679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2681 = 8'h6d == _match_key_qbytes_4_T_2 ? phv_data_109 : _GEN_2680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2682 = 8'h6e == _match_key_qbytes_4_T_2 ? phv_data_110 : _GEN_2681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2683 = 8'h6f == _match_key_qbytes_4_T_2 ? phv_data_111 : _GEN_2682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2684 = 8'h70 == _match_key_qbytes_4_T_2 ? phv_data_112 : _GEN_2683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2685 = 8'h71 == _match_key_qbytes_4_T_2 ? phv_data_113 : _GEN_2684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2686 = 8'h72 == _match_key_qbytes_4_T_2 ? phv_data_114 : _GEN_2685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2687 = 8'h73 == _match_key_qbytes_4_T_2 ? phv_data_115 : _GEN_2686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2688 = 8'h74 == _match_key_qbytes_4_T_2 ? phv_data_116 : _GEN_2687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2689 = 8'h75 == _match_key_qbytes_4_T_2 ? phv_data_117 : _GEN_2688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2690 = 8'h76 == _match_key_qbytes_4_T_2 ? phv_data_118 : _GEN_2689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2691 = 8'h77 == _match_key_qbytes_4_T_2 ? phv_data_119 : _GEN_2690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2692 = 8'h78 == _match_key_qbytes_4_T_2 ? phv_data_120 : _GEN_2691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2693 = 8'h79 == _match_key_qbytes_4_T_2 ? phv_data_121 : _GEN_2692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2694 = 8'h7a == _match_key_qbytes_4_T_2 ? phv_data_122 : _GEN_2693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2695 = 8'h7b == _match_key_qbytes_4_T_2 ? phv_data_123 : _GEN_2694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2696 = 8'h7c == _match_key_qbytes_4_T_2 ? phv_data_124 : _GEN_2695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2697 = 8'h7d == _match_key_qbytes_4_T_2 ? phv_data_125 : _GEN_2696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2698 = 8'h7e == _match_key_qbytes_4_T_2 ? phv_data_126 : _GEN_2697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2699 = 8'h7f == _match_key_qbytes_4_T_2 ? phv_data_127 : _GEN_2698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2700 = 8'h80 == _match_key_qbytes_4_T_2 ? phv_data_128 : _GEN_2699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2701 = 8'h81 == _match_key_qbytes_4_T_2 ? phv_data_129 : _GEN_2700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2702 = 8'h82 == _match_key_qbytes_4_T_2 ? phv_data_130 : _GEN_2701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2703 = 8'h83 == _match_key_qbytes_4_T_2 ? phv_data_131 : _GEN_2702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2704 = 8'h84 == _match_key_qbytes_4_T_2 ? phv_data_132 : _GEN_2703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2705 = 8'h85 == _match_key_qbytes_4_T_2 ? phv_data_133 : _GEN_2704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2706 = 8'h86 == _match_key_qbytes_4_T_2 ? phv_data_134 : _GEN_2705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2707 = 8'h87 == _match_key_qbytes_4_T_2 ? phv_data_135 : _GEN_2706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2708 = 8'h88 == _match_key_qbytes_4_T_2 ? phv_data_136 : _GEN_2707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2709 = 8'h89 == _match_key_qbytes_4_T_2 ? phv_data_137 : _GEN_2708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2710 = 8'h8a == _match_key_qbytes_4_T_2 ? phv_data_138 : _GEN_2709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2711 = 8'h8b == _match_key_qbytes_4_T_2 ? phv_data_139 : _GEN_2710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2712 = 8'h8c == _match_key_qbytes_4_T_2 ? phv_data_140 : _GEN_2711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2713 = 8'h8d == _match_key_qbytes_4_T_2 ? phv_data_141 : _GEN_2712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2714 = 8'h8e == _match_key_qbytes_4_T_2 ? phv_data_142 : _GEN_2713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2715 = 8'h8f == _match_key_qbytes_4_T_2 ? phv_data_143 : _GEN_2714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2716 = 8'h90 == _match_key_qbytes_4_T_2 ? phv_data_144 : _GEN_2715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2717 = 8'h91 == _match_key_qbytes_4_T_2 ? phv_data_145 : _GEN_2716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2718 = 8'h92 == _match_key_qbytes_4_T_2 ? phv_data_146 : _GEN_2717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2719 = 8'h93 == _match_key_qbytes_4_T_2 ? phv_data_147 : _GEN_2718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2720 = 8'h94 == _match_key_qbytes_4_T_2 ? phv_data_148 : _GEN_2719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2721 = 8'h95 == _match_key_qbytes_4_T_2 ? phv_data_149 : _GEN_2720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2722 = 8'h96 == _match_key_qbytes_4_T_2 ? phv_data_150 : _GEN_2721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2723 = 8'h97 == _match_key_qbytes_4_T_2 ? phv_data_151 : _GEN_2722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2724 = 8'h98 == _match_key_qbytes_4_T_2 ? phv_data_152 : _GEN_2723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2725 = 8'h99 == _match_key_qbytes_4_T_2 ? phv_data_153 : _GEN_2724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2726 = 8'h9a == _match_key_qbytes_4_T_2 ? phv_data_154 : _GEN_2725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2727 = 8'h9b == _match_key_qbytes_4_T_2 ? phv_data_155 : _GEN_2726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2728 = 8'h9c == _match_key_qbytes_4_T_2 ? phv_data_156 : _GEN_2727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2729 = 8'h9d == _match_key_qbytes_4_T_2 ? phv_data_157 : _GEN_2728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2730 = 8'h9e == _match_key_qbytes_4_T_2 ? phv_data_158 : _GEN_2729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2731 = 8'h9f == _match_key_qbytes_4_T_2 ? phv_data_159 : _GEN_2730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2733 = 8'h1 == local_offset_4 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2734 = 8'h2 == local_offset_4 ? phv_data_2 : _GEN_2733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2735 = 8'h3 == local_offset_4 ? phv_data_3 : _GEN_2734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2736 = 8'h4 == local_offset_4 ? phv_data_4 : _GEN_2735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2737 = 8'h5 == local_offset_4 ? phv_data_5 : _GEN_2736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2738 = 8'h6 == local_offset_4 ? phv_data_6 : _GEN_2737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2739 = 8'h7 == local_offset_4 ? phv_data_7 : _GEN_2738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2740 = 8'h8 == local_offset_4 ? phv_data_8 : _GEN_2739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2741 = 8'h9 == local_offset_4 ? phv_data_9 : _GEN_2740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2742 = 8'ha == local_offset_4 ? phv_data_10 : _GEN_2741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2743 = 8'hb == local_offset_4 ? phv_data_11 : _GEN_2742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2744 = 8'hc == local_offset_4 ? phv_data_12 : _GEN_2743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2745 = 8'hd == local_offset_4 ? phv_data_13 : _GEN_2744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2746 = 8'he == local_offset_4 ? phv_data_14 : _GEN_2745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2747 = 8'hf == local_offset_4 ? phv_data_15 : _GEN_2746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2748 = 8'h10 == local_offset_4 ? phv_data_16 : _GEN_2747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2749 = 8'h11 == local_offset_4 ? phv_data_17 : _GEN_2748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2750 = 8'h12 == local_offset_4 ? phv_data_18 : _GEN_2749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2751 = 8'h13 == local_offset_4 ? phv_data_19 : _GEN_2750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2752 = 8'h14 == local_offset_4 ? phv_data_20 : _GEN_2751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2753 = 8'h15 == local_offset_4 ? phv_data_21 : _GEN_2752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2754 = 8'h16 == local_offset_4 ? phv_data_22 : _GEN_2753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2755 = 8'h17 == local_offset_4 ? phv_data_23 : _GEN_2754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2756 = 8'h18 == local_offset_4 ? phv_data_24 : _GEN_2755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2757 = 8'h19 == local_offset_4 ? phv_data_25 : _GEN_2756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2758 = 8'h1a == local_offset_4 ? phv_data_26 : _GEN_2757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2759 = 8'h1b == local_offset_4 ? phv_data_27 : _GEN_2758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2760 = 8'h1c == local_offset_4 ? phv_data_28 : _GEN_2759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2761 = 8'h1d == local_offset_4 ? phv_data_29 : _GEN_2760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2762 = 8'h1e == local_offset_4 ? phv_data_30 : _GEN_2761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2763 = 8'h1f == local_offset_4 ? phv_data_31 : _GEN_2762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2764 = 8'h20 == local_offset_4 ? phv_data_32 : _GEN_2763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2765 = 8'h21 == local_offset_4 ? phv_data_33 : _GEN_2764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2766 = 8'h22 == local_offset_4 ? phv_data_34 : _GEN_2765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2767 = 8'h23 == local_offset_4 ? phv_data_35 : _GEN_2766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2768 = 8'h24 == local_offset_4 ? phv_data_36 : _GEN_2767; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2769 = 8'h25 == local_offset_4 ? phv_data_37 : _GEN_2768; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2770 = 8'h26 == local_offset_4 ? phv_data_38 : _GEN_2769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2771 = 8'h27 == local_offset_4 ? phv_data_39 : _GEN_2770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2772 = 8'h28 == local_offset_4 ? phv_data_40 : _GEN_2771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2773 = 8'h29 == local_offset_4 ? phv_data_41 : _GEN_2772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2774 = 8'h2a == local_offset_4 ? phv_data_42 : _GEN_2773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2775 = 8'h2b == local_offset_4 ? phv_data_43 : _GEN_2774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2776 = 8'h2c == local_offset_4 ? phv_data_44 : _GEN_2775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2777 = 8'h2d == local_offset_4 ? phv_data_45 : _GEN_2776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2778 = 8'h2e == local_offset_4 ? phv_data_46 : _GEN_2777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2779 = 8'h2f == local_offset_4 ? phv_data_47 : _GEN_2778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2780 = 8'h30 == local_offset_4 ? phv_data_48 : _GEN_2779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2781 = 8'h31 == local_offset_4 ? phv_data_49 : _GEN_2780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2782 = 8'h32 == local_offset_4 ? phv_data_50 : _GEN_2781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2783 = 8'h33 == local_offset_4 ? phv_data_51 : _GEN_2782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2784 = 8'h34 == local_offset_4 ? phv_data_52 : _GEN_2783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2785 = 8'h35 == local_offset_4 ? phv_data_53 : _GEN_2784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2786 = 8'h36 == local_offset_4 ? phv_data_54 : _GEN_2785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2787 = 8'h37 == local_offset_4 ? phv_data_55 : _GEN_2786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2788 = 8'h38 == local_offset_4 ? phv_data_56 : _GEN_2787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2789 = 8'h39 == local_offset_4 ? phv_data_57 : _GEN_2788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2790 = 8'h3a == local_offset_4 ? phv_data_58 : _GEN_2789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2791 = 8'h3b == local_offset_4 ? phv_data_59 : _GEN_2790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2792 = 8'h3c == local_offset_4 ? phv_data_60 : _GEN_2791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2793 = 8'h3d == local_offset_4 ? phv_data_61 : _GEN_2792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2794 = 8'h3e == local_offset_4 ? phv_data_62 : _GEN_2793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2795 = 8'h3f == local_offset_4 ? phv_data_63 : _GEN_2794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2796 = 8'h40 == local_offset_4 ? phv_data_64 : _GEN_2795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2797 = 8'h41 == local_offset_4 ? phv_data_65 : _GEN_2796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2798 = 8'h42 == local_offset_4 ? phv_data_66 : _GEN_2797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2799 = 8'h43 == local_offset_4 ? phv_data_67 : _GEN_2798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2800 = 8'h44 == local_offset_4 ? phv_data_68 : _GEN_2799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2801 = 8'h45 == local_offset_4 ? phv_data_69 : _GEN_2800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2802 = 8'h46 == local_offset_4 ? phv_data_70 : _GEN_2801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2803 = 8'h47 == local_offset_4 ? phv_data_71 : _GEN_2802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2804 = 8'h48 == local_offset_4 ? phv_data_72 : _GEN_2803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2805 = 8'h49 == local_offset_4 ? phv_data_73 : _GEN_2804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2806 = 8'h4a == local_offset_4 ? phv_data_74 : _GEN_2805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2807 = 8'h4b == local_offset_4 ? phv_data_75 : _GEN_2806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2808 = 8'h4c == local_offset_4 ? phv_data_76 : _GEN_2807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2809 = 8'h4d == local_offset_4 ? phv_data_77 : _GEN_2808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2810 = 8'h4e == local_offset_4 ? phv_data_78 : _GEN_2809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2811 = 8'h4f == local_offset_4 ? phv_data_79 : _GEN_2810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2812 = 8'h50 == local_offset_4 ? phv_data_80 : _GEN_2811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2813 = 8'h51 == local_offset_4 ? phv_data_81 : _GEN_2812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2814 = 8'h52 == local_offset_4 ? phv_data_82 : _GEN_2813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2815 = 8'h53 == local_offset_4 ? phv_data_83 : _GEN_2814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2816 = 8'h54 == local_offset_4 ? phv_data_84 : _GEN_2815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2817 = 8'h55 == local_offset_4 ? phv_data_85 : _GEN_2816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2818 = 8'h56 == local_offset_4 ? phv_data_86 : _GEN_2817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2819 = 8'h57 == local_offset_4 ? phv_data_87 : _GEN_2818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2820 = 8'h58 == local_offset_4 ? phv_data_88 : _GEN_2819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2821 = 8'h59 == local_offset_4 ? phv_data_89 : _GEN_2820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2822 = 8'h5a == local_offset_4 ? phv_data_90 : _GEN_2821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2823 = 8'h5b == local_offset_4 ? phv_data_91 : _GEN_2822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2824 = 8'h5c == local_offset_4 ? phv_data_92 : _GEN_2823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2825 = 8'h5d == local_offset_4 ? phv_data_93 : _GEN_2824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2826 = 8'h5e == local_offset_4 ? phv_data_94 : _GEN_2825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2827 = 8'h5f == local_offset_4 ? phv_data_95 : _GEN_2826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2828 = 8'h60 == local_offset_4 ? phv_data_96 : _GEN_2827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2829 = 8'h61 == local_offset_4 ? phv_data_97 : _GEN_2828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2830 = 8'h62 == local_offset_4 ? phv_data_98 : _GEN_2829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2831 = 8'h63 == local_offset_4 ? phv_data_99 : _GEN_2830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2832 = 8'h64 == local_offset_4 ? phv_data_100 : _GEN_2831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2833 = 8'h65 == local_offset_4 ? phv_data_101 : _GEN_2832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2834 = 8'h66 == local_offset_4 ? phv_data_102 : _GEN_2833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2835 = 8'h67 == local_offset_4 ? phv_data_103 : _GEN_2834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2836 = 8'h68 == local_offset_4 ? phv_data_104 : _GEN_2835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2837 = 8'h69 == local_offset_4 ? phv_data_105 : _GEN_2836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2838 = 8'h6a == local_offset_4 ? phv_data_106 : _GEN_2837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2839 = 8'h6b == local_offset_4 ? phv_data_107 : _GEN_2838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2840 = 8'h6c == local_offset_4 ? phv_data_108 : _GEN_2839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2841 = 8'h6d == local_offset_4 ? phv_data_109 : _GEN_2840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2842 = 8'h6e == local_offset_4 ? phv_data_110 : _GEN_2841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2843 = 8'h6f == local_offset_4 ? phv_data_111 : _GEN_2842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2844 = 8'h70 == local_offset_4 ? phv_data_112 : _GEN_2843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2845 = 8'h71 == local_offset_4 ? phv_data_113 : _GEN_2844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2846 = 8'h72 == local_offset_4 ? phv_data_114 : _GEN_2845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2847 = 8'h73 == local_offset_4 ? phv_data_115 : _GEN_2846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2848 = 8'h74 == local_offset_4 ? phv_data_116 : _GEN_2847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2849 = 8'h75 == local_offset_4 ? phv_data_117 : _GEN_2848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2850 = 8'h76 == local_offset_4 ? phv_data_118 : _GEN_2849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2851 = 8'h77 == local_offset_4 ? phv_data_119 : _GEN_2850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2852 = 8'h78 == local_offset_4 ? phv_data_120 : _GEN_2851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2853 = 8'h79 == local_offset_4 ? phv_data_121 : _GEN_2852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2854 = 8'h7a == local_offset_4 ? phv_data_122 : _GEN_2853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2855 = 8'h7b == local_offset_4 ? phv_data_123 : _GEN_2854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2856 = 8'h7c == local_offset_4 ? phv_data_124 : _GEN_2855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2857 = 8'h7d == local_offset_4 ? phv_data_125 : _GEN_2856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2858 = 8'h7e == local_offset_4 ? phv_data_126 : _GEN_2857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2859 = 8'h7f == local_offset_4 ? phv_data_127 : _GEN_2858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2860 = 8'h80 == local_offset_4 ? phv_data_128 : _GEN_2859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2861 = 8'h81 == local_offset_4 ? phv_data_129 : _GEN_2860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2862 = 8'h82 == local_offset_4 ? phv_data_130 : _GEN_2861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2863 = 8'h83 == local_offset_4 ? phv_data_131 : _GEN_2862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2864 = 8'h84 == local_offset_4 ? phv_data_132 : _GEN_2863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2865 = 8'h85 == local_offset_4 ? phv_data_133 : _GEN_2864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2866 = 8'h86 == local_offset_4 ? phv_data_134 : _GEN_2865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2867 = 8'h87 == local_offset_4 ? phv_data_135 : _GEN_2866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2868 = 8'h88 == local_offset_4 ? phv_data_136 : _GEN_2867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2869 = 8'h89 == local_offset_4 ? phv_data_137 : _GEN_2868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2870 = 8'h8a == local_offset_4 ? phv_data_138 : _GEN_2869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2871 = 8'h8b == local_offset_4 ? phv_data_139 : _GEN_2870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2872 = 8'h8c == local_offset_4 ? phv_data_140 : _GEN_2871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2873 = 8'h8d == local_offset_4 ? phv_data_141 : _GEN_2872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2874 = 8'h8e == local_offset_4 ? phv_data_142 : _GEN_2873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2875 = 8'h8f == local_offset_4 ? phv_data_143 : _GEN_2874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2876 = 8'h90 == local_offset_4 ? phv_data_144 : _GEN_2875; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2877 = 8'h91 == local_offset_4 ? phv_data_145 : _GEN_2876; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2878 = 8'h92 == local_offset_4 ? phv_data_146 : _GEN_2877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2879 = 8'h93 == local_offset_4 ? phv_data_147 : _GEN_2878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2880 = 8'h94 == local_offset_4 ? phv_data_148 : _GEN_2879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2881 = 8'h95 == local_offset_4 ? phv_data_149 : _GEN_2880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2882 = 8'h96 == local_offset_4 ? phv_data_150 : _GEN_2881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2883 = 8'h97 == local_offset_4 ? phv_data_151 : _GEN_2882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2884 = 8'h98 == local_offset_4 ? phv_data_152 : _GEN_2883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2885 = 8'h99 == local_offset_4 ? phv_data_153 : _GEN_2884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2886 = 8'h9a == local_offset_4 ? phv_data_154 : _GEN_2885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2887 = 8'h9b == local_offset_4 ? phv_data_155 : _GEN_2886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2888 = 8'h9c == local_offset_4 ? phv_data_156 : _GEN_2887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2889 = 8'h9d == local_offset_4 ? phv_data_157 : _GEN_2888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2890 = 8'h9e == local_offset_4 ? phv_data_158 : _GEN_2889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2891 = 8'h9f == local_offset_4 ? phv_data_159 : _GEN_2890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2893 = 8'h1 == _match_key_qbytes_4_T ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2894 = 8'h2 == _match_key_qbytes_4_T ? phv_data_2 : _GEN_2893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2895 = 8'h3 == _match_key_qbytes_4_T ? phv_data_3 : _GEN_2894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2896 = 8'h4 == _match_key_qbytes_4_T ? phv_data_4 : _GEN_2895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2897 = 8'h5 == _match_key_qbytes_4_T ? phv_data_5 : _GEN_2896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2898 = 8'h6 == _match_key_qbytes_4_T ? phv_data_6 : _GEN_2897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2899 = 8'h7 == _match_key_qbytes_4_T ? phv_data_7 : _GEN_2898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2900 = 8'h8 == _match_key_qbytes_4_T ? phv_data_8 : _GEN_2899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2901 = 8'h9 == _match_key_qbytes_4_T ? phv_data_9 : _GEN_2900; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2902 = 8'ha == _match_key_qbytes_4_T ? phv_data_10 : _GEN_2901; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2903 = 8'hb == _match_key_qbytes_4_T ? phv_data_11 : _GEN_2902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2904 = 8'hc == _match_key_qbytes_4_T ? phv_data_12 : _GEN_2903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2905 = 8'hd == _match_key_qbytes_4_T ? phv_data_13 : _GEN_2904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2906 = 8'he == _match_key_qbytes_4_T ? phv_data_14 : _GEN_2905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2907 = 8'hf == _match_key_qbytes_4_T ? phv_data_15 : _GEN_2906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2908 = 8'h10 == _match_key_qbytes_4_T ? phv_data_16 : _GEN_2907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2909 = 8'h11 == _match_key_qbytes_4_T ? phv_data_17 : _GEN_2908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2910 = 8'h12 == _match_key_qbytes_4_T ? phv_data_18 : _GEN_2909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2911 = 8'h13 == _match_key_qbytes_4_T ? phv_data_19 : _GEN_2910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2912 = 8'h14 == _match_key_qbytes_4_T ? phv_data_20 : _GEN_2911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2913 = 8'h15 == _match_key_qbytes_4_T ? phv_data_21 : _GEN_2912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2914 = 8'h16 == _match_key_qbytes_4_T ? phv_data_22 : _GEN_2913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2915 = 8'h17 == _match_key_qbytes_4_T ? phv_data_23 : _GEN_2914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2916 = 8'h18 == _match_key_qbytes_4_T ? phv_data_24 : _GEN_2915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2917 = 8'h19 == _match_key_qbytes_4_T ? phv_data_25 : _GEN_2916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2918 = 8'h1a == _match_key_qbytes_4_T ? phv_data_26 : _GEN_2917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2919 = 8'h1b == _match_key_qbytes_4_T ? phv_data_27 : _GEN_2918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2920 = 8'h1c == _match_key_qbytes_4_T ? phv_data_28 : _GEN_2919; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2921 = 8'h1d == _match_key_qbytes_4_T ? phv_data_29 : _GEN_2920; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2922 = 8'h1e == _match_key_qbytes_4_T ? phv_data_30 : _GEN_2921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2923 = 8'h1f == _match_key_qbytes_4_T ? phv_data_31 : _GEN_2922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2924 = 8'h20 == _match_key_qbytes_4_T ? phv_data_32 : _GEN_2923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2925 = 8'h21 == _match_key_qbytes_4_T ? phv_data_33 : _GEN_2924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2926 = 8'h22 == _match_key_qbytes_4_T ? phv_data_34 : _GEN_2925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2927 = 8'h23 == _match_key_qbytes_4_T ? phv_data_35 : _GEN_2926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2928 = 8'h24 == _match_key_qbytes_4_T ? phv_data_36 : _GEN_2927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2929 = 8'h25 == _match_key_qbytes_4_T ? phv_data_37 : _GEN_2928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2930 = 8'h26 == _match_key_qbytes_4_T ? phv_data_38 : _GEN_2929; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2931 = 8'h27 == _match_key_qbytes_4_T ? phv_data_39 : _GEN_2930; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2932 = 8'h28 == _match_key_qbytes_4_T ? phv_data_40 : _GEN_2931; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2933 = 8'h29 == _match_key_qbytes_4_T ? phv_data_41 : _GEN_2932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2934 = 8'h2a == _match_key_qbytes_4_T ? phv_data_42 : _GEN_2933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2935 = 8'h2b == _match_key_qbytes_4_T ? phv_data_43 : _GEN_2934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2936 = 8'h2c == _match_key_qbytes_4_T ? phv_data_44 : _GEN_2935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2937 = 8'h2d == _match_key_qbytes_4_T ? phv_data_45 : _GEN_2936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2938 = 8'h2e == _match_key_qbytes_4_T ? phv_data_46 : _GEN_2937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2939 = 8'h2f == _match_key_qbytes_4_T ? phv_data_47 : _GEN_2938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2940 = 8'h30 == _match_key_qbytes_4_T ? phv_data_48 : _GEN_2939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2941 = 8'h31 == _match_key_qbytes_4_T ? phv_data_49 : _GEN_2940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2942 = 8'h32 == _match_key_qbytes_4_T ? phv_data_50 : _GEN_2941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2943 = 8'h33 == _match_key_qbytes_4_T ? phv_data_51 : _GEN_2942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2944 = 8'h34 == _match_key_qbytes_4_T ? phv_data_52 : _GEN_2943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2945 = 8'h35 == _match_key_qbytes_4_T ? phv_data_53 : _GEN_2944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2946 = 8'h36 == _match_key_qbytes_4_T ? phv_data_54 : _GEN_2945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2947 = 8'h37 == _match_key_qbytes_4_T ? phv_data_55 : _GEN_2946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2948 = 8'h38 == _match_key_qbytes_4_T ? phv_data_56 : _GEN_2947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2949 = 8'h39 == _match_key_qbytes_4_T ? phv_data_57 : _GEN_2948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2950 = 8'h3a == _match_key_qbytes_4_T ? phv_data_58 : _GEN_2949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2951 = 8'h3b == _match_key_qbytes_4_T ? phv_data_59 : _GEN_2950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2952 = 8'h3c == _match_key_qbytes_4_T ? phv_data_60 : _GEN_2951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2953 = 8'h3d == _match_key_qbytes_4_T ? phv_data_61 : _GEN_2952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2954 = 8'h3e == _match_key_qbytes_4_T ? phv_data_62 : _GEN_2953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2955 = 8'h3f == _match_key_qbytes_4_T ? phv_data_63 : _GEN_2954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2956 = 8'h40 == _match_key_qbytes_4_T ? phv_data_64 : _GEN_2955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2957 = 8'h41 == _match_key_qbytes_4_T ? phv_data_65 : _GEN_2956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2958 = 8'h42 == _match_key_qbytes_4_T ? phv_data_66 : _GEN_2957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2959 = 8'h43 == _match_key_qbytes_4_T ? phv_data_67 : _GEN_2958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2960 = 8'h44 == _match_key_qbytes_4_T ? phv_data_68 : _GEN_2959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2961 = 8'h45 == _match_key_qbytes_4_T ? phv_data_69 : _GEN_2960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2962 = 8'h46 == _match_key_qbytes_4_T ? phv_data_70 : _GEN_2961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2963 = 8'h47 == _match_key_qbytes_4_T ? phv_data_71 : _GEN_2962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2964 = 8'h48 == _match_key_qbytes_4_T ? phv_data_72 : _GEN_2963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2965 = 8'h49 == _match_key_qbytes_4_T ? phv_data_73 : _GEN_2964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2966 = 8'h4a == _match_key_qbytes_4_T ? phv_data_74 : _GEN_2965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2967 = 8'h4b == _match_key_qbytes_4_T ? phv_data_75 : _GEN_2966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2968 = 8'h4c == _match_key_qbytes_4_T ? phv_data_76 : _GEN_2967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2969 = 8'h4d == _match_key_qbytes_4_T ? phv_data_77 : _GEN_2968; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2970 = 8'h4e == _match_key_qbytes_4_T ? phv_data_78 : _GEN_2969; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2971 = 8'h4f == _match_key_qbytes_4_T ? phv_data_79 : _GEN_2970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2972 = 8'h50 == _match_key_qbytes_4_T ? phv_data_80 : _GEN_2971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2973 = 8'h51 == _match_key_qbytes_4_T ? phv_data_81 : _GEN_2972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2974 = 8'h52 == _match_key_qbytes_4_T ? phv_data_82 : _GEN_2973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2975 = 8'h53 == _match_key_qbytes_4_T ? phv_data_83 : _GEN_2974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2976 = 8'h54 == _match_key_qbytes_4_T ? phv_data_84 : _GEN_2975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2977 = 8'h55 == _match_key_qbytes_4_T ? phv_data_85 : _GEN_2976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2978 = 8'h56 == _match_key_qbytes_4_T ? phv_data_86 : _GEN_2977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2979 = 8'h57 == _match_key_qbytes_4_T ? phv_data_87 : _GEN_2978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2980 = 8'h58 == _match_key_qbytes_4_T ? phv_data_88 : _GEN_2979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2981 = 8'h59 == _match_key_qbytes_4_T ? phv_data_89 : _GEN_2980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2982 = 8'h5a == _match_key_qbytes_4_T ? phv_data_90 : _GEN_2981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2983 = 8'h5b == _match_key_qbytes_4_T ? phv_data_91 : _GEN_2982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2984 = 8'h5c == _match_key_qbytes_4_T ? phv_data_92 : _GEN_2983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2985 = 8'h5d == _match_key_qbytes_4_T ? phv_data_93 : _GEN_2984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2986 = 8'h5e == _match_key_qbytes_4_T ? phv_data_94 : _GEN_2985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2987 = 8'h5f == _match_key_qbytes_4_T ? phv_data_95 : _GEN_2986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2988 = 8'h60 == _match_key_qbytes_4_T ? phv_data_96 : _GEN_2987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2989 = 8'h61 == _match_key_qbytes_4_T ? phv_data_97 : _GEN_2988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2990 = 8'h62 == _match_key_qbytes_4_T ? phv_data_98 : _GEN_2989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2991 = 8'h63 == _match_key_qbytes_4_T ? phv_data_99 : _GEN_2990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2992 = 8'h64 == _match_key_qbytes_4_T ? phv_data_100 : _GEN_2991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2993 = 8'h65 == _match_key_qbytes_4_T ? phv_data_101 : _GEN_2992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2994 = 8'h66 == _match_key_qbytes_4_T ? phv_data_102 : _GEN_2993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2995 = 8'h67 == _match_key_qbytes_4_T ? phv_data_103 : _GEN_2994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2996 = 8'h68 == _match_key_qbytes_4_T ? phv_data_104 : _GEN_2995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2997 = 8'h69 == _match_key_qbytes_4_T ? phv_data_105 : _GEN_2996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2998 = 8'h6a == _match_key_qbytes_4_T ? phv_data_106 : _GEN_2997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2999 = 8'h6b == _match_key_qbytes_4_T ? phv_data_107 : _GEN_2998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3000 = 8'h6c == _match_key_qbytes_4_T ? phv_data_108 : _GEN_2999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3001 = 8'h6d == _match_key_qbytes_4_T ? phv_data_109 : _GEN_3000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3002 = 8'h6e == _match_key_qbytes_4_T ? phv_data_110 : _GEN_3001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3003 = 8'h6f == _match_key_qbytes_4_T ? phv_data_111 : _GEN_3002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3004 = 8'h70 == _match_key_qbytes_4_T ? phv_data_112 : _GEN_3003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3005 = 8'h71 == _match_key_qbytes_4_T ? phv_data_113 : _GEN_3004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3006 = 8'h72 == _match_key_qbytes_4_T ? phv_data_114 : _GEN_3005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3007 = 8'h73 == _match_key_qbytes_4_T ? phv_data_115 : _GEN_3006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3008 = 8'h74 == _match_key_qbytes_4_T ? phv_data_116 : _GEN_3007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3009 = 8'h75 == _match_key_qbytes_4_T ? phv_data_117 : _GEN_3008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3010 = 8'h76 == _match_key_qbytes_4_T ? phv_data_118 : _GEN_3009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3011 = 8'h77 == _match_key_qbytes_4_T ? phv_data_119 : _GEN_3010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3012 = 8'h78 == _match_key_qbytes_4_T ? phv_data_120 : _GEN_3011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3013 = 8'h79 == _match_key_qbytes_4_T ? phv_data_121 : _GEN_3012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3014 = 8'h7a == _match_key_qbytes_4_T ? phv_data_122 : _GEN_3013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3015 = 8'h7b == _match_key_qbytes_4_T ? phv_data_123 : _GEN_3014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3016 = 8'h7c == _match_key_qbytes_4_T ? phv_data_124 : _GEN_3015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3017 = 8'h7d == _match_key_qbytes_4_T ? phv_data_125 : _GEN_3016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3018 = 8'h7e == _match_key_qbytes_4_T ? phv_data_126 : _GEN_3017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3019 = 8'h7f == _match_key_qbytes_4_T ? phv_data_127 : _GEN_3018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3020 = 8'h80 == _match_key_qbytes_4_T ? phv_data_128 : _GEN_3019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3021 = 8'h81 == _match_key_qbytes_4_T ? phv_data_129 : _GEN_3020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3022 = 8'h82 == _match_key_qbytes_4_T ? phv_data_130 : _GEN_3021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3023 = 8'h83 == _match_key_qbytes_4_T ? phv_data_131 : _GEN_3022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3024 = 8'h84 == _match_key_qbytes_4_T ? phv_data_132 : _GEN_3023; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3025 = 8'h85 == _match_key_qbytes_4_T ? phv_data_133 : _GEN_3024; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3026 = 8'h86 == _match_key_qbytes_4_T ? phv_data_134 : _GEN_3025; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3027 = 8'h87 == _match_key_qbytes_4_T ? phv_data_135 : _GEN_3026; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3028 = 8'h88 == _match_key_qbytes_4_T ? phv_data_136 : _GEN_3027; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3029 = 8'h89 == _match_key_qbytes_4_T ? phv_data_137 : _GEN_3028; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3030 = 8'h8a == _match_key_qbytes_4_T ? phv_data_138 : _GEN_3029; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3031 = 8'h8b == _match_key_qbytes_4_T ? phv_data_139 : _GEN_3030; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3032 = 8'h8c == _match_key_qbytes_4_T ? phv_data_140 : _GEN_3031; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3033 = 8'h8d == _match_key_qbytes_4_T ? phv_data_141 : _GEN_3032; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3034 = 8'h8e == _match_key_qbytes_4_T ? phv_data_142 : _GEN_3033; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3035 = 8'h8f == _match_key_qbytes_4_T ? phv_data_143 : _GEN_3034; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3036 = 8'h90 == _match_key_qbytes_4_T ? phv_data_144 : _GEN_3035; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3037 = 8'h91 == _match_key_qbytes_4_T ? phv_data_145 : _GEN_3036; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3038 = 8'h92 == _match_key_qbytes_4_T ? phv_data_146 : _GEN_3037; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3039 = 8'h93 == _match_key_qbytes_4_T ? phv_data_147 : _GEN_3038; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3040 = 8'h94 == _match_key_qbytes_4_T ? phv_data_148 : _GEN_3039; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3041 = 8'h95 == _match_key_qbytes_4_T ? phv_data_149 : _GEN_3040; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3042 = 8'h96 == _match_key_qbytes_4_T ? phv_data_150 : _GEN_3041; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3043 = 8'h97 == _match_key_qbytes_4_T ? phv_data_151 : _GEN_3042; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3044 = 8'h98 == _match_key_qbytes_4_T ? phv_data_152 : _GEN_3043; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3045 = 8'h99 == _match_key_qbytes_4_T ? phv_data_153 : _GEN_3044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3046 = 8'h9a == _match_key_qbytes_4_T ? phv_data_154 : _GEN_3045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3047 = 8'h9b == _match_key_qbytes_4_T ? phv_data_155 : _GEN_3046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3048 = 8'h9c == _match_key_qbytes_4_T ? phv_data_156 : _GEN_3047; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3049 = 8'h9d == _match_key_qbytes_4_T ? phv_data_157 : _GEN_3048; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3050 = 8'h9e == _match_key_qbytes_4_T ? phv_data_158 : _GEN_3049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3051 = 8'h9f == _match_key_qbytes_4_T ? phv_data_159 : _GEN_3050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3053 = 8'h1 == _match_key_qbytes_4_T_1 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3054 = 8'h2 == _match_key_qbytes_4_T_1 ? phv_data_2 : _GEN_3053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3055 = 8'h3 == _match_key_qbytes_4_T_1 ? phv_data_3 : _GEN_3054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3056 = 8'h4 == _match_key_qbytes_4_T_1 ? phv_data_4 : _GEN_3055; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3057 = 8'h5 == _match_key_qbytes_4_T_1 ? phv_data_5 : _GEN_3056; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3058 = 8'h6 == _match_key_qbytes_4_T_1 ? phv_data_6 : _GEN_3057; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3059 = 8'h7 == _match_key_qbytes_4_T_1 ? phv_data_7 : _GEN_3058; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3060 = 8'h8 == _match_key_qbytes_4_T_1 ? phv_data_8 : _GEN_3059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3061 = 8'h9 == _match_key_qbytes_4_T_1 ? phv_data_9 : _GEN_3060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3062 = 8'ha == _match_key_qbytes_4_T_1 ? phv_data_10 : _GEN_3061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3063 = 8'hb == _match_key_qbytes_4_T_1 ? phv_data_11 : _GEN_3062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3064 = 8'hc == _match_key_qbytes_4_T_1 ? phv_data_12 : _GEN_3063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3065 = 8'hd == _match_key_qbytes_4_T_1 ? phv_data_13 : _GEN_3064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3066 = 8'he == _match_key_qbytes_4_T_1 ? phv_data_14 : _GEN_3065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3067 = 8'hf == _match_key_qbytes_4_T_1 ? phv_data_15 : _GEN_3066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3068 = 8'h10 == _match_key_qbytes_4_T_1 ? phv_data_16 : _GEN_3067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3069 = 8'h11 == _match_key_qbytes_4_T_1 ? phv_data_17 : _GEN_3068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3070 = 8'h12 == _match_key_qbytes_4_T_1 ? phv_data_18 : _GEN_3069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3071 = 8'h13 == _match_key_qbytes_4_T_1 ? phv_data_19 : _GEN_3070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3072 = 8'h14 == _match_key_qbytes_4_T_1 ? phv_data_20 : _GEN_3071; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3073 = 8'h15 == _match_key_qbytes_4_T_1 ? phv_data_21 : _GEN_3072; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3074 = 8'h16 == _match_key_qbytes_4_T_1 ? phv_data_22 : _GEN_3073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3075 = 8'h17 == _match_key_qbytes_4_T_1 ? phv_data_23 : _GEN_3074; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3076 = 8'h18 == _match_key_qbytes_4_T_1 ? phv_data_24 : _GEN_3075; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3077 = 8'h19 == _match_key_qbytes_4_T_1 ? phv_data_25 : _GEN_3076; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3078 = 8'h1a == _match_key_qbytes_4_T_1 ? phv_data_26 : _GEN_3077; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3079 = 8'h1b == _match_key_qbytes_4_T_1 ? phv_data_27 : _GEN_3078; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3080 = 8'h1c == _match_key_qbytes_4_T_1 ? phv_data_28 : _GEN_3079; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3081 = 8'h1d == _match_key_qbytes_4_T_1 ? phv_data_29 : _GEN_3080; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3082 = 8'h1e == _match_key_qbytes_4_T_1 ? phv_data_30 : _GEN_3081; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3083 = 8'h1f == _match_key_qbytes_4_T_1 ? phv_data_31 : _GEN_3082; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3084 = 8'h20 == _match_key_qbytes_4_T_1 ? phv_data_32 : _GEN_3083; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3085 = 8'h21 == _match_key_qbytes_4_T_1 ? phv_data_33 : _GEN_3084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3086 = 8'h22 == _match_key_qbytes_4_T_1 ? phv_data_34 : _GEN_3085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3087 = 8'h23 == _match_key_qbytes_4_T_1 ? phv_data_35 : _GEN_3086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3088 = 8'h24 == _match_key_qbytes_4_T_1 ? phv_data_36 : _GEN_3087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3089 = 8'h25 == _match_key_qbytes_4_T_1 ? phv_data_37 : _GEN_3088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3090 = 8'h26 == _match_key_qbytes_4_T_1 ? phv_data_38 : _GEN_3089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3091 = 8'h27 == _match_key_qbytes_4_T_1 ? phv_data_39 : _GEN_3090; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3092 = 8'h28 == _match_key_qbytes_4_T_1 ? phv_data_40 : _GEN_3091; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3093 = 8'h29 == _match_key_qbytes_4_T_1 ? phv_data_41 : _GEN_3092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3094 = 8'h2a == _match_key_qbytes_4_T_1 ? phv_data_42 : _GEN_3093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3095 = 8'h2b == _match_key_qbytes_4_T_1 ? phv_data_43 : _GEN_3094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3096 = 8'h2c == _match_key_qbytes_4_T_1 ? phv_data_44 : _GEN_3095; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3097 = 8'h2d == _match_key_qbytes_4_T_1 ? phv_data_45 : _GEN_3096; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3098 = 8'h2e == _match_key_qbytes_4_T_1 ? phv_data_46 : _GEN_3097; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3099 = 8'h2f == _match_key_qbytes_4_T_1 ? phv_data_47 : _GEN_3098; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3100 = 8'h30 == _match_key_qbytes_4_T_1 ? phv_data_48 : _GEN_3099; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3101 = 8'h31 == _match_key_qbytes_4_T_1 ? phv_data_49 : _GEN_3100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3102 = 8'h32 == _match_key_qbytes_4_T_1 ? phv_data_50 : _GEN_3101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3103 = 8'h33 == _match_key_qbytes_4_T_1 ? phv_data_51 : _GEN_3102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3104 = 8'h34 == _match_key_qbytes_4_T_1 ? phv_data_52 : _GEN_3103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3105 = 8'h35 == _match_key_qbytes_4_T_1 ? phv_data_53 : _GEN_3104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3106 = 8'h36 == _match_key_qbytes_4_T_1 ? phv_data_54 : _GEN_3105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3107 = 8'h37 == _match_key_qbytes_4_T_1 ? phv_data_55 : _GEN_3106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3108 = 8'h38 == _match_key_qbytes_4_T_1 ? phv_data_56 : _GEN_3107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3109 = 8'h39 == _match_key_qbytes_4_T_1 ? phv_data_57 : _GEN_3108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3110 = 8'h3a == _match_key_qbytes_4_T_1 ? phv_data_58 : _GEN_3109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3111 = 8'h3b == _match_key_qbytes_4_T_1 ? phv_data_59 : _GEN_3110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3112 = 8'h3c == _match_key_qbytes_4_T_1 ? phv_data_60 : _GEN_3111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3113 = 8'h3d == _match_key_qbytes_4_T_1 ? phv_data_61 : _GEN_3112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3114 = 8'h3e == _match_key_qbytes_4_T_1 ? phv_data_62 : _GEN_3113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3115 = 8'h3f == _match_key_qbytes_4_T_1 ? phv_data_63 : _GEN_3114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3116 = 8'h40 == _match_key_qbytes_4_T_1 ? phv_data_64 : _GEN_3115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3117 = 8'h41 == _match_key_qbytes_4_T_1 ? phv_data_65 : _GEN_3116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3118 = 8'h42 == _match_key_qbytes_4_T_1 ? phv_data_66 : _GEN_3117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3119 = 8'h43 == _match_key_qbytes_4_T_1 ? phv_data_67 : _GEN_3118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3120 = 8'h44 == _match_key_qbytes_4_T_1 ? phv_data_68 : _GEN_3119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3121 = 8'h45 == _match_key_qbytes_4_T_1 ? phv_data_69 : _GEN_3120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3122 = 8'h46 == _match_key_qbytes_4_T_1 ? phv_data_70 : _GEN_3121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3123 = 8'h47 == _match_key_qbytes_4_T_1 ? phv_data_71 : _GEN_3122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3124 = 8'h48 == _match_key_qbytes_4_T_1 ? phv_data_72 : _GEN_3123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3125 = 8'h49 == _match_key_qbytes_4_T_1 ? phv_data_73 : _GEN_3124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3126 = 8'h4a == _match_key_qbytes_4_T_1 ? phv_data_74 : _GEN_3125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3127 = 8'h4b == _match_key_qbytes_4_T_1 ? phv_data_75 : _GEN_3126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3128 = 8'h4c == _match_key_qbytes_4_T_1 ? phv_data_76 : _GEN_3127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3129 = 8'h4d == _match_key_qbytes_4_T_1 ? phv_data_77 : _GEN_3128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3130 = 8'h4e == _match_key_qbytes_4_T_1 ? phv_data_78 : _GEN_3129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3131 = 8'h4f == _match_key_qbytes_4_T_1 ? phv_data_79 : _GEN_3130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3132 = 8'h50 == _match_key_qbytes_4_T_1 ? phv_data_80 : _GEN_3131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3133 = 8'h51 == _match_key_qbytes_4_T_1 ? phv_data_81 : _GEN_3132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3134 = 8'h52 == _match_key_qbytes_4_T_1 ? phv_data_82 : _GEN_3133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3135 = 8'h53 == _match_key_qbytes_4_T_1 ? phv_data_83 : _GEN_3134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3136 = 8'h54 == _match_key_qbytes_4_T_1 ? phv_data_84 : _GEN_3135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3137 = 8'h55 == _match_key_qbytes_4_T_1 ? phv_data_85 : _GEN_3136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3138 = 8'h56 == _match_key_qbytes_4_T_1 ? phv_data_86 : _GEN_3137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3139 = 8'h57 == _match_key_qbytes_4_T_1 ? phv_data_87 : _GEN_3138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3140 = 8'h58 == _match_key_qbytes_4_T_1 ? phv_data_88 : _GEN_3139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3141 = 8'h59 == _match_key_qbytes_4_T_1 ? phv_data_89 : _GEN_3140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3142 = 8'h5a == _match_key_qbytes_4_T_1 ? phv_data_90 : _GEN_3141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3143 = 8'h5b == _match_key_qbytes_4_T_1 ? phv_data_91 : _GEN_3142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3144 = 8'h5c == _match_key_qbytes_4_T_1 ? phv_data_92 : _GEN_3143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3145 = 8'h5d == _match_key_qbytes_4_T_1 ? phv_data_93 : _GEN_3144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3146 = 8'h5e == _match_key_qbytes_4_T_1 ? phv_data_94 : _GEN_3145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3147 = 8'h5f == _match_key_qbytes_4_T_1 ? phv_data_95 : _GEN_3146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3148 = 8'h60 == _match_key_qbytes_4_T_1 ? phv_data_96 : _GEN_3147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3149 = 8'h61 == _match_key_qbytes_4_T_1 ? phv_data_97 : _GEN_3148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3150 = 8'h62 == _match_key_qbytes_4_T_1 ? phv_data_98 : _GEN_3149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3151 = 8'h63 == _match_key_qbytes_4_T_1 ? phv_data_99 : _GEN_3150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3152 = 8'h64 == _match_key_qbytes_4_T_1 ? phv_data_100 : _GEN_3151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3153 = 8'h65 == _match_key_qbytes_4_T_1 ? phv_data_101 : _GEN_3152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3154 = 8'h66 == _match_key_qbytes_4_T_1 ? phv_data_102 : _GEN_3153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3155 = 8'h67 == _match_key_qbytes_4_T_1 ? phv_data_103 : _GEN_3154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3156 = 8'h68 == _match_key_qbytes_4_T_1 ? phv_data_104 : _GEN_3155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3157 = 8'h69 == _match_key_qbytes_4_T_1 ? phv_data_105 : _GEN_3156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3158 = 8'h6a == _match_key_qbytes_4_T_1 ? phv_data_106 : _GEN_3157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3159 = 8'h6b == _match_key_qbytes_4_T_1 ? phv_data_107 : _GEN_3158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3160 = 8'h6c == _match_key_qbytes_4_T_1 ? phv_data_108 : _GEN_3159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3161 = 8'h6d == _match_key_qbytes_4_T_1 ? phv_data_109 : _GEN_3160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3162 = 8'h6e == _match_key_qbytes_4_T_1 ? phv_data_110 : _GEN_3161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3163 = 8'h6f == _match_key_qbytes_4_T_1 ? phv_data_111 : _GEN_3162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3164 = 8'h70 == _match_key_qbytes_4_T_1 ? phv_data_112 : _GEN_3163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3165 = 8'h71 == _match_key_qbytes_4_T_1 ? phv_data_113 : _GEN_3164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3166 = 8'h72 == _match_key_qbytes_4_T_1 ? phv_data_114 : _GEN_3165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3167 = 8'h73 == _match_key_qbytes_4_T_1 ? phv_data_115 : _GEN_3166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3168 = 8'h74 == _match_key_qbytes_4_T_1 ? phv_data_116 : _GEN_3167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3169 = 8'h75 == _match_key_qbytes_4_T_1 ? phv_data_117 : _GEN_3168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3170 = 8'h76 == _match_key_qbytes_4_T_1 ? phv_data_118 : _GEN_3169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3171 = 8'h77 == _match_key_qbytes_4_T_1 ? phv_data_119 : _GEN_3170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3172 = 8'h78 == _match_key_qbytes_4_T_1 ? phv_data_120 : _GEN_3171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3173 = 8'h79 == _match_key_qbytes_4_T_1 ? phv_data_121 : _GEN_3172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3174 = 8'h7a == _match_key_qbytes_4_T_1 ? phv_data_122 : _GEN_3173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3175 = 8'h7b == _match_key_qbytes_4_T_1 ? phv_data_123 : _GEN_3174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3176 = 8'h7c == _match_key_qbytes_4_T_1 ? phv_data_124 : _GEN_3175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3177 = 8'h7d == _match_key_qbytes_4_T_1 ? phv_data_125 : _GEN_3176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3178 = 8'h7e == _match_key_qbytes_4_T_1 ? phv_data_126 : _GEN_3177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3179 = 8'h7f == _match_key_qbytes_4_T_1 ? phv_data_127 : _GEN_3178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3180 = 8'h80 == _match_key_qbytes_4_T_1 ? phv_data_128 : _GEN_3179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3181 = 8'h81 == _match_key_qbytes_4_T_1 ? phv_data_129 : _GEN_3180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3182 = 8'h82 == _match_key_qbytes_4_T_1 ? phv_data_130 : _GEN_3181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3183 = 8'h83 == _match_key_qbytes_4_T_1 ? phv_data_131 : _GEN_3182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3184 = 8'h84 == _match_key_qbytes_4_T_1 ? phv_data_132 : _GEN_3183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3185 = 8'h85 == _match_key_qbytes_4_T_1 ? phv_data_133 : _GEN_3184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3186 = 8'h86 == _match_key_qbytes_4_T_1 ? phv_data_134 : _GEN_3185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3187 = 8'h87 == _match_key_qbytes_4_T_1 ? phv_data_135 : _GEN_3186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3188 = 8'h88 == _match_key_qbytes_4_T_1 ? phv_data_136 : _GEN_3187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3189 = 8'h89 == _match_key_qbytes_4_T_1 ? phv_data_137 : _GEN_3188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3190 = 8'h8a == _match_key_qbytes_4_T_1 ? phv_data_138 : _GEN_3189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3191 = 8'h8b == _match_key_qbytes_4_T_1 ? phv_data_139 : _GEN_3190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3192 = 8'h8c == _match_key_qbytes_4_T_1 ? phv_data_140 : _GEN_3191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3193 = 8'h8d == _match_key_qbytes_4_T_1 ? phv_data_141 : _GEN_3192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3194 = 8'h8e == _match_key_qbytes_4_T_1 ? phv_data_142 : _GEN_3193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3195 = 8'h8f == _match_key_qbytes_4_T_1 ? phv_data_143 : _GEN_3194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3196 = 8'h90 == _match_key_qbytes_4_T_1 ? phv_data_144 : _GEN_3195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3197 = 8'h91 == _match_key_qbytes_4_T_1 ? phv_data_145 : _GEN_3196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3198 = 8'h92 == _match_key_qbytes_4_T_1 ? phv_data_146 : _GEN_3197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3199 = 8'h93 == _match_key_qbytes_4_T_1 ? phv_data_147 : _GEN_3198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3200 = 8'h94 == _match_key_qbytes_4_T_1 ? phv_data_148 : _GEN_3199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3201 = 8'h95 == _match_key_qbytes_4_T_1 ? phv_data_149 : _GEN_3200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3202 = 8'h96 == _match_key_qbytes_4_T_1 ? phv_data_150 : _GEN_3201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3203 = 8'h97 == _match_key_qbytes_4_T_1 ? phv_data_151 : _GEN_3202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3204 = 8'h98 == _match_key_qbytes_4_T_1 ? phv_data_152 : _GEN_3203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3205 = 8'h99 == _match_key_qbytes_4_T_1 ? phv_data_153 : _GEN_3204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3206 = 8'h9a == _match_key_qbytes_4_T_1 ? phv_data_154 : _GEN_3205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3207 = 8'h9b == _match_key_qbytes_4_T_1 ? phv_data_155 : _GEN_3206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3208 = 8'h9c == _match_key_qbytes_4_T_1 ? phv_data_156 : _GEN_3207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3209 = 8'h9d == _match_key_qbytes_4_T_1 ? phv_data_157 : _GEN_3208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3210 = 8'h9e == _match_key_qbytes_4_T_1 ? phv_data_158 : _GEN_3209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3211 = 8'h9f == _match_key_qbytes_4_T_1 ? phv_data_159 : _GEN_3210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [31:0] _match_key_qbytes_4_T_3 = {_GEN_3051,_GEN_3211,_GEN_2731,_GEN_2891}; // @[Cat.scala 30:58]
  wire [31:0] match_key_qbytes_4 = local_offset_4 < end_offset ? _match_key_qbytes_4_T_3 : 32'h0; // @[matcher.scala 88:54 matcher.scala 89:45 matcher.scala 97:45]
  wire [7:0] local_offset_5 = 8'h14 + read_key_offset; // @[matcher.scala 87:77]
  wire [5:0] match_key_qbytes_5_hi = local_offset_5[7:2]; // @[matcher.scala 91:54]
  wire [7:0] _match_key_qbytes_5_T = {match_key_qbytes_5_hi,2'h3}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_5_T_1 = {match_key_qbytes_5_hi,2'h2}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_5_T_2 = {match_key_qbytes_5_hi,2'h1}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_3214 = 8'h1 == _match_key_qbytes_5_T_2 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3215 = 8'h2 == _match_key_qbytes_5_T_2 ? phv_data_2 : _GEN_3214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3216 = 8'h3 == _match_key_qbytes_5_T_2 ? phv_data_3 : _GEN_3215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3217 = 8'h4 == _match_key_qbytes_5_T_2 ? phv_data_4 : _GEN_3216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3218 = 8'h5 == _match_key_qbytes_5_T_2 ? phv_data_5 : _GEN_3217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3219 = 8'h6 == _match_key_qbytes_5_T_2 ? phv_data_6 : _GEN_3218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3220 = 8'h7 == _match_key_qbytes_5_T_2 ? phv_data_7 : _GEN_3219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3221 = 8'h8 == _match_key_qbytes_5_T_2 ? phv_data_8 : _GEN_3220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3222 = 8'h9 == _match_key_qbytes_5_T_2 ? phv_data_9 : _GEN_3221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3223 = 8'ha == _match_key_qbytes_5_T_2 ? phv_data_10 : _GEN_3222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3224 = 8'hb == _match_key_qbytes_5_T_2 ? phv_data_11 : _GEN_3223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3225 = 8'hc == _match_key_qbytes_5_T_2 ? phv_data_12 : _GEN_3224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3226 = 8'hd == _match_key_qbytes_5_T_2 ? phv_data_13 : _GEN_3225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3227 = 8'he == _match_key_qbytes_5_T_2 ? phv_data_14 : _GEN_3226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3228 = 8'hf == _match_key_qbytes_5_T_2 ? phv_data_15 : _GEN_3227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3229 = 8'h10 == _match_key_qbytes_5_T_2 ? phv_data_16 : _GEN_3228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3230 = 8'h11 == _match_key_qbytes_5_T_2 ? phv_data_17 : _GEN_3229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3231 = 8'h12 == _match_key_qbytes_5_T_2 ? phv_data_18 : _GEN_3230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3232 = 8'h13 == _match_key_qbytes_5_T_2 ? phv_data_19 : _GEN_3231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3233 = 8'h14 == _match_key_qbytes_5_T_2 ? phv_data_20 : _GEN_3232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3234 = 8'h15 == _match_key_qbytes_5_T_2 ? phv_data_21 : _GEN_3233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3235 = 8'h16 == _match_key_qbytes_5_T_2 ? phv_data_22 : _GEN_3234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3236 = 8'h17 == _match_key_qbytes_5_T_2 ? phv_data_23 : _GEN_3235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3237 = 8'h18 == _match_key_qbytes_5_T_2 ? phv_data_24 : _GEN_3236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3238 = 8'h19 == _match_key_qbytes_5_T_2 ? phv_data_25 : _GEN_3237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3239 = 8'h1a == _match_key_qbytes_5_T_2 ? phv_data_26 : _GEN_3238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3240 = 8'h1b == _match_key_qbytes_5_T_2 ? phv_data_27 : _GEN_3239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3241 = 8'h1c == _match_key_qbytes_5_T_2 ? phv_data_28 : _GEN_3240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3242 = 8'h1d == _match_key_qbytes_5_T_2 ? phv_data_29 : _GEN_3241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3243 = 8'h1e == _match_key_qbytes_5_T_2 ? phv_data_30 : _GEN_3242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3244 = 8'h1f == _match_key_qbytes_5_T_2 ? phv_data_31 : _GEN_3243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3245 = 8'h20 == _match_key_qbytes_5_T_2 ? phv_data_32 : _GEN_3244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3246 = 8'h21 == _match_key_qbytes_5_T_2 ? phv_data_33 : _GEN_3245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3247 = 8'h22 == _match_key_qbytes_5_T_2 ? phv_data_34 : _GEN_3246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3248 = 8'h23 == _match_key_qbytes_5_T_2 ? phv_data_35 : _GEN_3247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3249 = 8'h24 == _match_key_qbytes_5_T_2 ? phv_data_36 : _GEN_3248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3250 = 8'h25 == _match_key_qbytes_5_T_2 ? phv_data_37 : _GEN_3249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3251 = 8'h26 == _match_key_qbytes_5_T_2 ? phv_data_38 : _GEN_3250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3252 = 8'h27 == _match_key_qbytes_5_T_2 ? phv_data_39 : _GEN_3251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3253 = 8'h28 == _match_key_qbytes_5_T_2 ? phv_data_40 : _GEN_3252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3254 = 8'h29 == _match_key_qbytes_5_T_2 ? phv_data_41 : _GEN_3253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3255 = 8'h2a == _match_key_qbytes_5_T_2 ? phv_data_42 : _GEN_3254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3256 = 8'h2b == _match_key_qbytes_5_T_2 ? phv_data_43 : _GEN_3255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3257 = 8'h2c == _match_key_qbytes_5_T_2 ? phv_data_44 : _GEN_3256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3258 = 8'h2d == _match_key_qbytes_5_T_2 ? phv_data_45 : _GEN_3257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3259 = 8'h2e == _match_key_qbytes_5_T_2 ? phv_data_46 : _GEN_3258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3260 = 8'h2f == _match_key_qbytes_5_T_2 ? phv_data_47 : _GEN_3259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3261 = 8'h30 == _match_key_qbytes_5_T_2 ? phv_data_48 : _GEN_3260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3262 = 8'h31 == _match_key_qbytes_5_T_2 ? phv_data_49 : _GEN_3261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3263 = 8'h32 == _match_key_qbytes_5_T_2 ? phv_data_50 : _GEN_3262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3264 = 8'h33 == _match_key_qbytes_5_T_2 ? phv_data_51 : _GEN_3263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3265 = 8'h34 == _match_key_qbytes_5_T_2 ? phv_data_52 : _GEN_3264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3266 = 8'h35 == _match_key_qbytes_5_T_2 ? phv_data_53 : _GEN_3265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3267 = 8'h36 == _match_key_qbytes_5_T_2 ? phv_data_54 : _GEN_3266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3268 = 8'h37 == _match_key_qbytes_5_T_2 ? phv_data_55 : _GEN_3267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3269 = 8'h38 == _match_key_qbytes_5_T_2 ? phv_data_56 : _GEN_3268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3270 = 8'h39 == _match_key_qbytes_5_T_2 ? phv_data_57 : _GEN_3269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3271 = 8'h3a == _match_key_qbytes_5_T_2 ? phv_data_58 : _GEN_3270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3272 = 8'h3b == _match_key_qbytes_5_T_2 ? phv_data_59 : _GEN_3271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3273 = 8'h3c == _match_key_qbytes_5_T_2 ? phv_data_60 : _GEN_3272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3274 = 8'h3d == _match_key_qbytes_5_T_2 ? phv_data_61 : _GEN_3273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3275 = 8'h3e == _match_key_qbytes_5_T_2 ? phv_data_62 : _GEN_3274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3276 = 8'h3f == _match_key_qbytes_5_T_2 ? phv_data_63 : _GEN_3275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3277 = 8'h40 == _match_key_qbytes_5_T_2 ? phv_data_64 : _GEN_3276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3278 = 8'h41 == _match_key_qbytes_5_T_2 ? phv_data_65 : _GEN_3277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3279 = 8'h42 == _match_key_qbytes_5_T_2 ? phv_data_66 : _GEN_3278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3280 = 8'h43 == _match_key_qbytes_5_T_2 ? phv_data_67 : _GEN_3279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3281 = 8'h44 == _match_key_qbytes_5_T_2 ? phv_data_68 : _GEN_3280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3282 = 8'h45 == _match_key_qbytes_5_T_2 ? phv_data_69 : _GEN_3281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3283 = 8'h46 == _match_key_qbytes_5_T_2 ? phv_data_70 : _GEN_3282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3284 = 8'h47 == _match_key_qbytes_5_T_2 ? phv_data_71 : _GEN_3283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3285 = 8'h48 == _match_key_qbytes_5_T_2 ? phv_data_72 : _GEN_3284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3286 = 8'h49 == _match_key_qbytes_5_T_2 ? phv_data_73 : _GEN_3285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3287 = 8'h4a == _match_key_qbytes_5_T_2 ? phv_data_74 : _GEN_3286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3288 = 8'h4b == _match_key_qbytes_5_T_2 ? phv_data_75 : _GEN_3287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3289 = 8'h4c == _match_key_qbytes_5_T_2 ? phv_data_76 : _GEN_3288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3290 = 8'h4d == _match_key_qbytes_5_T_2 ? phv_data_77 : _GEN_3289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3291 = 8'h4e == _match_key_qbytes_5_T_2 ? phv_data_78 : _GEN_3290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3292 = 8'h4f == _match_key_qbytes_5_T_2 ? phv_data_79 : _GEN_3291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3293 = 8'h50 == _match_key_qbytes_5_T_2 ? phv_data_80 : _GEN_3292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3294 = 8'h51 == _match_key_qbytes_5_T_2 ? phv_data_81 : _GEN_3293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3295 = 8'h52 == _match_key_qbytes_5_T_2 ? phv_data_82 : _GEN_3294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3296 = 8'h53 == _match_key_qbytes_5_T_2 ? phv_data_83 : _GEN_3295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3297 = 8'h54 == _match_key_qbytes_5_T_2 ? phv_data_84 : _GEN_3296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3298 = 8'h55 == _match_key_qbytes_5_T_2 ? phv_data_85 : _GEN_3297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3299 = 8'h56 == _match_key_qbytes_5_T_2 ? phv_data_86 : _GEN_3298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3300 = 8'h57 == _match_key_qbytes_5_T_2 ? phv_data_87 : _GEN_3299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3301 = 8'h58 == _match_key_qbytes_5_T_2 ? phv_data_88 : _GEN_3300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3302 = 8'h59 == _match_key_qbytes_5_T_2 ? phv_data_89 : _GEN_3301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3303 = 8'h5a == _match_key_qbytes_5_T_2 ? phv_data_90 : _GEN_3302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3304 = 8'h5b == _match_key_qbytes_5_T_2 ? phv_data_91 : _GEN_3303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3305 = 8'h5c == _match_key_qbytes_5_T_2 ? phv_data_92 : _GEN_3304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3306 = 8'h5d == _match_key_qbytes_5_T_2 ? phv_data_93 : _GEN_3305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3307 = 8'h5e == _match_key_qbytes_5_T_2 ? phv_data_94 : _GEN_3306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3308 = 8'h5f == _match_key_qbytes_5_T_2 ? phv_data_95 : _GEN_3307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3309 = 8'h60 == _match_key_qbytes_5_T_2 ? phv_data_96 : _GEN_3308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3310 = 8'h61 == _match_key_qbytes_5_T_2 ? phv_data_97 : _GEN_3309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3311 = 8'h62 == _match_key_qbytes_5_T_2 ? phv_data_98 : _GEN_3310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3312 = 8'h63 == _match_key_qbytes_5_T_2 ? phv_data_99 : _GEN_3311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3313 = 8'h64 == _match_key_qbytes_5_T_2 ? phv_data_100 : _GEN_3312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3314 = 8'h65 == _match_key_qbytes_5_T_2 ? phv_data_101 : _GEN_3313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3315 = 8'h66 == _match_key_qbytes_5_T_2 ? phv_data_102 : _GEN_3314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3316 = 8'h67 == _match_key_qbytes_5_T_2 ? phv_data_103 : _GEN_3315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3317 = 8'h68 == _match_key_qbytes_5_T_2 ? phv_data_104 : _GEN_3316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3318 = 8'h69 == _match_key_qbytes_5_T_2 ? phv_data_105 : _GEN_3317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3319 = 8'h6a == _match_key_qbytes_5_T_2 ? phv_data_106 : _GEN_3318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3320 = 8'h6b == _match_key_qbytes_5_T_2 ? phv_data_107 : _GEN_3319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3321 = 8'h6c == _match_key_qbytes_5_T_2 ? phv_data_108 : _GEN_3320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3322 = 8'h6d == _match_key_qbytes_5_T_2 ? phv_data_109 : _GEN_3321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3323 = 8'h6e == _match_key_qbytes_5_T_2 ? phv_data_110 : _GEN_3322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3324 = 8'h6f == _match_key_qbytes_5_T_2 ? phv_data_111 : _GEN_3323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3325 = 8'h70 == _match_key_qbytes_5_T_2 ? phv_data_112 : _GEN_3324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3326 = 8'h71 == _match_key_qbytes_5_T_2 ? phv_data_113 : _GEN_3325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3327 = 8'h72 == _match_key_qbytes_5_T_2 ? phv_data_114 : _GEN_3326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3328 = 8'h73 == _match_key_qbytes_5_T_2 ? phv_data_115 : _GEN_3327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3329 = 8'h74 == _match_key_qbytes_5_T_2 ? phv_data_116 : _GEN_3328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3330 = 8'h75 == _match_key_qbytes_5_T_2 ? phv_data_117 : _GEN_3329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3331 = 8'h76 == _match_key_qbytes_5_T_2 ? phv_data_118 : _GEN_3330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3332 = 8'h77 == _match_key_qbytes_5_T_2 ? phv_data_119 : _GEN_3331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3333 = 8'h78 == _match_key_qbytes_5_T_2 ? phv_data_120 : _GEN_3332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3334 = 8'h79 == _match_key_qbytes_5_T_2 ? phv_data_121 : _GEN_3333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3335 = 8'h7a == _match_key_qbytes_5_T_2 ? phv_data_122 : _GEN_3334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3336 = 8'h7b == _match_key_qbytes_5_T_2 ? phv_data_123 : _GEN_3335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3337 = 8'h7c == _match_key_qbytes_5_T_2 ? phv_data_124 : _GEN_3336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3338 = 8'h7d == _match_key_qbytes_5_T_2 ? phv_data_125 : _GEN_3337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3339 = 8'h7e == _match_key_qbytes_5_T_2 ? phv_data_126 : _GEN_3338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3340 = 8'h7f == _match_key_qbytes_5_T_2 ? phv_data_127 : _GEN_3339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3341 = 8'h80 == _match_key_qbytes_5_T_2 ? phv_data_128 : _GEN_3340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3342 = 8'h81 == _match_key_qbytes_5_T_2 ? phv_data_129 : _GEN_3341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3343 = 8'h82 == _match_key_qbytes_5_T_2 ? phv_data_130 : _GEN_3342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3344 = 8'h83 == _match_key_qbytes_5_T_2 ? phv_data_131 : _GEN_3343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3345 = 8'h84 == _match_key_qbytes_5_T_2 ? phv_data_132 : _GEN_3344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3346 = 8'h85 == _match_key_qbytes_5_T_2 ? phv_data_133 : _GEN_3345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3347 = 8'h86 == _match_key_qbytes_5_T_2 ? phv_data_134 : _GEN_3346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3348 = 8'h87 == _match_key_qbytes_5_T_2 ? phv_data_135 : _GEN_3347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3349 = 8'h88 == _match_key_qbytes_5_T_2 ? phv_data_136 : _GEN_3348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3350 = 8'h89 == _match_key_qbytes_5_T_2 ? phv_data_137 : _GEN_3349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3351 = 8'h8a == _match_key_qbytes_5_T_2 ? phv_data_138 : _GEN_3350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3352 = 8'h8b == _match_key_qbytes_5_T_2 ? phv_data_139 : _GEN_3351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3353 = 8'h8c == _match_key_qbytes_5_T_2 ? phv_data_140 : _GEN_3352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3354 = 8'h8d == _match_key_qbytes_5_T_2 ? phv_data_141 : _GEN_3353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3355 = 8'h8e == _match_key_qbytes_5_T_2 ? phv_data_142 : _GEN_3354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3356 = 8'h8f == _match_key_qbytes_5_T_2 ? phv_data_143 : _GEN_3355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3357 = 8'h90 == _match_key_qbytes_5_T_2 ? phv_data_144 : _GEN_3356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3358 = 8'h91 == _match_key_qbytes_5_T_2 ? phv_data_145 : _GEN_3357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3359 = 8'h92 == _match_key_qbytes_5_T_2 ? phv_data_146 : _GEN_3358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3360 = 8'h93 == _match_key_qbytes_5_T_2 ? phv_data_147 : _GEN_3359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3361 = 8'h94 == _match_key_qbytes_5_T_2 ? phv_data_148 : _GEN_3360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3362 = 8'h95 == _match_key_qbytes_5_T_2 ? phv_data_149 : _GEN_3361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3363 = 8'h96 == _match_key_qbytes_5_T_2 ? phv_data_150 : _GEN_3362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3364 = 8'h97 == _match_key_qbytes_5_T_2 ? phv_data_151 : _GEN_3363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3365 = 8'h98 == _match_key_qbytes_5_T_2 ? phv_data_152 : _GEN_3364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3366 = 8'h99 == _match_key_qbytes_5_T_2 ? phv_data_153 : _GEN_3365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3367 = 8'h9a == _match_key_qbytes_5_T_2 ? phv_data_154 : _GEN_3366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3368 = 8'h9b == _match_key_qbytes_5_T_2 ? phv_data_155 : _GEN_3367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3369 = 8'h9c == _match_key_qbytes_5_T_2 ? phv_data_156 : _GEN_3368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3370 = 8'h9d == _match_key_qbytes_5_T_2 ? phv_data_157 : _GEN_3369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3371 = 8'h9e == _match_key_qbytes_5_T_2 ? phv_data_158 : _GEN_3370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3372 = 8'h9f == _match_key_qbytes_5_T_2 ? phv_data_159 : _GEN_3371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3374 = 8'h1 == local_offset_5 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3375 = 8'h2 == local_offset_5 ? phv_data_2 : _GEN_3374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3376 = 8'h3 == local_offset_5 ? phv_data_3 : _GEN_3375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3377 = 8'h4 == local_offset_5 ? phv_data_4 : _GEN_3376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3378 = 8'h5 == local_offset_5 ? phv_data_5 : _GEN_3377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3379 = 8'h6 == local_offset_5 ? phv_data_6 : _GEN_3378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3380 = 8'h7 == local_offset_5 ? phv_data_7 : _GEN_3379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3381 = 8'h8 == local_offset_5 ? phv_data_8 : _GEN_3380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3382 = 8'h9 == local_offset_5 ? phv_data_9 : _GEN_3381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3383 = 8'ha == local_offset_5 ? phv_data_10 : _GEN_3382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3384 = 8'hb == local_offset_5 ? phv_data_11 : _GEN_3383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3385 = 8'hc == local_offset_5 ? phv_data_12 : _GEN_3384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3386 = 8'hd == local_offset_5 ? phv_data_13 : _GEN_3385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3387 = 8'he == local_offset_5 ? phv_data_14 : _GEN_3386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3388 = 8'hf == local_offset_5 ? phv_data_15 : _GEN_3387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3389 = 8'h10 == local_offset_5 ? phv_data_16 : _GEN_3388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3390 = 8'h11 == local_offset_5 ? phv_data_17 : _GEN_3389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3391 = 8'h12 == local_offset_5 ? phv_data_18 : _GEN_3390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3392 = 8'h13 == local_offset_5 ? phv_data_19 : _GEN_3391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3393 = 8'h14 == local_offset_5 ? phv_data_20 : _GEN_3392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3394 = 8'h15 == local_offset_5 ? phv_data_21 : _GEN_3393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3395 = 8'h16 == local_offset_5 ? phv_data_22 : _GEN_3394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3396 = 8'h17 == local_offset_5 ? phv_data_23 : _GEN_3395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3397 = 8'h18 == local_offset_5 ? phv_data_24 : _GEN_3396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3398 = 8'h19 == local_offset_5 ? phv_data_25 : _GEN_3397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3399 = 8'h1a == local_offset_5 ? phv_data_26 : _GEN_3398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3400 = 8'h1b == local_offset_5 ? phv_data_27 : _GEN_3399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3401 = 8'h1c == local_offset_5 ? phv_data_28 : _GEN_3400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3402 = 8'h1d == local_offset_5 ? phv_data_29 : _GEN_3401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3403 = 8'h1e == local_offset_5 ? phv_data_30 : _GEN_3402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3404 = 8'h1f == local_offset_5 ? phv_data_31 : _GEN_3403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3405 = 8'h20 == local_offset_5 ? phv_data_32 : _GEN_3404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3406 = 8'h21 == local_offset_5 ? phv_data_33 : _GEN_3405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3407 = 8'h22 == local_offset_5 ? phv_data_34 : _GEN_3406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3408 = 8'h23 == local_offset_5 ? phv_data_35 : _GEN_3407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3409 = 8'h24 == local_offset_5 ? phv_data_36 : _GEN_3408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3410 = 8'h25 == local_offset_5 ? phv_data_37 : _GEN_3409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3411 = 8'h26 == local_offset_5 ? phv_data_38 : _GEN_3410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3412 = 8'h27 == local_offset_5 ? phv_data_39 : _GEN_3411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3413 = 8'h28 == local_offset_5 ? phv_data_40 : _GEN_3412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3414 = 8'h29 == local_offset_5 ? phv_data_41 : _GEN_3413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3415 = 8'h2a == local_offset_5 ? phv_data_42 : _GEN_3414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3416 = 8'h2b == local_offset_5 ? phv_data_43 : _GEN_3415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3417 = 8'h2c == local_offset_5 ? phv_data_44 : _GEN_3416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3418 = 8'h2d == local_offset_5 ? phv_data_45 : _GEN_3417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3419 = 8'h2e == local_offset_5 ? phv_data_46 : _GEN_3418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3420 = 8'h2f == local_offset_5 ? phv_data_47 : _GEN_3419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3421 = 8'h30 == local_offset_5 ? phv_data_48 : _GEN_3420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3422 = 8'h31 == local_offset_5 ? phv_data_49 : _GEN_3421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3423 = 8'h32 == local_offset_5 ? phv_data_50 : _GEN_3422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3424 = 8'h33 == local_offset_5 ? phv_data_51 : _GEN_3423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3425 = 8'h34 == local_offset_5 ? phv_data_52 : _GEN_3424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3426 = 8'h35 == local_offset_5 ? phv_data_53 : _GEN_3425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3427 = 8'h36 == local_offset_5 ? phv_data_54 : _GEN_3426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3428 = 8'h37 == local_offset_5 ? phv_data_55 : _GEN_3427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3429 = 8'h38 == local_offset_5 ? phv_data_56 : _GEN_3428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3430 = 8'h39 == local_offset_5 ? phv_data_57 : _GEN_3429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3431 = 8'h3a == local_offset_5 ? phv_data_58 : _GEN_3430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3432 = 8'h3b == local_offset_5 ? phv_data_59 : _GEN_3431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3433 = 8'h3c == local_offset_5 ? phv_data_60 : _GEN_3432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3434 = 8'h3d == local_offset_5 ? phv_data_61 : _GEN_3433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3435 = 8'h3e == local_offset_5 ? phv_data_62 : _GEN_3434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3436 = 8'h3f == local_offset_5 ? phv_data_63 : _GEN_3435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3437 = 8'h40 == local_offset_5 ? phv_data_64 : _GEN_3436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3438 = 8'h41 == local_offset_5 ? phv_data_65 : _GEN_3437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3439 = 8'h42 == local_offset_5 ? phv_data_66 : _GEN_3438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3440 = 8'h43 == local_offset_5 ? phv_data_67 : _GEN_3439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3441 = 8'h44 == local_offset_5 ? phv_data_68 : _GEN_3440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3442 = 8'h45 == local_offset_5 ? phv_data_69 : _GEN_3441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3443 = 8'h46 == local_offset_5 ? phv_data_70 : _GEN_3442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3444 = 8'h47 == local_offset_5 ? phv_data_71 : _GEN_3443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3445 = 8'h48 == local_offset_5 ? phv_data_72 : _GEN_3444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3446 = 8'h49 == local_offset_5 ? phv_data_73 : _GEN_3445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3447 = 8'h4a == local_offset_5 ? phv_data_74 : _GEN_3446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3448 = 8'h4b == local_offset_5 ? phv_data_75 : _GEN_3447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3449 = 8'h4c == local_offset_5 ? phv_data_76 : _GEN_3448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3450 = 8'h4d == local_offset_5 ? phv_data_77 : _GEN_3449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3451 = 8'h4e == local_offset_5 ? phv_data_78 : _GEN_3450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3452 = 8'h4f == local_offset_5 ? phv_data_79 : _GEN_3451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3453 = 8'h50 == local_offset_5 ? phv_data_80 : _GEN_3452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3454 = 8'h51 == local_offset_5 ? phv_data_81 : _GEN_3453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3455 = 8'h52 == local_offset_5 ? phv_data_82 : _GEN_3454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3456 = 8'h53 == local_offset_5 ? phv_data_83 : _GEN_3455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3457 = 8'h54 == local_offset_5 ? phv_data_84 : _GEN_3456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3458 = 8'h55 == local_offset_5 ? phv_data_85 : _GEN_3457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3459 = 8'h56 == local_offset_5 ? phv_data_86 : _GEN_3458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3460 = 8'h57 == local_offset_5 ? phv_data_87 : _GEN_3459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3461 = 8'h58 == local_offset_5 ? phv_data_88 : _GEN_3460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3462 = 8'h59 == local_offset_5 ? phv_data_89 : _GEN_3461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3463 = 8'h5a == local_offset_5 ? phv_data_90 : _GEN_3462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3464 = 8'h5b == local_offset_5 ? phv_data_91 : _GEN_3463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3465 = 8'h5c == local_offset_5 ? phv_data_92 : _GEN_3464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3466 = 8'h5d == local_offset_5 ? phv_data_93 : _GEN_3465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3467 = 8'h5e == local_offset_5 ? phv_data_94 : _GEN_3466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3468 = 8'h5f == local_offset_5 ? phv_data_95 : _GEN_3467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3469 = 8'h60 == local_offset_5 ? phv_data_96 : _GEN_3468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3470 = 8'h61 == local_offset_5 ? phv_data_97 : _GEN_3469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3471 = 8'h62 == local_offset_5 ? phv_data_98 : _GEN_3470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3472 = 8'h63 == local_offset_5 ? phv_data_99 : _GEN_3471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3473 = 8'h64 == local_offset_5 ? phv_data_100 : _GEN_3472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3474 = 8'h65 == local_offset_5 ? phv_data_101 : _GEN_3473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3475 = 8'h66 == local_offset_5 ? phv_data_102 : _GEN_3474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3476 = 8'h67 == local_offset_5 ? phv_data_103 : _GEN_3475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3477 = 8'h68 == local_offset_5 ? phv_data_104 : _GEN_3476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3478 = 8'h69 == local_offset_5 ? phv_data_105 : _GEN_3477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3479 = 8'h6a == local_offset_5 ? phv_data_106 : _GEN_3478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3480 = 8'h6b == local_offset_5 ? phv_data_107 : _GEN_3479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3481 = 8'h6c == local_offset_5 ? phv_data_108 : _GEN_3480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3482 = 8'h6d == local_offset_5 ? phv_data_109 : _GEN_3481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3483 = 8'h6e == local_offset_5 ? phv_data_110 : _GEN_3482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3484 = 8'h6f == local_offset_5 ? phv_data_111 : _GEN_3483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3485 = 8'h70 == local_offset_5 ? phv_data_112 : _GEN_3484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3486 = 8'h71 == local_offset_5 ? phv_data_113 : _GEN_3485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3487 = 8'h72 == local_offset_5 ? phv_data_114 : _GEN_3486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3488 = 8'h73 == local_offset_5 ? phv_data_115 : _GEN_3487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3489 = 8'h74 == local_offset_5 ? phv_data_116 : _GEN_3488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3490 = 8'h75 == local_offset_5 ? phv_data_117 : _GEN_3489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3491 = 8'h76 == local_offset_5 ? phv_data_118 : _GEN_3490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3492 = 8'h77 == local_offset_5 ? phv_data_119 : _GEN_3491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3493 = 8'h78 == local_offset_5 ? phv_data_120 : _GEN_3492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3494 = 8'h79 == local_offset_5 ? phv_data_121 : _GEN_3493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3495 = 8'h7a == local_offset_5 ? phv_data_122 : _GEN_3494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3496 = 8'h7b == local_offset_5 ? phv_data_123 : _GEN_3495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3497 = 8'h7c == local_offset_5 ? phv_data_124 : _GEN_3496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3498 = 8'h7d == local_offset_5 ? phv_data_125 : _GEN_3497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3499 = 8'h7e == local_offset_5 ? phv_data_126 : _GEN_3498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3500 = 8'h7f == local_offset_5 ? phv_data_127 : _GEN_3499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3501 = 8'h80 == local_offset_5 ? phv_data_128 : _GEN_3500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3502 = 8'h81 == local_offset_5 ? phv_data_129 : _GEN_3501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3503 = 8'h82 == local_offset_5 ? phv_data_130 : _GEN_3502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3504 = 8'h83 == local_offset_5 ? phv_data_131 : _GEN_3503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3505 = 8'h84 == local_offset_5 ? phv_data_132 : _GEN_3504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3506 = 8'h85 == local_offset_5 ? phv_data_133 : _GEN_3505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3507 = 8'h86 == local_offset_5 ? phv_data_134 : _GEN_3506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3508 = 8'h87 == local_offset_5 ? phv_data_135 : _GEN_3507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3509 = 8'h88 == local_offset_5 ? phv_data_136 : _GEN_3508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3510 = 8'h89 == local_offset_5 ? phv_data_137 : _GEN_3509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3511 = 8'h8a == local_offset_5 ? phv_data_138 : _GEN_3510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3512 = 8'h8b == local_offset_5 ? phv_data_139 : _GEN_3511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3513 = 8'h8c == local_offset_5 ? phv_data_140 : _GEN_3512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3514 = 8'h8d == local_offset_5 ? phv_data_141 : _GEN_3513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3515 = 8'h8e == local_offset_5 ? phv_data_142 : _GEN_3514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3516 = 8'h8f == local_offset_5 ? phv_data_143 : _GEN_3515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3517 = 8'h90 == local_offset_5 ? phv_data_144 : _GEN_3516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3518 = 8'h91 == local_offset_5 ? phv_data_145 : _GEN_3517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3519 = 8'h92 == local_offset_5 ? phv_data_146 : _GEN_3518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3520 = 8'h93 == local_offset_5 ? phv_data_147 : _GEN_3519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3521 = 8'h94 == local_offset_5 ? phv_data_148 : _GEN_3520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3522 = 8'h95 == local_offset_5 ? phv_data_149 : _GEN_3521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3523 = 8'h96 == local_offset_5 ? phv_data_150 : _GEN_3522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3524 = 8'h97 == local_offset_5 ? phv_data_151 : _GEN_3523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3525 = 8'h98 == local_offset_5 ? phv_data_152 : _GEN_3524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3526 = 8'h99 == local_offset_5 ? phv_data_153 : _GEN_3525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3527 = 8'h9a == local_offset_5 ? phv_data_154 : _GEN_3526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3528 = 8'h9b == local_offset_5 ? phv_data_155 : _GEN_3527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3529 = 8'h9c == local_offset_5 ? phv_data_156 : _GEN_3528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3530 = 8'h9d == local_offset_5 ? phv_data_157 : _GEN_3529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3531 = 8'h9e == local_offset_5 ? phv_data_158 : _GEN_3530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3532 = 8'h9f == local_offset_5 ? phv_data_159 : _GEN_3531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3534 = 8'h1 == _match_key_qbytes_5_T ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3535 = 8'h2 == _match_key_qbytes_5_T ? phv_data_2 : _GEN_3534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3536 = 8'h3 == _match_key_qbytes_5_T ? phv_data_3 : _GEN_3535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3537 = 8'h4 == _match_key_qbytes_5_T ? phv_data_4 : _GEN_3536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3538 = 8'h5 == _match_key_qbytes_5_T ? phv_data_5 : _GEN_3537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3539 = 8'h6 == _match_key_qbytes_5_T ? phv_data_6 : _GEN_3538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3540 = 8'h7 == _match_key_qbytes_5_T ? phv_data_7 : _GEN_3539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3541 = 8'h8 == _match_key_qbytes_5_T ? phv_data_8 : _GEN_3540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3542 = 8'h9 == _match_key_qbytes_5_T ? phv_data_9 : _GEN_3541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3543 = 8'ha == _match_key_qbytes_5_T ? phv_data_10 : _GEN_3542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3544 = 8'hb == _match_key_qbytes_5_T ? phv_data_11 : _GEN_3543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3545 = 8'hc == _match_key_qbytes_5_T ? phv_data_12 : _GEN_3544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3546 = 8'hd == _match_key_qbytes_5_T ? phv_data_13 : _GEN_3545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3547 = 8'he == _match_key_qbytes_5_T ? phv_data_14 : _GEN_3546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3548 = 8'hf == _match_key_qbytes_5_T ? phv_data_15 : _GEN_3547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3549 = 8'h10 == _match_key_qbytes_5_T ? phv_data_16 : _GEN_3548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3550 = 8'h11 == _match_key_qbytes_5_T ? phv_data_17 : _GEN_3549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3551 = 8'h12 == _match_key_qbytes_5_T ? phv_data_18 : _GEN_3550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3552 = 8'h13 == _match_key_qbytes_5_T ? phv_data_19 : _GEN_3551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3553 = 8'h14 == _match_key_qbytes_5_T ? phv_data_20 : _GEN_3552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3554 = 8'h15 == _match_key_qbytes_5_T ? phv_data_21 : _GEN_3553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3555 = 8'h16 == _match_key_qbytes_5_T ? phv_data_22 : _GEN_3554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3556 = 8'h17 == _match_key_qbytes_5_T ? phv_data_23 : _GEN_3555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3557 = 8'h18 == _match_key_qbytes_5_T ? phv_data_24 : _GEN_3556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3558 = 8'h19 == _match_key_qbytes_5_T ? phv_data_25 : _GEN_3557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3559 = 8'h1a == _match_key_qbytes_5_T ? phv_data_26 : _GEN_3558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3560 = 8'h1b == _match_key_qbytes_5_T ? phv_data_27 : _GEN_3559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3561 = 8'h1c == _match_key_qbytes_5_T ? phv_data_28 : _GEN_3560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3562 = 8'h1d == _match_key_qbytes_5_T ? phv_data_29 : _GEN_3561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3563 = 8'h1e == _match_key_qbytes_5_T ? phv_data_30 : _GEN_3562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3564 = 8'h1f == _match_key_qbytes_5_T ? phv_data_31 : _GEN_3563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3565 = 8'h20 == _match_key_qbytes_5_T ? phv_data_32 : _GEN_3564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3566 = 8'h21 == _match_key_qbytes_5_T ? phv_data_33 : _GEN_3565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3567 = 8'h22 == _match_key_qbytes_5_T ? phv_data_34 : _GEN_3566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3568 = 8'h23 == _match_key_qbytes_5_T ? phv_data_35 : _GEN_3567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3569 = 8'h24 == _match_key_qbytes_5_T ? phv_data_36 : _GEN_3568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3570 = 8'h25 == _match_key_qbytes_5_T ? phv_data_37 : _GEN_3569; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3571 = 8'h26 == _match_key_qbytes_5_T ? phv_data_38 : _GEN_3570; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3572 = 8'h27 == _match_key_qbytes_5_T ? phv_data_39 : _GEN_3571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3573 = 8'h28 == _match_key_qbytes_5_T ? phv_data_40 : _GEN_3572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3574 = 8'h29 == _match_key_qbytes_5_T ? phv_data_41 : _GEN_3573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3575 = 8'h2a == _match_key_qbytes_5_T ? phv_data_42 : _GEN_3574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3576 = 8'h2b == _match_key_qbytes_5_T ? phv_data_43 : _GEN_3575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3577 = 8'h2c == _match_key_qbytes_5_T ? phv_data_44 : _GEN_3576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3578 = 8'h2d == _match_key_qbytes_5_T ? phv_data_45 : _GEN_3577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3579 = 8'h2e == _match_key_qbytes_5_T ? phv_data_46 : _GEN_3578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3580 = 8'h2f == _match_key_qbytes_5_T ? phv_data_47 : _GEN_3579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3581 = 8'h30 == _match_key_qbytes_5_T ? phv_data_48 : _GEN_3580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3582 = 8'h31 == _match_key_qbytes_5_T ? phv_data_49 : _GEN_3581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3583 = 8'h32 == _match_key_qbytes_5_T ? phv_data_50 : _GEN_3582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3584 = 8'h33 == _match_key_qbytes_5_T ? phv_data_51 : _GEN_3583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3585 = 8'h34 == _match_key_qbytes_5_T ? phv_data_52 : _GEN_3584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3586 = 8'h35 == _match_key_qbytes_5_T ? phv_data_53 : _GEN_3585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3587 = 8'h36 == _match_key_qbytes_5_T ? phv_data_54 : _GEN_3586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3588 = 8'h37 == _match_key_qbytes_5_T ? phv_data_55 : _GEN_3587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3589 = 8'h38 == _match_key_qbytes_5_T ? phv_data_56 : _GEN_3588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3590 = 8'h39 == _match_key_qbytes_5_T ? phv_data_57 : _GEN_3589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3591 = 8'h3a == _match_key_qbytes_5_T ? phv_data_58 : _GEN_3590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3592 = 8'h3b == _match_key_qbytes_5_T ? phv_data_59 : _GEN_3591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3593 = 8'h3c == _match_key_qbytes_5_T ? phv_data_60 : _GEN_3592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3594 = 8'h3d == _match_key_qbytes_5_T ? phv_data_61 : _GEN_3593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3595 = 8'h3e == _match_key_qbytes_5_T ? phv_data_62 : _GEN_3594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3596 = 8'h3f == _match_key_qbytes_5_T ? phv_data_63 : _GEN_3595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3597 = 8'h40 == _match_key_qbytes_5_T ? phv_data_64 : _GEN_3596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3598 = 8'h41 == _match_key_qbytes_5_T ? phv_data_65 : _GEN_3597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3599 = 8'h42 == _match_key_qbytes_5_T ? phv_data_66 : _GEN_3598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3600 = 8'h43 == _match_key_qbytes_5_T ? phv_data_67 : _GEN_3599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3601 = 8'h44 == _match_key_qbytes_5_T ? phv_data_68 : _GEN_3600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3602 = 8'h45 == _match_key_qbytes_5_T ? phv_data_69 : _GEN_3601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3603 = 8'h46 == _match_key_qbytes_5_T ? phv_data_70 : _GEN_3602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3604 = 8'h47 == _match_key_qbytes_5_T ? phv_data_71 : _GEN_3603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3605 = 8'h48 == _match_key_qbytes_5_T ? phv_data_72 : _GEN_3604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3606 = 8'h49 == _match_key_qbytes_5_T ? phv_data_73 : _GEN_3605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3607 = 8'h4a == _match_key_qbytes_5_T ? phv_data_74 : _GEN_3606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3608 = 8'h4b == _match_key_qbytes_5_T ? phv_data_75 : _GEN_3607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3609 = 8'h4c == _match_key_qbytes_5_T ? phv_data_76 : _GEN_3608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3610 = 8'h4d == _match_key_qbytes_5_T ? phv_data_77 : _GEN_3609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3611 = 8'h4e == _match_key_qbytes_5_T ? phv_data_78 : _GEN_3610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3612 = 8'h4f == _match_key_qbytes_5_T ? phv_data_79 : _GEN_3611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3613 = 8'h50 == _match_key_qbytes_5_T ? phv_data_80 : _GEN_3612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3614 = 8'h51 == _match_key_qbytes_5_T ? phv_data_81 : _GEN_3613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3615 = 8'h52 == _match_key_qbytes_5_T ? phv_data_82 : _GEN_3614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3616 = 8'h53 == _match_key_qbytes_5_T ? phv_data_83 : _GEN_3615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3617 = 8'h54 == _match_key_qbytes_5_T ? phv_data_84 : _GEN_3616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3618 = 8'h55 == _match_key_qbytes_5_T ? phv_data_85 : _GEN_3617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3619 = 8'h56 == _match_key_qbytes_5_T ? phv_data_86 : _GEN_3618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3620 = 8'h57 == _match_key_qbytes_5_T ? phv_data_87 : _GEN_3619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3621 = 8'h58 == _match_key_qbytes_5_T ? phv_data_88 : _GEN_3620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3622 = 8'h59 == _match_key_qbytes_5_T ? phv_data_89 : _GEN_3621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3623 = 8'h5a == _match_key_qbytes_5_T ? phv_data_90 : _GEN_3622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3624 = 8'h5b == _match_key_qbytes_5_T ? phv_data_91 : _GEN_3623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3625 = 8'h5c == _match_key_qbytes_5_T ? phv_data_92 : _GEN_3624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3626 = 8'h5d == _match_key_qbytes_5_T ? phv_data_93 : _GEN_3625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3627 = 8'h5e == _match_key_qbytes_5_T ? phv_data_94 : _GEN_3626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3628 = 8'h5f == _match_key_qbytes_5_T ? phv_data_95 : _GEN_3627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3629 = 8'h60 == _match_key_qbytes_5_T ? phv_data_96 : _GEN_3628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3630 = 8'h61 == _match_key_qbytes_5_T ? phv_data_97 : _GEN_3629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3631 = 8'h62 == _match_key_qbytes_5_T ? phv_data_98 : _GEN_3630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3632 = 8'h63 == _match_key_qbytes_5_T ? phv_data_99 : _GEN_3631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3633 = 8'h64 == _match_key_qbytes_5_T ? phv_data_100 : _GEN_3632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3634 = 8'h65 == _match_key_qbytes_5_T ? phv_data_101 : _GEN_3633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3635 = 8'h66 == _match_key_qbytes_5_T ? phv_data_102 : _GEN_3634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3636 = 8'h67 == _match_key_qbytes_5_T ? phv_data_103 : _GEN_3635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3637 = 8'h68 == _match_key_qbytes_5_T ? phv_data_104 : _GEN_3636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3638 = 8'h69 == _match_key_qbytes_5_T ? phv_data_105 : _GEN_3637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3639 = 8'h6a == _match_key_qbytes_5_T ? phv_data_106 : _GEN_3638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3640 = 8'h6b == _match_key_qbytes_5_T ? phv_data_107 : _GEN_3639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3641 = 8'h6c == _match_key_qbytes_5_T ? phv_data_108 : _GEN_3640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3642 = 8'h6d == _match_key_qbytes_5_T ? phv_data_109 : _GEN_3641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3643 = 8'h6e == _match_key_qbytes_5_T ? phv_data_110 : _GEN_3642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3644 = 8'h6f == _match_key_qbytes_5_T ? phv_data_111 : _GEN_3643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3645 = 8'h70 == _match_key_qbytes_5_T ? phv_data_112 : _GEN_3644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3646 = 8'h71 == _match_key_qbytes_5_T ? phv_data_113 : _GEN_3645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3647 = 8'h72 == _match_key_qbytes_5_T ? phv_data_114 : _GEN_3646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3648 = 8'h73 == _match_key_qbytes_5_T ? phv_data_115 : _GEN_3647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3649 = 8'h74 == _match_key_qbytes_5_T ? phv_data_116 : _GEN_3648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3650 = 8'h75 == _match_key_qbytes_5_T ? phv_data_117 : _GEN_3649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3651 = 8'h76 == _match_key_qbytes_5_T ? phv_data_118 : _GEN_3650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3652 = 8'h77 == _match_key_qbytes_5_T ? phv_data_119 : _GEN_3651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3653 = 8'h78 == _match_key_qbytes_5_T ? phv_data_120 : _GEN_3652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3654 = 8'h79 == _match_key_qbytes_5_T ? phv_data_121 : _GEN_3653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3655 = 8'h7a == _match_key_qbytes_5_T ? phv_data_122 : _GEN_3654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3656 = 8'h7b == _match_key_qbytes_5_T ? phv_data_123 : _GEN_3655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3657 = 8'h7c == _match_key_qbytes_5_T ? phv_data_124 : _GEN_3656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3658 = 8'h7d == _match_key_qbytes_5_T ? phv_data_125 : _GEN_3657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3659 = 8'h7e == _match_key_qbytes_5_T ? phv_data_126 : _GEN_3658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3660 = 8'h7f == _match_key_qbytes_5_T ? phv_data_127 : _GEN_3659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3661 = 8'h80 == _match_key_qbytes_5_T ? phv_data_128 : _GEN_3660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3662 = 8'h81 == _match_key_qbytes_5_T ? phv_data_129 : _GEN_3661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3663 = 8'h82 == _match_key_qbytes_5_T ? phv_data_130 : _GEN_3662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3664 = 8'h83 == _match_key_qbytes_5_T ? phv_data_131 : _GEN_3663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3665 = 8'h84 == _match_key_qbytes_5_T ? phv_data_132 : _GEN_3664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3666 = 8'h85 == _match_key_qbytes_5_T ? phv_data_133 : _GEN_3665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3667 = 8'h86 == _match_key_qbytes_5_T ? phv_data_134 : _GEN_3666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3668 = 8'h87 == _match_key_qbytes_5_T ? phv_data_135 : _GEN_3667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3669 = 8'h88 == _match_key_qbytes_5_T ? phv_data_136 : _GEN_3668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3670 = 8'h89 == _match_key_qbytes_5_T ? phv_data_137 : _GEN_3669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3671 = 8'h8a == _match_key_qbytes_5_T ? phv_data_138 : _GEN_3670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3672 = 8'h8b == _match_key_qbytes_5_T ? phv_data_139 : _GEN_3671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3673 = 8'h8c == _match_key_qbytes_5_T ? phv_data_140 : _GEN_3672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3674 = 8'h8d == _match_key_qbytes_5_T ? phv_data_141 : _GEN_3673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3675 = 8'h8e == _match_key_qbytes_5_T ? phv_data_142 : _GEN_3674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3676 = 8'h8f == _match_key_qbytes_5_T ? phv_data_143 : _GEN_3675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3677 = 8'h90 == _match_key_qbytes_5_T ? phv_data_144 : _GEN_3676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3678 = 8'h91 == _match_key_qbytes_5_T ? phv_data_145 : _GEN_3677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3679 = 8'h92 == _match_key_qbytes_5_T ? phv_data_146 : _GEN_3678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3680 = 8'h93 == _match_key_qbytes_5_T ? phv_data_147 : _GEN_3679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3681 = 8'h94 == _match_key_qbytes_5_T ? phv_data_148 : _GEN_3680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3682 = 8'h95 == _match_key_qbytes_5_T ? phv_data_149 : _GEN_3681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3683 = 8'h96 == _match_key_qbytes_5_T ? phv_data_150 : _GEN_3682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3684 = 8'h97 == _match_key_qbytes_5_T ? phv_data_151 : _GEN_3683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3685 = 8'h98 == _match_key_qbytes_5_T ? phv_data_152 : _GEN_3684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3686 = 8'h99 == _match_key_qbytes_5_T ? phv_data_153 : _GEN_3685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3687 = 8'h9a == _match_key_qbytes_5_T ? phv_data_154 : _GEN_3686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3688 = 8'h9b == _match_key_qbytes_5_T ? phv_data_155 : _GEN_3687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3689 = 8'h9c == _match_key_qbytes_5_T ? phv_data_156 : _GEN_3688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3690 = 8'h9d == _match_key_qbytes_5_T ? phv_data_157 : _GEN_3689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3691 = 8'h9e == _match_key_qbytes_5_T ? phv_data_158 : _GEN_3690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3692 = 8'h9f == _match_key_qbytes_5_T ? phv_data_159 : _GEN_3691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3694 = 8'h1 == _match_key_qbytes_5_T_1 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3695 = 8'h2 == _match_key_qbytes_5_T_1 ? phv_data_2 : _GEN_3694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3696 = 8'h3 == _match_key_qbytes_5_T_1 ? phv_data_3 : _GEN_3695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3697 = 8'h4 == _match_key_qbytes_5_T_1 ? phv_data_4 : _GEN_3696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3698 = 8'h5 == _match_key_qbytes_5_T_1 ? phv_data_5 : _GEN_3697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3699 = 8'h6 == _match_key_qbytes_5_T_1 ? phv_data_6 : _GEN_3698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3700 = 8'h7 == _match_key_qbytes_5_T_1 ? phv_data_7 : _GEN_3699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3701 = 8'h8 == _match_key_qbytes_5_T_1 ? phv_data_8 : _GEN_3700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3702 = 8'h9 == _match_key_qbytes_5_T_1 ? phv_data_9 : _GEN_3701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3703 = 8'ha == _match_key_qbytes_5_T_1 ? phv_data_10 : _GEN_3702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3704 = 8'hb == _match_key_qbytes_5_T_1 ? phv_data_11 : _GEN_3703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3705 = 8'hc == _match_key_qbytes_5_T_1 ? phv_data_12 : _GEN_3704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3706 = 8'hd == _match_key_qbytes_5_T_1 ? phv_data_13 : _GEN_3705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3707 = 8'he == _match_key_qbytes_5_T_1 ? phv_data_14 : _GEN_3706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3708 = 8'hf == _match_key_qbytes_5_T_1 ? phv_data_15 : _GEN_3707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3709 = 8'h10 == _match_key_qbytes_5_T_1 ? phv_data_16 : _GEN_3708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3710 = 8'h11 == _match_key_qbytes_5_T_1 ? phv_data_17 : _GEN_3709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3711 = 8'h12 == _match_key_qbytes_5_T_1 ? phv_data_18 : _GEN_3710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3712 = 8'h13 == _match_key_qbytes_5_T_1 ? phv_data_19 : _GEN_3711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3713 = 8'h14 == _match_key_qbytes_5_T_1 ? phv_data_20 : _GEN_3712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3714 = 8'h15 == _match_key_qbytes_5_T_1 ? phv_data_21 : _GEN_3713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3715 = 8'h16 == _match_key_qbytes_5_T_1 ? phv_data_22 : _GEN_3714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3716 = 8'h17 == _match_key_qbytes_5_T_1 ? phv_data_23 : _GEN_3715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3717 = 8'h18 == _match_key_qbytes_5_T_1 ? phv_data_24 : _GEN_3716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3718 = 8'h19 == _match_key_qbytes_5_T_1 ? phv_data_25 : _GEN_3717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3719 = 8'h1a == _match_key_qbytes_5_T_1 ? phv_data_26 : _GEN_3718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3720 = 8'h1b == _match_key_qbytes_5_T_1 ? phv_data_27 : _GEN_3719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3721 = 8'h1c == _match_key_qbytes_5_T_1 ? phv_data_28 : _GEN_3720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3722 = 8'h1d == _match_key_qbytes_5_T_1 ? phv_data_29 : _GEN_3721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3723 = 8'h1e == _match_key_qbytes_5_T_1 ? phv_data_30 : _GEN_3722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3724 = 8'h1f == _match_key_qbytes_5_T_1 ? phv_data_31 : _GEN_3723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3725 = 8'h20 == _match_key_qbytes_5_T_1 ? phv_data_32 : _GEN_3724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3726 = 8'h21 == _match_key_qbytes_5_T_1 ? phv_data_33 : _GEN_3725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3727 = 8'h22 == _match_key_qbytes_5_T_1 ? phv_data_34 : _GEN_3726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3728 = 8'h23 == _match_key_qbytes_5_T_1 ? phv_data_35 : _GEN_3727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3729 = 8'h24 == _match_key_qbytes_5_T_1 ? phv_data_36 : _GEN_3728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3730 = 8'h25 == _match_key_qbytes_5_T_1 ? phv_data_37 : _GEN_3729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3731 = 8'h26 == _match_key_qbytes_5_T_1 ? phv_data_38 : _GEN_3730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3732 = 8'h27 == _match_key_qbytes_5_T_1 ? phv_data_39 : _GEN_3731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3733 = 8'h28 == _match_key_qbytes_5_T_1 ? phv_data_40 : _GEN_3732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3734 = 8'h29 == _match_key_qbytes_5_T_1 ? phv_data_41 : _GEN_3733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3735 = 8'h2a == _match_key_qbytes_5_T_1 ? phv_data_42 : _GEN_3734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3736 = 8'h2b == _match_key_qbytes_5_T_1 ? phv_data_43 : _GEN_3735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3737 = 8'h2c == _match_key_qbytes_5_T_1 ? phv_data_44 : _GEN_3736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3738 = 8'h2d == _match_key_qbytes_5_T_1 ? phv_data_45 : _GEN_3737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3739 = 8'h2e == _match_key_qbytes_5_T_1 ? phv_data_46 : _GEN_3738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3740 = 8'h2f == _match_key_qbytes_5_T_1 ? phv_data_47 : _GEN_3739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3741 = 8'h30 == _match_key_qbytes_5_T_1 ? phv_data_48 : _GEN_3740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3742 = 8'h31 == _match_key_qbytes_5_T_1 ? phv_data_49 : _GEN_3741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3743 = 8'h32 == _match_key_qbytes_5_T_1 ? phv_data_50 : _GEN_3742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3744 = 8'h33 == _match_key_qbytes_5_T_1 ? phv_data_51 : _GEN_3743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3745 = 8'h34 == _match_key_qbytes_5_T_1 ? phv_data_52 : _GEN_3744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3746 = 8'h35 == _match_key_qbytes_5_T_1 ? phv_data_53 : _GEN_3745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3747 = 8'h36 == _match_key_qbytes_5_T_1 ? phv_data_54 : _GEN_3746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3748 = 8'h37 == _match_key_qbytes_5_T_1 ? phv_data_55 : _GEN_3747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3749 = 8'h38 == _match_key_qbytes_5_T_1 ? phv_data_56 : _GEN_3748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3750 = 8'h39 == _match_key_qbytes_5_T_1 ? phv_data_57 : _GEN_3749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3751 = 8'h3a == _match_key_qbytes_5_T_1 ? phv_data_58 : _GEN_3750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3752 = 8'h3b == _match_key_qbytes_5_T_1 ? phv_data_59 : _GEN_3751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3753 = 8'h3c == _match_key_qbytes_5_T_1 ? phv_data_60 : _GEN_3752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3754 = 8'h3d == _match_key_qbytes_5_T_1 ? phv_data_61 : _GEN_3753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3755 = 8'h3e == _match_key_qbytes_5_T_1 ? phv_data_62 : _GEN_3754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3756 = 8'h3f == _match_key_qbytes_5_T_1 ? phv_data_63 : _GEN_3755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3757 = 8'h40 == _match_key_qbytes_5_T_1 ? phv_data_64 : _GEN_3756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3758 = 8'h41 == _match_key_qbytes_5_T_1 ? phv_data_65 : _GEN_3757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3759 = 8'h42 == _match_key_qbytes_5_T_1 ? phv_data_66 : _GEN_3758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3760 = 8'h43 == _match_key_qbytes_5_T_1 ? phv_data_67 : _GEN_3759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3761 = 8'h44 == _match_key_qbytes_5_T_1 ? phv_data_68 : _GEN_3760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3762 = 8'h45 == _match_key_qbytes_5_T_1 ? phv_data_69 : _GEN_3761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3763 = 8'h46 == _match_key_qbytes_5_T_1 ? phv_data_70 : _GEN_3762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3764 = 8'h47 == _match_key_qbytes_5_T_1 ? phv_data_71 : _GEN_3763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3765 = 8'h48 == _match_key_qbytes_5_T_1 ? phv_data_72 : _GEN_3764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3766 = 8'h49 == _match_key_qbytes_5_T_1 ? phv_data_73 : _GEN_3765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3767 = 8'h4a == _match_key_qbytes_5_T_1 ? phv_data_74 : _GEN_3766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3768 = 8'h4b == _match_key_qbytes_5_T_1 ? phv_data_75 : _GEN_3767; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3769 = 8'h4c == _match_key_qbytes_5_T_1 ? phv_data_76 : _GEN_3768; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3770 = 8'h4d == _match_key_qbytes_5_T_1 ? phv_data_77 : _GEN_3769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3771 = 8'h4e == _match_key_qbytes_5_T_1 ? phv_data_78 : _GEN_3770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3772 = 8'h4f == _match_key_qbytes_5_T_1 ? phv_data_79 : _GEN_3771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3773 = 8'h50 == _match_key_qbytes_5_T_1 ? phv_data_80 : _GEN_3772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3774 = 8'h51 == _match_key_qbytes_5_T_1 ? phv_data_81 : _GEN_3773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3775 = 8'h52 == _match_key_qbytes_5_T_1 ? phv_data_82 : _GEN_3774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3776 = 8'h53 == _match_key_qbytes_5_T_1 ? phv_data_83 : _GEN_3775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3777 = 8'h54 == _match_key_qbytes_5_T_1 ? phv_data_84 : _GEN_3776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3778 = 8'h55 == _match_key_qbytes_5_T_1 ? phv_data_85 : _GEN_3777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3779 = 8'h56 == _match_key_qbytes_5_T_1 ? phv_data_86 : _GEN_3778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3780 = 8'h57 == _match_key_qbytes_5_T_1 ? phv_data_87 : _GEN_3779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3781 = 8'h58 == _match_key_qbytes_5_T_1 ? phv_data_88 : _GEN_3780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3782 = 8'h59 == _match_key_qbytes_5_T_1 ? phv_data_89 : _GEN_3781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3783 = 8'h5a == _match_key_qbytes_5_T_1 ? phv_data_90 : _GEN_3782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3784 = 8'h5b == _match_key_qbytes_5_T_1 ? phv_data_91 : _GEN_3783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3785 = 8'h5c == _match_key_qbytes_5_T_1 ? phv_data_92 : _GEN_3784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3786 = 8'h5d == _match_key_qbytes_5_T_1 ? phv_data_93 : _GEN_3785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3787 = 8'h5e == _match_key_qbytes_5_T_1 ? phv_data_94 : _GEN_3786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3788 = 8'h5f == _match_key_qbytes_5_T_1 ? phv_data_95 : _GEN_3787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3789 = 8'h60 == _match_key_qbytes_5_T_1 ? phv_data_96 : _GEN_3788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3790 = 8'h61 == _match_key_qbytes_5_T_1 ? phv_data_97 : _GEN_3789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3791 = 8'h62 == _match_key_qbytes_5_T_1 ? phv_data_98 : _GEN_3790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3792 = 8'h63 == _match_key_qbytes_5_T_1 ? phv_data_99 : _GEN_3791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3793 = 8'h64 == _match_key_qbytes_5_T_1 ? phv_data_100 : _GEN_3792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3794 = 8'h65 == _match_key_qbytes_5_T_1 ? phv_data_101 : _GEN_3793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3795 = 8'h66 == _match_key_qbytes_5_T_1 ? phv_data_102 : _GEN_3794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3796 = 8'h67 == _match_key_qbytes_5_T_1 ? phv_data_103 : _GEN_3795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3797 = 8'h68 == _match_key_qbytes_5_T_1 ? phv_data_104 : _GEN_3796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3798 = 8'h69 == _match_key_qbytes_5_T_1 ? phv_data_105 : _GEN_3797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3799 = 8'h6a == _match_key_qbytes_5_T_1 ? phv_data_106 : _GEN_3798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3800 = 8'h6b == _match_key_qbytes_5_T_1 ? phv_data_107 : _GEN_3799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3801 = 8'h6c == _match_key_qbytes_5_T_1 ? phv_data_108 : _GEN_3800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3802 = 8'h6d == _match_key_qbytes_5_T_1 ? phv_data_109 : _GEN_3801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3803 = 8'h6e == _match_key_qbytes_5_T_1 ? phv_data_110 : _GEN_3802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3804 = 8'h6f == _match_key_qbytes_5_T_1 ? phv_data_111 : _GEN_3803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3805 = 8'h70 == _match_key_qbytes_5_T_1 ? phv_data_112 : _GEN_3804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3806 = 8'h71 == _match_key_qbytes_5_T_1 ? phv_data_113 : _GEN_3805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3807 = 8'h72 == _match_key_qbytes_5_T_1 ? phv_data_114 : _GEN_3806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3808 = 8'h73 == _match_key_qbytes_5_T_1 ? phv_data_115 : _GEN_3807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3809 = 8'h74 == _match_key_qbytes_5_T_1 ? phv_data_116 : _GEN_3808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3810 = 8'h75 == _match_key_qbytes_5_T_1 ? phv_data_117 : _GEN_3809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3811 = 8'h76 == _match_key_qbytes_5_T_1 ? phv_data_118 : _GEN_3810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3812 = 8'h77 == _match_key_qbytes_5_T_1 ? phv_data_119 : _GEN_3811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3813 = 8'h78 == _match_key_qbytes_5_T_1 ? phv_data_120 : _GEN_3812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3814 = 8'h79 == _match_key_qbytes_5_T_1 ? phv_data_121 : _GEN_3813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3815 = 8'h7a == _match_key_qbytes_5_T_1 ? phv_data_122 : _GEN_3814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3816 = 8'h7b == _match_key_qbytes_5_T_1 ? phv_data_123 : _GEN_3815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3817 = 8'h7c == _match_key_qbytes_5_T_1 ? phv_data_124 : _GEN_3816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3818 = 8'h7d == _match_key_qbytes_5_T_1 ? phv_data_125 : _GEN_3817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3819 = 8'h7e == _match_key_qbytes_5_T_1 ? phv_data_126 : _GEN_3818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3820 = 8'h7f == _match_key_qbytes_5_T_1 ? phv_data_127 : _GEN_3819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3821 = 8'h80 == _match_key_qbytes_5_T_1 ? phv_data_128 : _GEN_3820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3822 = 8'h81 == _match_key_qbytes_5_T_1 ? phv_data_129 : _GEN_3821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3823 = 8'h82 == _match_key_qbytes_5_T_1 ? phv_data_130 : _GEN_3822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3824 = 8'h83 == _match_key_qbytes_5_T_1 ? phv_data_131 : _GEN_3823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3825 = 8'h84 == _match_key_qbytes_5_T_1 ? phv_data_132 : _GEN_3824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3826 = 8'h85 == _match_key_qbytes_5_T_1 ? phv_data_133 : _GEN_3825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3827 = 8'h86 == _match_key_qbytes_5_T_1 ? phv_data_134 : _GEN_3826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3828 = 8'h87 == _match_key_qbytes_5_T_1 ? phv_data_135 : _GEN_3827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3829 = 8'h88 == _match_key_qbytes_5_T_1 ? phv_data_136 : _GEN_3828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3830 = 8'h89 == _match_key_qbytes_5_T_1 ? phv_data_137 : _GEN_3829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3831 = 8'h8a == _match_key_qbytes_5_T_1 ? phv_data_138 : _GEN_3830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3832 = 8'h8b == _match_key_qbytes_5_T_1 ? phv_data_139 : _GEN_3831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3833 = 8'h8c == _match_key_qbytes_5_T_1 ? phv_data_140 : _GEN_3832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3834 = 8'h8d == _match_key_qbytes_5_T_1 ? phv_data_141 : _GEN_3833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3835 = 8'h8e == _match_key_qbytes_5_T_1 ? phv_data_142 : _GEN_3834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3836 = 8'h8f == _match_key_qbytes_5_T_1 ? phv_data_143 : _GEN_3835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3837 = 8'h90 == _match_key_qbytes_5_T_1 ? phv_data_144 : _GEN_3836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3838 = 8'h91 == _match_key_qbytes_5_T_1 ? phv_data_145 : _GEN_3837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3839 = 8'h92 == _match_key_qbytes_5_T_1 ? phv_data_146 : _GEN_3838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3840 = 8'h93 == _match_key_qbytes_5_T_1 ? phv_data_147 : _GEN_3839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3841 = 8'h94 == _match_key_qbytes_5_T_1 ? phv_data_148 : _GEN_3840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3842 = 8'h95 == _match_key_qbytes_5_T_1 ? phv_data_149 : _GEN_3841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3843 = 8'h96 == _match_key_qbytes_5_T_1 ? phv_data_150 : _GEN_3842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3844 = 8'h97 == _match_key_qbytes_5_T_1 ? phv_data_151 : _GEN_3843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3845 = 8'h98 == _match_key_qbytes_5_T_1 ? phv_data_152 : _GEN_3844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3846 = 8'h99 == _match_key_qbytes_5_T_1 ? phv_data_153 : _GEN_3845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3847 = 8'h9a == _match_key_qbytes_5_T_1 ? phv_data_154 : _GEN_3846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3848 = 8'h9b == _match_key_qbytes_5_T_1 ? phv_data_155 : _GEN_3847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3849 = 8'h9c == _match_key_qbytes_5_T_1 ? phv_data_156 : _GEN_3848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3850 = 8'h9d == _match_key_qbytes_5_T_1 ? phv_data_157 : _GEN_3849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3851 = 8'h9e == _match_key_qbytes_5_T_1 ? phv_data_158 : _GEN_3850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3852 = 8'h9f == _match_key_qbytes_5_T_1 ? phv_data_159 : _GEN_3851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [31:0] _match_key_qbytes_5_T_3 = {_GEN_3692,_GEN_3852,_GEN_3372,_GEN_3532}; // @[Cat.scala 30:58]
  wire [31:0] match_key_qbytes_5 = local_offset_5 < end_offset ? _match_key_qbytes_5_T_3 : 32'h0; // @[matcher.scala 88:54 matcher.scala 89:45 matcher.scala 97:45]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_96 = phv_data_96; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_97 = phv_data_97; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_98 = phv_data_98; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_99 = phv_data_99; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_100 = phv_data_100; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_101 = phv_data_101; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_102 = phv_data_102; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_103 = phv_data_103; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_104 = phv_data_104; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_105 = phv_data_105; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_106 = phv_data_106; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_107 = phv_data_107; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_108 = phv_data_108; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_109 = phv_data_109; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_110 = phv_data_110; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_111 = phv_data_111; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_112 = phv_data_112; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_113 = phv_data_113; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_114 = phv_data_114; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_115 = phv_data_115; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_116 = phv_data_116; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_117 = phv_data_117; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_118 = phv_data_118; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_119 = phv_data_119; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_120 = phv_data_120; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_121 = phv_data_121; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_122 = phv_data_122; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_123 = phv_data_123; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_124 = phv_data_124; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_125 = phv_data_125; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_126 = phv_data_126; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_127 = phv_data_127; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_128 = phv_data_128; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_129 = phv_data_129; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_130 = phv_data_130; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_131 = phv_data_131; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_132 = phv_data_132; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_133 = phv_data_133; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_134 = phv_data_134; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_135 = phv_data_135; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_136 = phv_data_136; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_137 = phv_data_137; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_138 = phv_data_138; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_139 = phv_data_139; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_140 = phv_data_140; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_141 = phv_data_141; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_142 = phv_data_142; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_143 = phv_data_143; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_144 = phv_data_144; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_145 = phv_data_145; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_146 = phv_data_146; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_147 = phv_data_147; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_148 = phv_data_148; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_149 = phv_data_149; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_150 = phv_data_150; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_151 = phv_data_151; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_152 = phv_data_152; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_153 = phv_data_153; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_154 = phv_data_154; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_155 = phv_data_155; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_156 = phv_data_156; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_157 = phv_data_157; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_158 = phv_data_158; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_159 = phv_data_159; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[matcher.scala 69:29]
  assign io_bias_out = key_offset[1:0]; // @[matcher.scala 79:38]
  assign io_match_key_bytes_0 = phv_is_valid_processor ? match_key_qbytes_0[7:0] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_1 = phv_is_valid_processor ? match_key_qbytes_0[15:8] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_2 = phv_is_valid_processor ? match_key_qbytes_0[23:16] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_3 = phv_is_valid_processor ? match_key_qbytes_0[31:24] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_4 = phv_is_valid_processor ? match_key_qbytes_1[7:0] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_5 = phv_is_valid_processor ? match_key_qbytes_1[15:8] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_6 = phv_is_valid_processor ? match_key_qbytes_1[23:16] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_7 = phv_is_valid_processor ? match_key_qbytes_1[31:24] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_8 = phv_is_valid_processor ? match_key_qbytes_2[7:0] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_9 = phv_is_valid_processor ? match_key_qbytes_2[15:8] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_10 = phv_is_valid_processor ? match_key_qbytes_2[23:16] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_11 = phv_is_valid_processor ? match_key_qbytes_2[31:24] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_12 = phv_is_valid_processor ? match_key_qbytes_3[7:0] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_13 = phv_is_valid_processor ? match_key_qbytes_3[15:8] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_14 = phv_is_valid_processor ? match_key_qbytes_3[23:16] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_15 = phv_is_valid_processor ? match_key_qbytes_3[31:24] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_16 = phv_is_valid_processor ? match_key_qbytes_4[7:0] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_17 = phv_is_valid_processor ? match_key_qbytes_4[15:8] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_18 = phv_is_valid_processor ? match_key_qbytes_4[23:16] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_19 = phv_is_valid_processor ? match_key_qbytes_4[31:24] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_20 = phv_is_valid_processor ? match_key_qbytes_5[7:0] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_21 = phv_is_valid_processor ? match_key_qbytes_5[15:8] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_22 = phv_is_valid_processor ? match_key_qbytes_5[23:16] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_23 = phv_is_valid_processor ? match_key_qbytes_5[31:24] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[matcher.scala 68:17]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[matcher.scala 68:17]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[matcher.scala 68:17]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[matcher.scala 68:17]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[matcher.scala 68:17]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[matcher.scala 68:17]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[matcher.scala 68:17]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[matcher.scala 68:17]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[matcher.scala 68:17]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[matcher.scala 68:17]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[matcher.scala 68:17]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[matcher.scala 68:17]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[matcher.scala 68:17]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[matcher.scala 68:17]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[matcher.scala 68:17]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[matcher.scala 68:17]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[matcher.scala 68:17]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[matcher.scala 68:17]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[matcher.scala 68:17]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[matcher.scala 68:17]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[matcher.scala 68:17]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[matcher.scala 68:17]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[matcher.scala 68:17]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[matcher.scala 68:17]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[matcher.scala 68:17]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[matcher.scala 68:17]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[matcher.scala 68:17]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[matcher.scala 68:17]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[matcher.scala 68:17]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[matcher.scala 68:17]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[matcher.scala 68:17]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[matcher.scala 68:17]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[matcher.scala 68:17]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[matcher.scala 68:17]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[matcher.scala 68:17]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[matcher.scala 68:17]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[matcher.scala 68:17]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[matcher.scala 68:17]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[matcher.scala 68:17]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[matcher.scala 68:17]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[matcher.scala 68:17]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[matcher.scala 68:17]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[matcher.scala 68:17]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[matcher.scala 68:17]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[matcher.scala 68:17]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[matcher.scala 68:17]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[matcher.scala 68:17]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[matcher.scala 68:17]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[matcher.scala 68:17]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[matcher.scala 68:17]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[matcher.scala 68:17]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[matcher.scala 68:17]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[matcher.scala 68:17]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[matcher.scala 68:17]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[matcher.scala 68:17]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[matcher.scala 68:17]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[matcher.scala 68:17]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[matcher.scala 68:17]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[matcher.scala 68:17]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[matcher.scala 68:17]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[matcher.scala 68:17]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[matcher.scala 68:17]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[matcher.scala 68:17]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[matcher.scala 68:17]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[matcher.scala 68:17]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[matcher.scala 68:17]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[matcher.scala 68:17]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[matcher.scala 68:17]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[matcher.scala 68:17]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[matcher.scala 68:17]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[matcher.scala 68:17]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[matcher.scala 68:17]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[matcher.scala 68:17]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[matcher.scala 68:17]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[matcher.scala 68:17]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[matcher.scala 68:17]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[matcher.scala 68:17]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[matcher.scala 68:17]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[matcher.scala 68:17]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[matcher.scala 68:17]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[matcher.scala 68:17]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[matcher.scala 68:17]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[matcher.scala 68:17]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[matcher.scala 68:17]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[matcher.scala 68:17]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[matcher.scala 68:17]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[matcher.scala 68:17]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[matcher.scala 68:17]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[matcher.scala 68:17]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[matcher.scala 68:17]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[matcher.scala 68:17]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[matcher.scala 68:17]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[matcher.scala 68:17]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[matcher.scala 68:17]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[matcher.scala 68:17]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[matcher.scala 68:17]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[matcher.scala 68:17]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[matcher.scala 68:17]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[matcher.scala 68:17]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[matcher.scala 68:17]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[matcher.scala 68:17]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[matcher.scala 68:17]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[matcher.scala 68:17]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[matcher.scala 68:17]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[matcher.scala 68:17]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[matcher.scala 68:17]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[matcher.scala 68:17]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[matcher.scala 68:17]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[matcher.scala 68:17]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[matcher.scala 68:17]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[matcher.scala 68:17]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[matcher.scala 68:17]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[matcher.scala 68:17]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[matcher.scala 68:17]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[matcher.scala 68:17]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[matcher.scala 68:17]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[matcher.scala 68:17]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[matcher.scala 68:17]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[matcher.scala 68:17]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[matcher.scala 68:17]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[matcher.scala 68:17]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[matcher.scala 68:17]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[matcher.scala 68:17]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[matcher.scala 68:17]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[matcher.scala 68:17]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[matcher.scala 68:17]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[matcher.scala 68:17]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[matcher.scala 68:17]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[matcher.scala 68:17]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[matcher.scala 68:17]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[matcher.scala 68:17]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[matcher.scala 68:17]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[matcher.scala 68:17]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[matcher.scala 68:17]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[matcher.scala 68:17]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[matcher.scala 68:17]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[matcher.scala 68:17]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[matcher.scala 68:17]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[matcher.scala 68:17]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[matcher.scala 68:17]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[matcher.scala 68:17]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[matcher.scala 68:17]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[matcher.scala 68:17]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[matcher.scala 68:17]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[matcher.scala 68:17]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[matcher.scala 68:17]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[matcher.scala 68:17]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[matcher.scala 68:17]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[matcher.scala 68:17]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[matcher.scala 68:17]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[matcher.scala 68:17]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[matcher.scala 68:17]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[matcher.scala 68:17]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[matcher.scala 68:17]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[matcher.scala 68:17]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[matcher.scala 68:17]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[matcher.scala 68:17]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[matcher.scala 68:17]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[matcher.scala 68:17]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[matcher.scala 68:17]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[matcher.scala 68:17]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[matcher.scala 68:17]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[matcher.scala 68:17]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[matcher.scala 68:17]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[matcher.scala 68:17]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[matcher.scala 68:17]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[matcher.scala 68:17]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[matcher.scala 68:17]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[matcher.scala 68:17]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[matcher.scala 68:17]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[matcher.scala 68:17]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[matcher.scala 68:17]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[matcher.scala 68:17]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[matcher.scala 68:17]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[matcher.scala 68:17]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[matcher.scala 68:17]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[matcher.scala 68:17]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[matcher.scala 68:17]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[matcher.scala 68:17]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[matcher.scala 68:17]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[matcher.scala 68:17]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[matcher.scala 68:17]
    key_offset <= io_key_offset_in; // @[matcher.scala 72:24]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_header_0 = _RAND_160[15:0];
  _RAND_161 = {1{`RANDOM}};
  phv_header_1 = _RAND_161[15:0];
  _RAND_162 = {1{`RANDOM}};
  phv_header_2 = _RAND_162[15:0];
  _RAND_163 = {1{`RANDOM}};
  phv_header_3 = _RAND_163[15:0];
  _RAND_164 = {1{`RANDOM}};
  phv_header_4 = _RAND_164[15:0];
  _RAND_165 = {1{`RANDOM}};
  phv_header_5 = _RAND_165[15:0];
  _RAND_166 = {1{`RANDOM}};
  phv_header_6 = _RAND_166[15:0];
  _RAND_167 = {1{`RANDOM}};
  phv_header_7 = _RAND_167[15:0];
  _RAND_168 = {1{`RANDOM}};
  phv_header_8 = _RAND_168[15:0];
  _RAND_169 = {1{`RANDOM}};
  phv_header_9 = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  phv_header_10 = _RAND_170[15:0];
  _RAND_171 = {1{`RANDOM}};
  phv_header_11 = _RAND_171[15:0];
  _RAND_172 = {1{`RANDOM}};
  phv_header_12 = _RAND_172[15:0];
  _RAND_173 = {1{`RANDOM}};
  phv_header_13 = _RAND_173[15:0];
  _RAND_174 = {1{`RANDOM}};
  phv_header_14 = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  phv_header_15 = _RAND_175[15:0];
  _RAND_176 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_178[15:0];
  _RAND_179 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_179[3:0];
  _RAND_180 = {1{`RANDOM}};
  phv_next_config_id = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  key_offset = _RAND_182[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
