module PrimitiveGetSource(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [1:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [1:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input  [7:0]  io_args_in_0,
  input  [7:0]  io_args_in_1,
  input  [7:0]  io_args_in_2,
  input  [7:0]  io_args_in_3,
  input  [7:0]  io_args_in_4,
  input  [7:0]  io_args_in_5,
  input  [7:0]  io_args_in_6,
  input  [31:0] io_vliw_in_0,
  input  [31:0] io_vliw_in_1,
  input  [31:0] io_vliw_in_2,
  input  [31:0] io_vliw_in_3,
  input  [7:0]  io_offset_in_0,
  input  [7:0]  io_offset_in_1,
  input  [7:0]  io_offset_in_2,
  input  [7:0]  io_offset_in_3,
  input  [7:0]  io_length_in_0,
  input  [7:0]  io_length_in_1,
  input  [7:0]  io_length_in_2,
  input  [7:0]  io_length_in_3,
  output [31:0] io_vliw_out_0,
  output [31:0] io_vliw_out_1,
  output [31:0] io_vliw_out_2,
  output [31:0] io_vliw_out_3,
  output [63:0] io_field_out_0,
  output [63:0] io_field_out_1,
  output [63:0] io_field_out_2,
  output [63:0] io_field_out_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[executor.scala 128:22]
  reg [7:0] phv_data_1; // @[executor.scala 128:22]
  reg [7:0] phv_data_2; // @[executor.scala 128:22]
  reg [7:0] phv_data_3; // @[executor.scala 128:22]
  reg [7:0] phv_data_4; // @[executor.scala 128:22]
  reg [7:0] phv_data_5; // @[executor.scala 128:22]
  reg [7:0] phv_data_6; // @[executor.scala 128:22]
  reg [7:0] phv_data_7; // @[executor.scala 128:22]
  reg [7:0] phv_data_8; // @[executor.scala 128:22]
  reg [7:0] phv_data_9; // @[executor.scala 128:22]
  reg [7:0] phv_data_10; // @[executor.scala 128:22]
  reg [7:0] phv_data_11; // @[executor.scala 128:22]
  reg [7:0] phv_data_12; // @[executor.scala 128:22]
  reg [7:0] phv_data_13; // @[executor.scala 128:22]
  reg [7:0] phv_data_14; // @[executor.scala 128:22]
  reg [7:0] phv_data_15; // @[executor.scala 128:22]
  reg [7:0] phv_data_16; // @[executor.scala 128:22]
  reg [7:0] phv_data_17; // @[executor.scala 128:22]
  reg [7:0] phv_data_18; // @[executor.scala 128:22]
  reg [7:0] phv_data_19; // @[executor.scala 128:22]
  reg [7:0] phv_data_20; // @[executor.scala 128:22]
  reg [7:0] phv_data_21; // @[executor.scala 128:22]
  reg [7:0] phv_data_22; // @[executor.scala 128:22]
  reg [7:0] phv_data_23; // @[executor.scala 128:22]
  reg [7:0] phv_data_24; // @[executor.scala 128:22]
  reg [7:0] phv_data_25; // @[executor.scala 128:22]
  reg [7:0] phv_data_26; // @[executor.scala 128:22]
  reg [7:0] phv_data_27; // @[executor.scala 128:22]
  reg [7:0] phv_data_28; // @[executor.scala 128:22]
  reg [7:0] phv_data_29; // @[executor.scala 128:22]
  reg [7:0] phv_data_30; // @[executor.scala 128:22]
  reg [7:0] phv_data_31; // @[executor.scala 128:22]
  reg [7:0] phv_data_32; // @[executor.scala 128:22]
  reg [7:0] phv_data_33; // @[executor.scala 128:22]
  reg [7:0] phv_data_34; // @[executor.scala 128:22]
  reg [7:0] phv_data_35; // @[executor.scala 128:22]
  reg [7:0] phv_data_36; // @[executor.scala 128:22]
  reg [7:0] phv_data_37; // @[executor.scala 128:22]
  reg [7:0] phv_data_38; // @[executor.scala 128:22]
  reg [7:0] phv_data_39; // @[executor.scala 128:22]
  reg [7:0] phv_data_40; // @[executor.scala 128:22]
  reg [7:0] phv_data_41; // @[executor.scala 128:22]
  reg [7:0] phv_data_42; // @[executor.scala 128:22]
  reg [7:0] phv_data_43; // @[executor.scala 128:22]
  reg [7:0] phv_data_44; // @[executor.scala 128:22]
  reg [7:0] phv_data_45; // @[executor.scala 128:22]
  reg [7:0] phv_data_46; // @[executor.scala 128:22]
  reg [7:0] phv_data_47; // @[executor.scala 128:22]
  reg [7:0] phv_data_48; // @[executor.scala 128:22]
  reg [7:0] phv_data_49; // @[executor.scala 128:22]
  reg [7:0] phv_data_50; // @[executor.scala 128:22]
  reg [7:0] phv_data_51; // @[executor.scala 128:22]
  reg [7:0] phv_data_52; // @[executor.scala 128:22]
  reg [7:0] phv_data_53; // @[executor.scala 128:22]
  reg [7:0] phv_data_54; // @[executor.scala 128:22]
  reg [7:0] phv_data_55; // @[executor.scala 128:22]
  reg [7:0] phv_data_56; // @[executor.scala 128:22]
  reg [7:0] phv_data_57; // @[executor.scala 128:22]
  reg [7:0] phv_data_58; // @[executor.scala 128:22]
  reg [7:0] phv_data_59; // @[executor.scala 128:22]
  reg [7:0] phv_data_60; // @[executor.scala 128:22]
  reg [7:0] phv_data_61; // @[executor.scala 128:22]
  reg [7:0] phv_data_62; // @[executor.scala 128:22]
  reg [7:0] phv_data_63; // @[executor.scala 128:22]
  reg [7:0] phv_data_64; // @[executor.scala 128:22]
  reg [7:0] phv_data_65; // @[executor.scala 128:22]
  reg [7:0] phv_data_66; // @[executor.scala 128:22]
  reg [7:0] phv_data_67; // @[executor.scala 128:22]
  reg [7:0] phv_data_68; // @[executor.scala 128:22]
  reg [7:0] phv_data_69; // @[executor.scala 128:22]
  reg [7:0] phv_data_70; // @[executor.scala 128:22]
  reg [7:0] phv_data_71; // @[executor.scala 128:22]
  reg [7:0] phv_data_72; // @[executor.scala 128:22]
  reg [7:0] phv_data_73; // @[executor.scala 128:22]
  reg [7:0] phv_data_74; // @[executor.scala 128:22]
  reg [7:0] phv_data_75; // @[executor.scala 128:22]
  reg [7:0] phv_data_76; // @[executor.scala 128:22]
  reg [7:0] phv_data_77; // @[executor.scala 128:22]
  reg [7:0] phv_data_78; // @[executor.scala 128:22]
  reg [7:0] phv_data_79; // @[executor.scala 128:22]
  reg [7:0] phv_data_80; // @[executor.scala 128:22]
  reg [7:0] phv_data_81; // @[executor.scala 128:22]
  reg [7:0] phv_data_82; // @[executor.scala 128:22]
  reg [7:0] phv_data_83; // @[executor.scala 128:22]
  reg [7:0] phv_data_84; // @[executor.scala 128:22]
  reg [7:0] phv_data_85; // @[executor.scala 128:22]
  reg [7:0] phv_data_86; // @[executor.scala 128:22]
  reg [7:0] phv_data_87; // @[executor.scala 128:22]
  reg [7:0] phv_data_88; // @[executor.scala 128:22]
  reg [7:0] phv_data_89; // @[executor.scala 128:22]
  reg [7:0] phv_data_90; // @[executor.scala 128:22]
  reg [7:0] phv_data_91; // @[executor.scala 128:22]
  reg [7:0] phv_data_92; // @[executor.scala 128:22]
  reg [7:0] phv_data_93; // @[executor.scala 128:22]
  reg [7:0] phv_data_94; // @[executor.scala 128:22]
  reg [7:0] phv_data_95; // @[executor.scala 128:22]
  reg [15:0] phv_header_0; // @[executor.scala 128:22]
  reg [15:0] phv_header_1; // @[executor.scala 128:22]
  reg [15:0] phv_header_2; // @[executor.scala 128:22]
  reg [15:0] phv_header_3; // @[executor.scala 128:22]
  reg [15:0] phv_header_4; // @[executor.scala 128:22]
  reg [15:0] phv_header_5; // @[executor.scala 128:22]
  reg [15:0] phv_header_6; // @[executor.scala 128:22]
  reg [15:0] phv_header_7; // @[executor.scala 128:22]
  reg [15:0] phv_header_8; // @[executor.scala 128:22]
  reg [15:0] phv_header_9; // @[executor.scala 128:22]
  reg [15:0] phv_header_10; // @[executor.scala 128:22]
  reg [15:0] phv_header_11; // @[executor.scala 128:22]
  reg [15:0] phv_header_12; // @[executor.scala 128:22]
  reg [15:0] phv_header_13; // @[executor.scala 128:22]
  reg [15:0] phv_header_14; // @[executor.scala 128:22]
  reg [15:0] phv_header_15; // @[executor.scala 128:22]
  reg [7:0] phv_parse_current_state; // @[executor.scala 128:22]
  reg [7:0] phv_parse_current_offset; // @[executor.scala 128:22]
  reg [15:0] phv_parse_transition_field; // @[executor.scala 128:22]
  reg [1:0] phv_next_processor_id; // @[executor.scala 128:22]
  reg  phv_next_config_id; // @[executor.scala 128:22]
  reg  phv_is_valid_processor; // @[executor.scala 128:22]
  reg [7:0] args_0; // @[executor.scala 132:23]
  reg [7:0] args_1; // @[executor.scala 132:23]
  reg [7:0] args_2; // @[executor.scala 132:23]
  reg [7:0] args_3; // @[executor.scala 132:23]
  reg [7:0] args_4; // @[executor.scala 132:23]
  reg [7:0] args_5; // @[executor.scala 132:23]
  reg [7:0] args_6; // @[executor.scala 132:23]
  reg [31:0] vliw_0; // @[executor.scala 135:23]
  reg [31:0] vliw_1; // @[executor.scala 135:23]
  reg [31:0] vliw_2; // @[executor.scala 135:23]
  reg [31:0] vliw_3; // @[executor.scala 135:23]
  reg [7:0] offset_0; // @[executor.scala 139:25]
  reg [7:0] offset_1; // @[executor.scala 139:25]
  reg [7:0] offset_2; // @[executor.scala 139:25]
  reg [7:0] offset_3; // @[executor.scala 139:25]
  reg [7:0] length_0; // @[executor.scala 140:25]
  reg [7:0] length_1; // @[executor.scala 140:25]
  reg [7:0] length_2; // @[executor.scala 140:25]
  reg [7:0] length_3; // @[executor.scala 140:25]
  wire [3:0] opcode = vliw_0[31:28]; // @[primitive.scala 9:44]
  wire [13:0] io_field_out_0_lo = vliw_0[13:0]; // @[primitive.scala 11:44]
  wire  from_header = length_0 != 8'h0; // @[executor.scala 151:45]
  wire [8:0] _total_offset_T = {{1'd0}, offset_0}; // @[executor.scala 158:57]
  wire [7:0] total_offset = _total_offset_T[7:0]; // @[executor.scala 158:57]
  wire [7:0] _GEN_1 = 7'h1 == total_offset[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2 = 7'h2 == total_offset[6:0] ? phv_data_2 : _GEN_1; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3 = 7'h3 == total_offset[6:0] ? phv_data_3 : _GEN_2; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_4 = 7'h4 == total_offset[6:0] ? phv_data_4 : _GEN_3; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_5 = 7'h5 == total_offset[6:0] ? phv_data_5 : _GEN_4; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_6 = 7'h6 == total_offset[6:0] ? phv_data_6 : _GEN_5; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_7 = 7'h7 == total_offset[6:0] ? phv_data_7 : _GEN_6; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_8 = 7'h8 == total_offset[6:0] ? phv_data_8 : _GEN_7; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_9 = 7'h9 == total_offset[6:0] ? phv_data_9 : _GEN_8; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_10 = 7'ha == total_offset[6:0] ? phv_data_10 : _GEN_9; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_11 = 7'hb == total_offset[6:0] ? phv_data_11 : _GEN_10; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_12 = 7'hc == total_offset[6:0] ? phv_data_12 : _GEN_11; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_13 = 7'hd == total_offset[6:0] ? phv_data_13 : _GEN_12; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_14 = 7'he == total_offset[6:0] ? phv_data_14 : _GEN_13; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_15 = 7'hf == total_offset[6:0] ? phv_data_15 : _GEN_14; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_16 = 7'h10 == total_offset[6:0] ? phv_data_16 : _GEN_15; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_17 = 7'h11 == total_offset[6:0] ? phv_data_17 : _GEN_16; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_18 = 7'h12 == total_offset[6:0] ? phv_data_18 : _GEN_17; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_19 = 7'h13 == total_offset[6:0] ? phv_data_19 : _GEN_18; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_20 = 7'h14 == total_offset[6:0] ? phv_data_20 : _GEN_19; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_21 = 7'h15 == total_offset[6:0] ? phv_data_21 : _GEN_20; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_22 = 7'h16 == total_offset[6:0] ? phv_data_22 : _GEN_21; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_23 = 7'h17 == total_offset[6:0] ? phv_data_23 : _GEN_22; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_24 = 7'h18 == total_offset[6:0] ? phv_data_24 : _GEN_23; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_25 = 7'h19 == total_offset[6:0] ? phv_data_25 : _GEN_24; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_26 = 7'h1a == total_offset[6:0] ? phv_data_26 : _GEN_25; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_27 = 7'h1b == total_offset[6:0] ? phv_data_27 : _GEN_26; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_28 = 7'h1c == total_offset[6:0] ? phv_data_28 : _GEN_27; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_29 = 7'h1d == total_offset[6:0] ? phv_data_29 : _GEN_28; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_30 = 7'h1e == total_offset[6:0] ? phv_data_30 : _GEN_29; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_31 = 7'h1f == total_offset[6:0] ? phv_data_31 : _GEN_30; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_32 = 7'h20 == total_offset[6:0] ? phv_data_32 : _GEN_31; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_33 = 7'h21 == total_offset[6:0] ? phv_data_33 : _GEN_32; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_34 = 7'h22 == total_offset[6:0] ? phv_data_34 : _GEN_33; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_35 = 7'h23 == total_offset[6:0] ? phv_data_35 : _GEN_34; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_36 = 7'h24 == total_offset[6:0] ? phv_data_36 : _GEN_35; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_37 = 7'h25 == total_offset[6:0] ? phv_data_37 : _GEN_36; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_38 = 7'h26 == total_offset[6:0] ? phv_data_38 : _GEN_37; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_39 = 7'h27 == total_offset[6:0] ? phv_data_39 : _GEN_38; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_40 = 7'h28 == total_offset[6:0] ? phv_data_40 : _GEN_39; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_41 = 7'h29 == total_offset[6:0] ? phv_data_41 : _GEN_40; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_42 = 7'h2a == total_offset[6:0] ? phv_data_42 : _GEN_41; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_43 = 7'h2b == total_offset[6:0] ? phv_data_43 : _GEN_42; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_44 = 7'h2c == total_offset[6:0] ? phv_data_44 : _GEN_43; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_45 = 7'h2d == total_offset[6:0] ? phv_data_45 : _GEN_44; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_46 = 7'h2e == total_offset[6:0] ? phv_data_46 : _GEN_45; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_47 = 7'h2f == total_offset[6:0] ? phv_data_47 : _GEN_46; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_48 = 7'h30 == total_offset[6:0] ? phv_data_48 : _GEN_47; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_49 = 7'h31 == total_offset[6:0] ? phv_data_49 : _GEN_48; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_50 = 7'h32 == total_offset[6:0] ? phv_data_50 : _GEN_49; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_51 = 7'h33 == total_offset[6:0] ? phv_data_51 : _GEN_50; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_52 = 7'h34 == total_offset[6:0] ? phv_data_52 : _GEN_51; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_53 = 7'h35 == total_offset[6:0] ? phv_data_53 : _GEN_52; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_54 = 7'h36 == total_offset[6:0] ? phv_data_54 : _GEN_53; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_55 = 7'h37 == total_offset[6:0] ? phv_data_55 : _GEN_54; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_56 = 7'h38 == total_offset[6:0] ? phv_data_56 : _GEN_55; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_57 = 7'h39 == total_offset[6:0] ? phv_data_57 : _GEN_56; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_58 = 7'h3a == total_offset[6:0] ? phv_data_58 : _GEN_57; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_59 = 7'h3b == total_offset[6:0] ? phv_data_59 : _GEN_58; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_60 = 7'h3c == total_offset[6:0] ? phv_data_60 : _GEN_59; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_61 = 7'h3d == total_offset[6:0] ? phv_data_61 : _GEN_60; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_62 = 7'h3e == total_offset[6:0] ? phv_data_62 : _GEN_61; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_63 = 7'h3f == total_offset[6:0] ? phv_data_63 : _GEN_62; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_64 = 7'h40 == total_offset[6:0] ? phv_data_64 : _GEN_63; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_65 = 7'h41 == total_offset[6:0] ? phv_data_65 : _GEN_64; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_66 = 7'h42 == total_offset[6:0] ? phv_data_66 : _GEN_65; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_67 = 7'h43 == total_offset[6:0] ? phv_data_67 : _GEN_66; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_68 = 7'h44 == total_offset[6:0] ? phv_data_68 : _GEN_67; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_69 = 7'h45 == total_offset[6:0] ? phv_data_69 : _GEN_68; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_70 = 7'h46 == total_offset[6:0] ? phv_data_70 : _GEN_69; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_71 = 7'h47 == total_offset[6:0] ? phv_data_71 : _GEN_70; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_72 = 7'h48 == total_offset[6:0] ? phv_data_72 : _GEN_71; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_73 = 7'h49 == total_offset[6:0] ? phv_data_73 : _GEN_72; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_74 = 7'h4a == total_offset[6:0] ? phv_data_74 : _GEN_73; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_75 = 7'h4b == total_offset[6:0] ? phv_data_75 : _GEN_74; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_76 = 7'h4c == total_offset[6:0] ? phv_data_76 : _GEN_75; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_77 = 7'h4d == total_offset[6:0] ? phv_data_77 : _GEN_76; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_78 = 7'h4e == total_offset[6:0] ? phv_data_78 : _GEN_77; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_79 = 7'h4f == total_offset[6:0] ? phv_data_79 : _GEN_78; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_80 = 7'h50 == total_offset[6:0] ? phv_data_80 : _GEN_79; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_81 = 7'h51 == total_offset[6:0] ? phv_data_81 : _GEN_80; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_82 = 7'h52 == total_offset[6:0] ? phv_data_82 : _GEN_81; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_83 = 7'h53 == total_offset[6:0] ? phv_data_83 : _GEN_82; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_84 = 7'h54 == total_offset[6:0] ? phv_data_84 : _GEN_83; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_85 = 7'h55 == total_offset[6:0] ? phv_data_85 : _GEN_84; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_86 = 7'h56 == total_offset[6:0] ? phv_data_86 : _GEN_85; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_87 = 7'h57 == total_offset[6:0] ? phv_data_87 : _GEN_86; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_88 = 7'h58 == total_offset[6:0] ? phv_data_88 : _GEN_87; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_89 = 7'h59 == total_offset[6:0] ? phv_data_89 : _GEN_88; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_90 = 7'h5a == total_offset[6:0] ? phv_data_90 : _GEN_89; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_91 = 7'h5b == total_offset[6:0] ? phv_data_91 : _GEN_90; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_92 = 7'h5c == total_offset[6:0] ? phv_data_92 : _GEN_91; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_93 = 7'h5d == total_offset[6:0] ? phv_data_93 : _GEN_92; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_94 = 7'h5e == total_offset[6:0] ? phv_data_94 : _GEN_93; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_95 = 7'h5f == total_offset[6:0] ? phv_data_95 : _GEN_94; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes__0 = 8'h0 < length_0 ? _GEN_95 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_1 = offset_0 + 8'h1; // @[executor.scala 158:57]
  wire [7:0] _GEN_98 = 7'h1 == total_offset_1[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_99 = 7'h2 == total_offset_1[6:0] ? phv_data_2 : _GEN_98; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_100 = 7'h3 == total_offset_1[6:0] ? phv_data_3 : _GEN_99; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_101 = 7'h4 == total_offset_1[6:0] ? phv_data_4 : _GEN_100; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_102 = 7'h5 == total_offset_1[6:0] ? phv_data_5 : _GEN_101; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_103 = 7'h6 == total_offset_1[6:0] ? phv_data_6 : _GEN_102; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_104 = 7'h7 == total_offset_1[6:0] ? phv_data_7 : _GEN_103; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_105 = 7'h8 == total_offset_1[6:0] ? phv_data_8 : _GEN_104; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_106 = 7'h9 == total_offset_1[6:0] ? phv_data_9 : _GEN_105; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_107 = 7'ha == total_offset_1[6:0] ? phv_data_10 : _GEN_106; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_108 = 7'hb == total_offset_1[6:0] ? phv_data_11 : _GEN_107; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_109 = 7'hc == total_offset_1[6:0] ? phv_data_12 : _GEN_108; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_110 = 7'hd == total_offset_1[6:0] ? phv_data_13 : _GEN_109; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_111 = 7'he == total_offset_1[6:0] ? phv_data_14 : _GEN_110; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_112 = 7'hf == total_offset_1[6:0] ? phv_data_15 : _GEN_111; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_113 = 7'h10 == total_offset_1[6:0] ? phv_data_16 : _GEN_112; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_114 = 7'h11 == total_offset_1[6:0] ? phv_data_17 : _GEN_113; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_115 = 7'h12 == total_offset_1[6:0] ? phv_data_18 : _GEN_114; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_116 = 7'h13 == total_offset_1[6:0] ? phv_data_19 : _GEN_115; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_117 = 7'h14 == total_offset_1[6:0] ? phv_data_20 : _GEN_116; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_118 = 7'h15 == total_offset_1[6:0] ? phv_data_21 : _GEN_117; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_119 = 7'h16 == total_offset_1[6:0] ? phv_data_22 : _GEN_118; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_120 = 7'h17 == total_offset_1[6:0] ? phv_data_23 : _GEN_119; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_121 = 7'h18 == total_offset_1[6:0] ? phv_data_24 : _GEN_120; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_122 = 7'h19 == total_offset_1[6:0] ? phv_data_25 : _GEN_121; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_123 = 7'h1a == total_offset_1[6:0] ? phv_data_26 : _GEN_122; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_124 = 7'h1b == total_offset_1[6:0] ? phv_data_27 : _GEN_123; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_125 = 7'h1c == total_offset_1[6:0] ? phv_data_28 : _GEN_124; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_126 = 7'h1d == total_offset_1[6:0] ? phv_data_29 : _GEN_125; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_127 = 7'h1e == total_offset_1[6:0] ? phv_data_30 : _GEN_126; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_128 = 7'h1f == total_offset_1[6:0] ? phv_data_31 : _GEN_127; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_129 = 7'h20 == total_offset_1[6:0] ? phv_data_32 : _GEN_128; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_130 = 7'h21 == total_offset_1[6:0] ? phv_data_33 : _GEN_129; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_131 = 7'h22 == total_offset_1[6:0] ? phv_data_34 : _GEN_130; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_132 = 7'h23 == total_offset_1[6:0] ? phv_data_35 : _GEN_131; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_133 = 7'h24 == total_offset_1[6:0] ? phv_data_36 : _GEN_132; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_134 = 7'h25 == total_offset_1[6:0] ? phv_data_37 : _GEN_133; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_135 = 7'h26 == total_offset_1[6:0] ? phv_data_38 : _GEN_134; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_136 = 7'h27 == total_offset_1[6:0] ? phv_data_39 : _GEN_135; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_137 = 7'h28 == total_offset_1[6:0] ? phv_data_40 : _GEN_136; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_138 = 7'h29 == total_offset_1[6:0] ? phv_data_41 : _GEN_137; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_139 = 7'h2a == total_offset_1[6:0] ? phv_data_42 : _GEN_138; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_140 = 7'h2b == total_offset_1[6:0] ? phv_data_43 : _GEN_139; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_141 = 7'h2c == total_offset_1[6:0] ? phv_data_44 : _GEN_140; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_142 = 7'h2d == total_offset_1[6:0] ? phv_data_45 : _GEN_141; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_143 = 7'h2e == total_offset_1[6:0] ? phv_data_46 : _GEN_142; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_144 = 7'h2f == total_offset_1[6:0] ? phv_data_47 : _GEN_143; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_145 = 7'h30 == total_offset_1[6:0] ? phv_data_48 : _GEN_144; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_146 = 7'h31 == total_offset_1[6:0] ? phv_data_49 : _GEN_145; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_147 = 7'h32 == total_offset_1[6:0] ? phv_data_50 : _GEN_146; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_148 = 7'h33 == total_offset_1[6:0] ? phv_data_51 : _GEN_147; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_149 = 7'h34 == total_offset_1[6:0] ? phv_data_52 : _GEN_148; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_150 = 7'h35 == total_offset_1[6:0] ? phv_data_53 : _GEN_149; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_151 = 7'h36 == total_offset_1[6:0] ? phv_data_54 : _GEN_150; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_152 = 7'h37 == total_offset_1[6:0] ? phv_data_55 : _GEN_151; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_153 = 7'h38 == total_offset_1[6:0] ? phv_data_56 : _GEN_152; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_154 = 7'h39 == total_offset_1[6:0] ? phv_data_57 : _GEN_153; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_155 = 7'h3a == total_offset_1[6:0] ? phv_data_58 : _GEN_154; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_156 = 7'h3b == total_offset_1[6:0] ? phv_data_59 : _GEN_155; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_157 = 7'h3c == total_offset_1[6:0] ? phv_data_60 : _GEN_156; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_158 = 7'h3d == total_offset_1[6:0] ? phv_data_61 : _GEN_157; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_159 = 7'h3e == total_offset_1[6:0] ? phv_data_62 : _GEN_158; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_160 = 7'h3f == total_offset_1[6:0] ? phv_data_63 : _GEN_159; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_161 = 7'h40 == total_offset_1[6:0] ? phv_data_64 : _GEN_160; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_162 = 7'h41 == total_offset_1[6:0] ? phv_data_65 : _GEN_161; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_163 = 7'h42 == total_offset_1[6:0] ? phv_data_66 : _GEN_162; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_164 = 7'h43 == total_offset_1[6:0] ? phv_data_67 : _GEN_163; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_165 = 7'h44 == total_offset_1[6:0] ? phv_data_68 : _GEN_164; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_166 = 7'h45 == total_offset_1[6:0] ? phv_data_69 : _GEN_165; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_167 = 7'h46 == total_offset_1[6:0] ? phv_data_70 : _GEN_166; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_168 = 7'h47 == total_offset_1[6:0] ? phv_data_71 : _GEN_167; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_169 = 7'h48 == total_offset_1[6:0] ? phv_data_72 : _GEN_168; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_170 = 7'h49 == total_offset_1[6:0] ? phv_data_73 : _GEN_169; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_171 = 7'h4a == total_offset_1[6:0] ? phv_data_74 : _GEN_170; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_172 = 7'h4b == total_offset_1[6:0] ? phv_data_75 : _GEN_171; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_173 = 7'h4c == total_offset_1[6:0] ? phv_data_76 : _GEN_172; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_174 = 7'h4d == total_offset_1[6:0] ? phv_data_77 : _GEN_173; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_175 = 7'h4e == total_offset_1[6:0] ? phv_data_78 : _GEN_174; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_176 = 7'h4f == total_offset_1[6:0] ? phv_data_79 : _GEN_175; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_177 = 7'h50 == total_offset_1[6:0] ? phv_data_80 : _GEN_176; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_178 = 7'h51 == total_offset_1[6:0] ? phv_data_81 : _GEN_177; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_179 = 7'h52 == total_offset_1[6:0] ? phv_data_82 : _GEN_178; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_180 = 7'h53 == total_offset_1[6:0] ? phv_data_83 : _GEN_179; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_181 = 7'h54 == total_offset_1[6:0] ? phv_data_84 : _GEN_180; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_182 = 7'h55 == total_offset_1[6:0] ? phv_data_85 : _GEN_181; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_183 = 7'h56 == total_offset_1[6:0] ? phv_data_86 : _GEN_182; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_184 = 7'h57 == total_offset_1[6:0] ? phv_data_87 : _GEN_183; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_185 = 7'h58 == total_offset_1[6:0] ? phv_data_88 : _GEN_184; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_186 = 7'h59 == total_offset_1[6:0] ? phv_data_89 : _GEN_185; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_187 = 7'h5a == total_offset_1[6:0] ? phv_data_90 : _GEN_186; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_188 = 7'h5b == total_offset_1[6:0] ? phv_data_91 : _GEN_187; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_189 = 7'h5c == total_offset_1[6:0] ? phv_data_92 : _GEN_188; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_190 = 7'h5d == total_offset_1[6:0] ? phv_data_93 : _GEN_189; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_191 = 7'h5e == total_offset_1[6:0] ? phv_data_94 : _GEN_190; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_192 = 7'h5f == total_offset_1[6:0] ? phv_data_95 : _GEN_191; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes__1 = 8'h1 < length_0 ? _GEN_192 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_2 = offset_0 + 8'h2; // @[executor.scala 158:57]
  wire [7:0] _GEN_195 = 7'h1 == total_offset_2[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_196 = 7'h2 == total_offset_2[6:0] ? phv_data_2 : _GEN_195; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_197 = 7'h3 == total_offset_2[6:0] ? phv_data_3 : _GEN_196; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_198 = 7'h4 == total_offset_2[6:0] ? phv_data_4 : _GEN_197; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_199 = 7'h5 == total_offset_2[6:0] ? phv_data_5 : _GEN_198; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_200 = 7'h6 == total_offset_2[6:0] ? phv_data_6 : _GEN_199; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_201 = 7'h7 == total_offset_2[6:0] ? phv_data_7 : _GEN_200; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_202 = 7'h8 == total_offset_2[6:0] ? phv_data_8 : _GEN_201; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_203 = 7'h9 == total_offset_2[6:0] ? phv_data_9 : _GEN_202; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_204 = 7'ha == total_offset_2[6:0] ? phv_data_10 : _GEN_203; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_205 = 7'hb == total_offset_2[6:0] ? phv_data_11 : _GEN_204; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_206 = 7'hc == total_offset_2[6:0] ? phv_data_12 : _GEN_205; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_207 = 7'hd == total_offset_2[6:0] ? phv_data_13 : _GEN_206; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_208 = 7'he == total_offset_2[6:0] ? phv_data_14 : _GEN_207; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_209 = 7'hf == total_offset_2[6:0] ? phv_data_15 : _GEN_208; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_210 = 7'h10 == total_offset_2[6:0] ? phv_data_16 : _GEN_209; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_211 = 7'h11 == total_offset_2[6:0] ? phv_data_17 : _GEN_210; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_212 = 7'h12 == total_offset_2[6:0] ? phv_data_18 : _GEN_211; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_213 = 7'h13 == total_offset_2[6:0] ? phv_data_19 : _GEN_212; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_214 = 7'h14 == total_offset_2[6:0] ? phv_data_20 : _GEN_213; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_215 = 7'h15 == total_offset_2[6:0] ? phv_data_21 : _GEN_214; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_216 = 7'h16 == total_offset_2[6:0] ? phv_data_22 : _GEN_215; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_217 = 7'h17 == total_offset_2[6:0] ? phv_data_23 : _GEN_216; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_218 = 7'h18 == total_offset_2[6:0] ? phv_data_24 : _GEN_217; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_219 = 7'h19 == total_offset_2[6:0] ? phv_data_25 : _GEN_218; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_220 = 7'h1a == total_offset_2[6:0] ? phv_data_26 : _GEN_219; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_221 = 7'h1b == total_offset_2[6:0] ? phv_data_27 : _GEN_220; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_222 = 7'h1c == total_offset_2[6:0] ? phv_data_28 : _GEN_221; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_223 = 7'h1d == total_offset_2[6:0] ? phv_data_29 : _GEN_222; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_224 = 7'h1e == total_offset_2[6:0] ? phv_data_30 : _GEN_223; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_225 = 7'h1f == total_offset_2[6:0] ? phv_data_31 : _GEN_224; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_226 = 7'h20 == total_offset_2[6:0] ? phv_data_32 : _GEN_225; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_227 = 7'h21 == total_offset_2[6:0] ? phv_data_33 : _GEN_226; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_228 = 7'h22 == total_offset_2[6:0] ? phv_data_34 : _GEN_227; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_229 = 7'h23 == total_offset_2[6:0] ? phv_data_35 : _GEN_228; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_230 = 7'h24 == total_offset_2[6:0] ? phv_data_36 : _GEN_229; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_231 = 7'h25 == total_offset_2[6:0] ? phv_data_37 : _GEN_230; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_232 = 7'h26 == total_offset_2[6:0] ? phv_data_38 : _GEN_231; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_233 = 7'h27 == total_offset_2[6:0] ? phv_data_39 : _GEN_232; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_234 = 7'h28 == total_offset_2[6:0] ? phv_data_40 : _GEN_233; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_235 = 7'h29 == total_offset_2[6:0] ? phv_data_41 : _GEN_234; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_236 = 7'h2a == total_offset_2[6:0] ? phv_data_42 : _GEN_235; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_237 = 7'h2b == total_offset_2[6:0] ? phv_data_43 : _GEN_236; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_238 = 7'h2c == total_offset_2[6:0] ? phv_data_44 : _GEN_237; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_239 = 7'h2d == total_offset_2[6:0] ? phv_data_45 : _GEN_238; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_240 = 7'h2e == total_offset_2[6:0] ? phv_data_46 : _GEN_239; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_241 = 7'h2f == total_offset_2[6:0] ? phv_data_47 : _GEN_240; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_242 = 7'h30 == total_offset_2[6:0] ? phv_data_48 : _GEN_241; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_243 = 7'h31 == total_offset_2[6:0] ? phv_data_49 : _GEN_242; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_244 = 7'h32 == total_offset_2[6:0] ? phv_data_50 : _GEN_243; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_245 = 7'h33 == total_offset_2[6:0] ? phv_data_51 : _GEN_244; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_246 = 7'h34 == total_offset_2[6:0] ? phv_data_52 : _GEN_245; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_247 = 7'h35 == total_offset_2[6:0] ? phv_data_53 : _GEN_246; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_248 = 7'h36 == total_offset_2[6:0] ? phv_data_54 : _GEN_247; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_249 = 7'h37 == total_offset_2[6:0] ? phv_data_55 : _GEN_248; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_250 = 7'h38 == total_offset_2[6:0] ? phv_data_56 : _GEN_249; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_251 = 7'h39 == total_offset_2[6:0] ? phv_data_57 : _GEN_250; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_252 = 7'h3a == total_offset_2[6:0] ? phv_data_58 : _GEN_251; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_253 = 7'h3b == total_offset_2[6:0] ? phv_data_59 : _GEN_252; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_254 = 7'h3c == total_offset_2[6:0] ? phv_data_60 : _GEN_253; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_255 = 7'h3d == total_offset_2[6:0] ? phv_data_61 : _GEN_254; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_256 = 7'h3e == total_offset_2[6:0] ? phv_data_62 : _GEN_255; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_257 = 7'h3f == total_offset_2[6:0] ? phv_data_63 : _GEN_256; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_258 = 7'h40 == total_offset_2[6:0] ? phv_data_64 : _GEN_257; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_259 = 7'h41 == total_offset_2[6:0] ? phv_data_65 : _GEN_258; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_260 = 7'h42 == total_offset_2[6:0] ? phv_data_66 : _GEN_259; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_261 = 7'h43 == total_offset_2[6:0] ? phv_data_67 : _GEN_260; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_262 = 7'h44 == total_offset_2[6:0] ? phv_data_68 : _GEN_261; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_263 = 7'h45 == total_offset_2[6:0] ? phv_data_69 : _GEN_262; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_264 = 7'h46 == total_offset_2[6:0] ? phv_data_70 : _GEN_263; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_265 = 7'h47 == total_offset_2[6:0] ? phv_data_71 : _GEN_264; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_266 = 7'h48 == total_offset_2[6:0] ? phv_data_72 : _GEN_265; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_267 = 7'h49 == total_offset_2[6:0] ? phv_data_73 : _GEN_266; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_268 = 7'h4a == total_offset_2[6:0] ? phv_data_74 : _GEN_267; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_269 = 7'h4b == total_offset_2[6:0] ? phv_data_75 : _GEN_268; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_270 = 7'h4c == total_offset_2[6:0] ? phv_data_76 : _GEN_269; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_271 = 7'h4d == total_offset_2[6:0] ? phv_data_77 : _GEN_270; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_272 = 7'h4e == total_offset_2[6:0] ? phv_data_78 : _GEN_271; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_273 = 7'h4f == total_offset_2[6:0] ? phv_data_79 : _GEN_272; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_274 = 7'h50 == total_offset_2[6:0] ? phv_data_80 : _GEN_273; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_275 = 7'h51 == total_offset_2[6:0] ? phv_data_81 : _GEN_274; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_276 = 7'h52 == total_offset_2[6:0] ? phv_data_82 : _GEN_275; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_277 = 7'h53 == total_offset_2[6:0] ? phv_data_83 : _GEN_276; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_278 = 7'h54 == total_offset_2[6:0] ? phv_data_84 : _GEN_277; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_279 = 7'h55 == total_offset_2[6:0] ? phv_data_85 : _GEN_278; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_280 = 7'h56 == total_offset_2[6:0] ? phv_data_86 : _GEN_279; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_281 = 7'h57 == total_offset_2[6:0] ? phv_data_87 : _GEN_280; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_282 = 7'h58 == total_offset_2[6:0] ? phv_data_88 : _GEN_281; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_283 = 7'h59 == total_offset_2[6:0] ? phv_data_89 : _GEN_282; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_284 = 7'h5a == total_offset_2[6:0] ? phv_data_90 : _GEN_283; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_285 = 7'h5b == total_offset_2[6:0] ? phv_data_91 : _GEN_284; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_286 = 7'h5c == total_offset_2[6:0] ? phv_data_92 : _GEN_285; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_287 = 7'h5d == total_offset_2[6:0] ? phv_data_93 : _GEN_286; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_288 = 7'h5e == total_offset_2[6:0] ? phv_data_94 : _GEN_287; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_289 = 7'h5f == total_offset_2[6:0] ? phv_data_95 : _GEN_288; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes__2 = 8'h2 < length_0 ? _GEN_289 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_3 = offset_0 + 8'h3; // @[executor.scala 158:57]
  wire [7:0] _GEN_292 = 7'h1 == total_offset_3[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_293 = 7'h2 == total_offset_3[6:0] ? phv_data_2 : _GEN_292; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_294 = 7'h3 == total_offset_3[6:0] ? phv_data_3 : _GEN_293; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_295 = 7'h4 == total_offset_3[6:0] ? phv_data_4 : _GEN_294; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_296 = 7'h5 == total_offset_3[6:0] ? phv_data_5 : _GEN_295; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_297 = 7'h6 == total_offset_3[6:0] ? phv_data_6 : _GEN_296; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_298 = 7'h7 == total_offset_3[6:0] ? phv_data_7 : _GEN_297; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_299 = 7'h8 == total_offset_3[6:0] ? phv_data_8 : _GEN_298; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_300 = 7'h9 == total_offset_3[6:0] ? phv_data_9 : _GEN_299; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_301 = 7'ha == total_offset_3[6:0] ? phv_data_10 : _GEN_300; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_302 = 7'hb == total_offset_3[6:0] ? phv_data_11 : _GEN_301; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_303 = 7'hc == total_offset_3[6:0] ? phv_data_12 : _GEN_302; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_304 = 7'hd == total_offset_3[6:0] ? phv_data_13 : _GEN_303; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_305 = 7'he == total_offset_3[6:0] ? phv_data_14 : _GEN_304; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_306 = 7'hf == total_offset_3[6:0] ? phv_data_15 : _GEN_305; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_307 = 7'h10 == total_offset_3[6:0] ? phv_data_16 : _GEN_306; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_308 = 7'h11 == total_offset_3[6:0] ? phv_data_17 : _GEN_307; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_309 = 7'h12 == total_offset_3[6:0] ? phv_data_18 : _GEN_308; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_310 = 7'h13 == total_offset_3[6:0] ? phv_data_19 : _GEN_309; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_311 = 7'h14 == total_offset_3[6:0] ? phv_data_20 : _GEN_310; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_312 = 7'h15 == total_offset_3[6:0] ? phv_data_21 : _GEN_311; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_313 = 7'h16 == total_offset_3[6:0] ? phv_data_22 : _GEN_312; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_314 = 7'h17 == total_offset_3[6:0] ? phv_data_23 : _GEN_313; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_315 = 7'h18 == total_offset_3[6:0] ? phv_data_24 : _GEN_314; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_316 = 7'h19 == total_offset_3[6:0] ? phv_data_25 : _GEN_315; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_317 = 7'h1a == total_offset_3[6:0] ? phv_data_26 : _GEN_316; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_318 = 7'h1b == total_offset_3[6:0] ? phv_data_27 : _GEN_317; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_319 = 7'h1c == total_offset_3[6:0] ? phv_data_28 : _GEN_318; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_320 = 7'h1d == total_offset_3[6:0] ? phv_data_29 : _GEN_319; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_321 = 7'h1e == total_offset_3[6:0] ? phv_data_30 : _GEN_320; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_322 = 7'h1f == total_offset_3[6:0] ? phv_data_31 : _GEN_321; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_323 = 7'h20 == total_offset_3[6:0] ? phv_data_32 : _GEN_322; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_324 = 7'h21 == total_offset_3[6:0] ? phv_data_33 : _GEN_323; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_325 = 7'h22 == total_offset_3[6:0] ? phv_data_34 : _GEN_324; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_326 = 7'h23 == total_offset_3[6:0] ? phv_data_35 : _GEN_325; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_327 = 7'h24 == total_offset_3[6:0] ? phv_data_36 : _GEN_326; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_328 = 7'h25 == total_offset_3[6:0] ? phv_data_37 : _GEN_327; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_329 = 7'h26 == total_offset_3[6:0] ? phv_data_38 : _GEN_328; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_330 = 7'h27 == total_offset_3[6:0] ? phv_data_39 : _GEN_329; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_331 = 7'h28 == total_offset_3[6:0] ? phv_data_40 : _GEN_330; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_332 = 7'h29 == total_offset_3[6:0] ? phv_data_41 : _GEN_331; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_333 = 7'h2a == total_offset_3[6:0] ? phv_data_42 : _GEN_332; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_334 = 7'h2b == total_offset_3[6:0] ? phv_data_43 : _GEN_333; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_335 = 7'h2c == total_offset_3[6:0] ? phv_data_44 : _GEN_334; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_336 = 7'h2d == total_offset_3[6:0] ? phv_data_45 : _GEN_335; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_337 = 7'h2e == total_offset_3[6:0] ? phv_data_46 : _GEN_336; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_338 = 7'h2f == total_offset_3[6:0] ? phv_data_47 : _GEN_337; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_339 = 7'h30 == total_offset_3[6:0] ? phv_data_48 : _GEN_338; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_340 = 7'h31 == total_offset_3[6:0] ? phv_data_49 : _GEN_339; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_341 = 7'h32 == total_offset_3[6:0] ? phv_data_50 : _GEN_340; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_342 = 7'h33 == total_offset_3[6:0] ? phv_data_51 : _GEN_341; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_343 = 7'h34 == total_offset_3[6:0] ? phv_data_52 : _GEN_342; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_344 = 7'h35 == total_offset_3[6:0] ? phv_data_53 : _GEN_343; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_345 = 7'h36 == total_offset_3[6:0] ? phv_data_54 : _GEN_344; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_346 = 7'h37 == total_offset_3[6:0] ? phv_data_55 : _GEN_345; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_347 = 7'h38 == total_offset_3[6:0] ? phv_data_56 : _GEN_346; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_348 = 7'h39 == total_offset_3[6:0] ? phv_data_57 : _GEN_347; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_349 = 7'h3a == total_offset_3[6:0] ? phv_data_58 : _GEN_348; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_350 = 7'h3b == total_offset_3[6:0] ? phv_data_59 : _GEN_349; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_351 = 7'h3c == total_offset_3[6:0] ? phv_data_60 : _GEN_350; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_352 = 7'h3d == total_offset_3[6:0] ? phv_data_61 : _GEN_351; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_353 = 7'h3e == total_offset_3[6:0] ? phv_data_62 : _GEN_352; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_354 = 7'h3f == total_offset_3[6:0] ? phv_data_63 : _GEN_353; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_355 = 7'h40 == total_offset_3[6:0] ? phv_data_64 : _GEN_354; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_356 = 7'h41 == total_offset_3[6:0] ? phv_data_65 : _GEN_355; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_357 = 7'h42 == total_offset_3[6:0] ? phv_data_66 : _GEN_356; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_358 = 7'h43 == total_offset_3[6:0] ? phv_data_67 : _GEN_357; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_359 = 7'h44 == total_offset_3[6:0] ? phv_data_68 : _GEN_358; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_360 = 7'h45 == total_offset_3[6:0] ? phv_data_69 : _GEN_359; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_361 = 7'h46 == total_offset_3[6:0] ? phv_data_70 : _GEN_360; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_362 = 7'h47 == total_offset_3[6:0] ? phv_data_71 : _GEN_361; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_363 = 7'h48 == total_offset_3[6:0] ? phv_data_72 : _GEN_362; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_364 = 7'h49 == total_offset_3[6:0] ? phv_data_73 : _GEN_363; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_365 = 7'h4a == total_offset_3[6:0] ? phv_data_74 : _GEN_364; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_366 = 7'h4b == total_offset_3[6:0] ? phv_data_75 : _GEN_365; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_367 = 7'h4c == total_offset_3[6:0] ? phv_data_76 : _GEN_366; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_368 = 7'h4d == total_offset_3[6:0] ? phv_data_77 : _GEN_367; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_369 = 7'h4e == total_offset_3[6:0] ? phv_data_78 : _GEN_368; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_370 = 7'h4f == total_offset_3[6:0] ? phv_data_79 : _GEN_369; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_371 = 7'h50 == total_offset_3[6:0] ? phv_data_80 : _GEN_370; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_372 = 7'h51 == total_offset_3[6:0] ? phv_data_81 : _GEN_371; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_373 = 7'h52 == total_offset_3[6:0] ? phv_data_82 : _GEN_372; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_374 = 7'h53 == total_offset_3[6:0] ? phv_data_83 : _GEN_373; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_375 = 7'h54 == total_offset_3[6:0] ? phv_data_84 : _GEN_374; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_376 = 7'h55 == total_offset_3[6:0] ? phv_data_85 : _GEN_375; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_377 = 7'h56 == total_offset_3[6:0] ? phv_data_86 : _GEN_376; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_378 = 7'h57 == total_offset_3[6:0] ? phv_data_87 : _GEN_377; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_379 = 7'h58 == total_offset_3[6:0] ? phv_data_88 : _GEN_378; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_380 = 7'h59 == total_offset_3[6:0] ? phv_data_89 : _GEN_379; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_381 = 7'h5a == total_offset_3[6:0] ? phv_data_90 : _GEN_380; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_382 = 7'h5b == total_offset_3[6:0] ? phv_data_91 : _GEN_381; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_383 = 7'h5c == total_offset_3[6:0] ? phv_data_92 : _GEN_382; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_384 = 7'h5d == total_offset_3[6:0] ? phv_data_93 : _GEN_383; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_385 = 7'h5e == total_offset_3[6:0] ? phv_data_94 : _GEN_384; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_386 = 7'h5f == total_offset_3[6:0] ? phv_data_95 : _GEN_385; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes__3 = 8'h3 < length_0 ? _GEN_386 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_4 = offset_0 + 8'h4; // @[executor.scala 158:57]
  wire [7:0] _GEN_389 = 7'h1 == total_offset_4[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_390 = 7'h2 == total_offset_4[6:0] ? phv_data_2 : _GEN_389; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_391 = 7'h3 == total_offset_4[6:0] ? phv_data_3 : _GEN_390; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_392 = 7'h4 == total_offset_4[6:0] ? phv_data_4 : _GEN_391; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_393 = 7'h5 == total_offset_4[6:0] ? phv_data_5 : _GEN_392; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_394 = 7'h6 == total_offset_4[6:0] ? phv_data_6 : _GEN_393; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_395 = 7'h7 == total_offset_4[6:0] ? phv_data_7 : _GEN_394; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_396 = 7'h8 == total_offset_4[6:0] ? phv_data_8 : _GEN_395; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_397 = 7'h9 == total_offset_4[6:0] ? phv_data_9 : _GEN_396; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_398 = 7'ha == total_offset_4[6:0] ? phv_data_10 : _GEN_397; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_399 = 7'hb == total_offset_4[6:0] ? phv_data_11 : _GEN_398; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_400 = 7'hc == total_offset_4[6:0] ? phv_data_12 : _GEN_399; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_401 = 7'hd == total_offset_4[6:0] ? phv_data_13 : _GEN_400; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_402 = 7'he == total_offset_4[6:0] ? phv_data_14 : _GEN_401; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_403 = 7'hf == total_offset_4[6:0] ? phv_data_15 : _GEN_402; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_404 = 7'h10 == total_offset_4[6:0] ? phv_data_16 : _GEN_403; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_405 = 7'h11 == total_offset_4[6:0] ? phv_data_17 : _GEN_404; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_406 = 7'h12 == total_offset_4[6:0] ? phv_data_18 : _GEN_405; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_407 = 7'h13 == total_offset_4[6:0] ? phv_data_19 : _GEN_406; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_408 = 7'h14 == total_offset_4[6:0] ? phv_data_20 : _GEN_407; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_409 = 7'h15 == total_offset_4[6:0] ? phv_data_21 : _GEN_408; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_410 = 7'h16 == total_offset_4[6:0] ? phv_data_22 : _GEN_409; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_411 = 7'h17 == total_offset_4[6:0] ? phv_data_23 : _GEN_410; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_412 = 7'h18 == total_offset_4[6:0] ? phv_data_24 : _GEN_411; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_413 = 7'h19 == total_offset_4[6:0] ? phv_data_25 : _GEN_412; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_414 = 7'h1a == total_offset_4[6:0] ? phv_data_26 : _GEN_413; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_415 = 7'h1b == total_offset_4[6:0] ? phv_data_27 : _GEN_414; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_416 = 7'h1c == total_offset_4[6:0] ? phv_data_28 : _GEN_415; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_417 = 7'h1d == total_offset_4[6:0] ? phv_data_29 : _GEN_416; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_418 = 7'h1e == total_offset_4[6:0] ? phv_data_30 : _GEN_417; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_419 = 7'h1f == total_offset_4[6:0] ? phv_data_31 : _GEN_418; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_420 = 7'h20 == total_offset_4[6:0] ? phv_data_32 : _GEN_419; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_421 = 7'h21 == total_offset_4[6:0] ? phv_data_33 : _GEN_420; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_422 = 7'h22 == total_offset_4[6:0] ? phv_data_34 : _GEN_421; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_423 = 7'h23 == total_offset_4[6:0] ? phv_data_35 : _GEN_422; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_424 = 7'h24 == total_offset_4[6:0] ? phv_data_36 : _GEN_423; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_425 = 7'h25 == total_offset_4[6:0] ? phv_data_37 : _GEN_424; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_426 = 7'h26 == total_offset_4[6:0] ? phv_data_38 : _GEN_425; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_427 = 7'h27 == total_offset_4[6:0] ? phv_data_39 : _GEN_426; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_428 = 7'h28 == total_offset_4[6:0] ? phv_data_40 : _GEN_427; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_429 = 7'h29 == total_offset_4[6:0] ? phv_data_41 : _GEN_428; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_430 = 7'h2a == total_offset_4[6:0] ? phv_data_42 : _GEN_429; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_431 = 7'h2b == total_offset_4[6:0] ? phv_data_43 : _GEN_430; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_432 = 7'h2c == total_offset_4[6:0] ? phv_data_44 : _GEN_431; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_433 = 7'h2d == total_offset_4[6:0] ? phv_data_45 : _GEN_432; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_434 = 7'h2e == total_offset_4[6:0] ? phv_data_46 : _GEN_433; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_435 = 7'h2f == total_offset_4[6:0] ? phv_data_47 : _GEN_434; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_436 = 7'h30 == total_offset_4[6:0] ? phv_data_48 : _GEN_435; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_437 = 7'h31 == total_offset_4[6:0] ? phv_data_49 : _GEN_436; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_438 = 7'h32 == total_offset_4[6:0] ? phv_data_50 : _GEN_437; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_439 = 7'h33 == total_offset_4[6:0] ? phv_data_51 : _GEN_438; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_440 = 7'h34 == total_offset_4[6:0] ? phv_data_52 : _GEN_439; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_441 = 7'h35 == total_offset_4[6:0] ? phv_data_53 : _GEN_440; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_442 = 7'h36 == total_offset_4[6:0] ? phv_data_54 : _GEN_441; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_443 = 7'h37 == total_offset_4[6:0] ? phv_data_55 : _GEN_442; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_444 = 7'h38 == total_offset_4[6:0] ? phv_data_56 : _GEN_443; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_445 = 7'h39 == total_offset_4[6:0] ? phv_data_57 : _GEN_444; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_446 = 7'h3a == total_offset_4[6:0] ? phv_data_58 : _GEN_445; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_447 = 7'h3b == total_offset_4[6:0] ? phv_data_59 : _GEN_446; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_448 = 7'h3c == total_offset_4[6:0] ? phv_data_60 : _GEN_447; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_449 = 7'h3d == total_offset_4[6:0] ? phv_data_61 : _GEN_448; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_450 = 7'h3e == total_offset_4[6:0] ? phv_data_62 : _GEN_449; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_451 = 7'h3f == total_offset_4[6:0] ? phv_data_63 : _GEN_450; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_452 = 7'h40 == total_offset_4[6:0] ? phv_data_64 : _GEN_451; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_453 = 7'h41 == total_offset_4[6:0] ? phv_data_65 : _GEN_452; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_454 = 7'h42 == total_offset_4[6:0] ? phv_data_66 : _GEN_453; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_455 = 7'h43 == total_offset_4[6:0] ? phv_data_67 : _GEN_454; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_456 = 7'h44 == total_offset_4[6:0] ? phv_data_68 : _GEN_455; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_457 = 7'h45 == total_offset_4[6:0] ? phv_data_69 : _GEN_456; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_458 = 7'h46 == total_offset_4[6:0] ? phv_data_70 : _GEN_457; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_459 = 7'h47 == total_offset_4[6:0] ? phv_data_71 : _GEN_458; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_460 = 7'h48 == total_offset_4[6:0] ? phv_data_72 : _GEN_459; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_461 = 7'h49 == total_offset_4[6:0] ? phv_data_73 : _GEN_460; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_462 = 7'h4a == total_offset_4[6:0] ? phv_data_74 : _GEN_461; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_463 = 7'h4b == total_offset_4[6:0] ? phv_data_75 : _GEN_462; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_464 = 7'h4c == total_offset_4[6:0] ? phv_data_76 : _GEN_463; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_465 = 7'h4d == total_offset_4[6:0] ? phv_data_77 : _GEN_464; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_466 = 7'h4e == total_offset_4[6:0] ? phv_data_78 : _GEN_465; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_467 = 7'h4f == total_offset_4[6:0] ? phv_data_79 : _GEN_466; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_468 = 7'h50 == total_offset_4[6:0] ? phv_data_80 : _GEN_467; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_469 = 7'h51 == total_offset_4[6:0] ? phv_data_81 : _GEN_468; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_470 = 7'h52 == total_offset_4[6:0] ? phv_data_82 : _GEN_469; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_471 = 7'h53 == total_offset_4[6:0] ? phv_data_83 : _GEN_470; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_472 = 7'h54 == total_offset_4[6:0] ? phv_data_84 : _GEN_471; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_473 = 7'h55 == total_offset_4[6:0] ? phv_data_85 : _GEN_472; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_474 = 7'h56 == total_offset_4[6:0] ? phv_data_86 : _GEN_473; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_475 = 7'h57 == total_offset_4[6:0] ? phv_data_87 : _GEN_474; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_476 = 7'h58 == total_offset_4[6:0] ? phv_data_88 : _GEN_475; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_477 = 7'h59 == total_offset_4[6:0] ? phv_data_89 : _GEN_476; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_478 = 7'h5a == total_offset_4[6:0] ? phv_data_90 : _GEN_477; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_479 = 7'h5b == total_offset_4[6:0] ? phv_data_91 : _GEN_478; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_480 = 7'h5c == total_offset_4[6:0] ? phv_data_92 : _GEN_479; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_481 = 7'h5d == total_offset_4[6:0] ? phv_data_93 : _GEN_480; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_482 = 7'h5e == total_offset_4[6:0] ? phv_data_94 : _GEN_481; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_483 = 7'h5f == total_offset_4[6:0] ? phv_data_95 : _GEN_482; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes__4 = 8'h4 < length_0 ? _GEN_483 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_5 = offset_0 + 8'h5; // @[executor.scala 158:57]
  wire [7:0] _GEN_486 = 7'h1 == total_offset_5[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_487 = 7'h2 == total_offset_5[6:0] ? phv_data_2 : _GEN_486; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_488 = 7'h3 == total_offset_5[6:0] ? phv_data_3 : _GEN_487; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_489 = 7'h4 == total_offset_5[6:0] ? phv_data_4 : _GEN_488; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_490 = 7'h5 == total_offset_5[6:0] ? phv_data_5 : _GEN_489; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_491 = 7'h6 == total_offset_5[6:0] ? phv_data_6 : _GEN_490; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_492 = 7'h7 == total_offset_5[6:0] ? phv_data_7 : _GEN_491; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_493 = 7'h8 == total_offset_5[6:0] ? phv_data_8 : _GEN_492; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_494 = 7'h9 == total_offset_5[6:0] ? phv_data_9 : _GEN_493; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_495 = 7'ha == total_offset_5[6:0] ? phv_data_10 : _GEN_494; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_496 = 7'hb == total_offset_5[6:0] ? phv_data_11 : _GEN_495; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_497 = 7'hc == total_offset_5[6:0] ? phv_data_12 : _GEN_496; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_498 = 7'hd == total_offset_5[6:0] ? phv_data_13 : _GEN_497; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_499 = 7'he == total_offset_5[6:0] ? phv_data_14 : _GEN_498; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_500 = 7'hf == total_offset_5[6:0] ? phv_data_15 : _GEN_499; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_501 = 7'h10 == total_offset_5[6:0] ? phv_data_16 : _GEN_500; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_502 = 7'h11 == total_offset_5[6:0] ? phv_data_17 : _GEN_501; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_503 = 7'h12 == total_offset_5[6:0] ? phv_data_18 : _GEN_502; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_504 = 7'h13 == total_offset_5[6:0] ? phv_data_19 : _GEN_503; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_505 = 7'h14 == total_offset_5[6:0] ? phv_data_20 : _GEN_504; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_506 = 7'h15 == total_offset_5[6:0] ? phv_data_21 : _GEN_505; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_507 = 7'h16 == total_offset_5[6:0] ? phv_data_22 : _GEN_506; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_508 = 7'h17 == total_offset_5[6:0] ? phv_data_23 : _GEN_507; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_509 = 7'h18 == total_offset_5[6:0] ? phv_data_24 : _GEN_508; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_510 = 7'h19 == total_offset_5[6:0] ? phv_data_25 : _GEN_509; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_511 = 7'h1a == total_offset_5[6:0] ? phv_data_26 : _GEN_510; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_512 = 7'h1b == total_offset_5[6:0] ? phv_data_27 : _GEN_511; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_513 = 7'h1c == total_offset_5[6:0] ? phv_data_28 : _GEN_512; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_514 = 7'h1d == total_offset_5[6:0] ? phv_data_29 : _GEN_513; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_515 = 7'h1e == total_offset_5[6:0] ? phv_data_30 : _GEN_514; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_516 = 7'h1f == total_offset_5[6:0] ? phv_data_31 : _GEN_515; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_517 = 7'h20 == total_offset_5[6:0] ? phv_data_32 : _GEN_516; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_518 = 7'h21 == total_offset_5[6:0] ? phv_data_33 : _GEN_517; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_519 = 7'h22 == total_offset_5[6:0] ? phv_data_34 : _GEN_518; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_520 = 7'h23 == total_offset_5[6:0] ? phv_data_35 : _GEN_519; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_521 = 7'h24 == total_offset_5[6:0] ? phv_data_36 : _GEN_520; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_522 = 7'h25 == total_offset_5[6:0] ? phv_data_37 : _GEN_521; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_523 = 7'h26 == total_offset_5[6:0] ? phv_data_38 : _GEN_522; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_524 = 7'h27 == total_offset_5[6:0] ? phv_data_39 : _GEN_523; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_525 = 7'h28 == total_offset_5[6:0] ? phv_data_40 : _GEN_524; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_526 = 7'h29 == total_offset_5[6:0] ? phv_data_41 : _GEN_525; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_527 = 7'h2a == total_offset_5[6:0] ? phv_data_42 : _GEN_526; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_528 = 7'h2b == total_offset_5[6:0] ? phv_data_43 : _GEN_527; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_529 = 7'h2c == total_offset_5[6:0] ? phv_data_44 : _GEN_528; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_530 = 7'h2d == total_offset_5[6:0] ? phv_data_45 : _GEN_529; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_531 = 7'h2e == total_offset_5[6:0] ? phv_data_46 : _GEN_530; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_532 = 7'h2f == total_offset_5[6:0] ? phv_data_47 : _GEN_531; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_533 = 7'h30 == total_offset_5[6:0] ? phv_data_48 : _GEN_532; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_534 = 7'h31 == total_offset_5[6:0] ? phv_data_49 : _GEN_533; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_535 = 7'h32 == total_offset_5[6:0] ? phv_data_50 : _GEN_534; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_536 = 7'h33 == total_offset_5[6:0] ? phv_data_51 : _GEN_535; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_537 = 7'h34 == total_offset_5[6:0] ? phv_data_52 : _GEN_536; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_538 = 7'h35 == total_offset_5[6:0] ? phv_data_53 : _GEN_537; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_539 = 7'h36 == total_offset_5[6:0] ? phv_data_54 : _GEN_538; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_540 = 7'h37 == total_offset_5[6:0] ? phv_data_55 : _GEN_539; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_541 = 7'h38 == total_offset_5[6:0] ? phv_data_56 : _GEN_540; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_542 = 7'h39 == total_offset_5[6:0] ? phv_data_57 : _GEN_541; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_543 = 7'h3a == total_offset_5[6:0] ? phv_data_58 : _GEN_542; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_544 = 7'h3b == total_offset_5[6:0] ? phv_data_59 : _GEN_543; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_545 = 7'h3c == total_offset_5[6:0] ? phv_data_60 : _GEN_544; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_546 = 7'h3d == total_offset_5[6:0] ? phv_data_61 : _GEN_545; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_547 = 7'h3e == total_offset_5[6:0] ? phv_data_62 : _GEN_546; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_548 = 7'h3f == total_offset_5[6:0] ? phv_data_63 : _GEN_547; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_549 = 7'h40 == total_offset_5[6:0] ? phv_data_64 : _GEN_548; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_550 = 7'h41 == total_offset_5[6:0] ? phv_data_65 : _GEN_549; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_551 = 7'h42 == total_offset_5[6:0] ? phv_data_66 : _GEN_550; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_552 = 7'h43 == total_offset_5[6:0] ? phv_data_67 : _GEN_551; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_553 = 7'h44 == total_offset_5[6:0] ? phv_data_68 : _GEN_552; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_554 = 7'h45 == total_offset_5[6:0] ? phv_data_69 : _GEN_553; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_555 = 7'h46 == total_offset_5[6:0] ? phv_data_70 : _GEN_554; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_556 = 7'h47 == total_offset_5[6:0] ? phv_data_71 : _GEN_555; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_557 = 7'h48 == total_offset_5[6:0] ? phv_data_72 : _GEN_556; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_558 = 7'h49 == total_offset_5[6:0] ? phv_data_73 : _GEN_557; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_559 = 7'h4a == total_offset_5[6:0] ? phv_data_74 : _GEN_558; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_560 = 7'h4b == total_offset_5[6:0] ? phv_data_75 : _GEN_559; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_561 = 7'h4c == total_offset_5[6:0] ? phv_data_76 : _GEN_560; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_562 = 7'h4d == total_offset_5[6:0] ? phv_data_77 : _GEN_561; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_563 = 7'h4e == total_offset_5[6:0] ? phv_data_78 : _GEN_562; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_564 = 7'h4f == total_offset_5[6:0] ? phv_data_79 : _GEN_563; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_565 = 7'h50 == total_offset_5[6:0] ? phv_data_80 : _GEN_564; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_566 = 7'h51 == total_offset_5[6:0] ? phv_data_81 : _GEN_565; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_567 = 7'h52 == total_offset_5[6:0] ? phv_data_82 : _GEN_566; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_568 = 7'h53 == total_offset_5[6:0] ? phv_data_83 : _GEN_567; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_569 = 7'h54 == total_offset_5[6:0] ? phv_data_84 : _GEN_568; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_570 = 7'h55 == total_offset_5[6:0] ? phv_data_85 : _GEN_569; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_571 = 7'h56 == total_offset_5[6:0] ? phv_data_86 : _GEN_570; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_572 = 7'h57 == total_offset_5[6:0] ? phv_data_87 : _GEN_571; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_573 = 7'h58 == total_offset_5[6:0] ? phv_data_88 : _GEN_572; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_574 = 7'h59 == total_offset_5[6:0] ? phv_data_89 : _GEN_573; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_575 = 7'h5a == total_offset_5[6:0] ? phv_data_90 : _GEN_574; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_576 = 7'h5b == total_offset_5[6:0] ? phv_data_91 : _GEN_575; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_577 = 7'h5c == total_offset_5[6:0] ? phv_data_92 : _GEN_576; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_578 = 7'h5d == total_offset_5[6:0] ? phv_data_93 : _GEN_577; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_579 = 7'h5e == total_offset_5[6:0] ? phv_data_94 : _GEN_578; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_580 = 7'h5f == total_offset_5[6:0] ? phv_data_95 : _GEN_579; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes__5 = 8'h5 < length_0 ? _GEN_580 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_6 = offset_0 + 8'h6; // @[executor.scala 158:57]
  wire [7:0] _GEN_583 = 7'h1 == total_offset_6[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_584 = 7'h2 == total_offset_6[6:0] ? phv_data_2 : _GEN_583; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_585 = 7'h3 == total_offset_6[6:0] ? phv_data_3 : _GEN_584; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_586 = 7'h4 == total_offset_6[6:0] ? phv_data_4 : _GEN_585; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_587 = 7'h5 == total_offset_6[6:0] ? phv_data_5 : _GEN_586; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_588 = 7'h6 == total_offset_6[6:0] ? phv_data_6 : _GEN_587; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_589 = 7'h7 == total_offset_6[6:0] ? phv_data_7 : _GEN_588; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_590 = 7'h8 == total_offset_6[6:0] ? phv_data_8 : _GEN_589; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_591 = 7'h9 == total_offset_6[6:0] ? phv_data_9 : _GEN_590; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_592 = 7'ha == total_offset_6[6:0] ? phv_data_10 : _GEN_591; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_593 = 7'hb == total_offset_6[6:0] ? phv_data_11 : _GEN_592; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_594 = 7'hc == total_offset_6[6:0] ? phv_data_12 : _GEN_593; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_595 = 7'hd == total_offset_6[6:0] ? phv_data_13 : _GEN_594; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_596 = 7'he == total_offset_6[6:0] ? phv_data_14 : _GEN_595; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_597 = 7'hf == total_offset_6[6:0] ? phv_data_15 : _GEN_596; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_598 = 7'h10 == total_offset_6[6:0] ? phv_data_16 : _GEN_597; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_599 = 7'h11 == total_offset_6[6:0] ? phv_data_17 : _GEN_598; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_600 = 7'h12 == total_offset_6[6:0] ? phv_data_18 : _GEN_599; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_601 = 7'h13 == total_offset_6[6:0] ? phv_data_19 : _GEN_600; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_602 = 7'h14 == total_offset_6[6:0] ? phv_data_20 : _GEN_601; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_603 = 7'h15 == total_offset_6[6:0] ? phv_data_21 : _GEN_602; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_604 = 7'h16 == total_offset_6[6:0] ? phv_data_22 : _GEN_603; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_605 = 7'h17 == total_offset_6[6:0] ? phv_data_23 : _GEN_604; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_606 = 7'h18 == total_offset_6[6:0] ? phv_data_24 : _GEN_605; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_607 = 7'h19 == total_offset_6[6:0] ? phv_data_25 : _GEN_606; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_608 = 7'h1a == total_offset_6[6:0] ? phv_data_26 : _GEN_607; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_609 = 7'h1b == total_offset_6[6:0] ? phv_data_27 : _GEN_608; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_610 = 7'h1c == total_offset_6[6:0] ? phv_data_28 : _GEN_609; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_611 = 7'h1d == total_offset_6[6:0] ? phv_data_29 : _GEN_610; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_612 = 7'h1e == total_offset_6[6:0] ? phv_data_30 : _GEN_611; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_613 = 7'h1f == total_offset_6[6:0] ? phv_data_31 : _GEN_612; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_614 = 7'h20 == total_offset_6[6:0] ? phv_data_32 : _GEN_613; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_615 = 7'h21 == total_offset_6[6:0] ? phv_data_33 : _GEN_614; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_616 = 7'h22 == total_offset_6[6:0] ? phv_data_34 : _GEN_615; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_617 = 7'h23 == total_offset_6[6:0] ? phv_data_35 : _GEN_616; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_618 = 7'h24 == total_offset_6[6:0] ? phv_data_36 : _GEN_617; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_619 = 7'h25 == total_offset_6[6:0] ? phv_data_37 : _GEN_618; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_620 = 7'h26 == total_offset_6[6:0] ? phv_data_38 : _GEN_619; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_621 = 7'h27 == total_offset_6[6:0] ? phv_data_39 : _GEN_620; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_622 = 7'h28 == total_offset_6[6:0] ? phv_data_40 : _GEN_621; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_623 = 7'h29 == total_offset_6[6:0] ? phv_data_41 : _GEN_622; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_624 = 7'h2a == total_offset_6[6:0] ? phv_data_42 : _GEN_623; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_625 = 7'h2b == total_offset_6[6:0] ? phv_data_43 : _GEN_624; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_626 = 7'h2c == total_offset_6[6:0] ? phv_data_44 : _GEN_625; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_627 = 7'h2d == total_offset_6[6:0] ? phv_data_45 : _GEN_626; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_628 = 7'h2e == total_offset_6[6:0] ? phv_data_46 : _GEN_627; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_629 = 7'h2f == total_offset_6[6:0] ? phv_data_47 : _GEN_628; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_630 = 7'h30 == total_offset_6[6:0] ? phv_data_48 : _GEN_629; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_631 = 7'h31 == total_offset_6[6:0] ? phv_data_49 : _GEN_630; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_632 = 7'h32 == total_offset_6[6:0] ? phv_data_50 : _GEN_631; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_633 = 7'h33 == total_offset_6[6:0] ? phv_data_51 : _GEN_632; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_634 = 7'h34 == total_offset_6[6:0] ? phv_data_52 : _GEN_633; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_635 = 7'h35 == total_offset_6[6:0] ? phv_data_53 : _GEN_634; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_636 = 7'h36 == total_offset_6[6:0] ? phv_data_54 : _GEN_635; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_637 = 7'h37 == total_offset_6[6:0] ? phv_data_55 : _GEN_636; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_638 = 7'h38 == total_offset_6[6:0] ? phv_data_56 : _GEN_637; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_639 = 7'h39 == total_offset_6[6:0] ? phv_data_57 : _GEN_638; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_640 = 7'h3a == total_offset_6[6:0] ? phv_data_58 : _GEN_639; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_641 = 7'h3b == total_offset_6[6:0] ? phv_data_59 : _GEN_640; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_642 = 7'h3c == total_offset_6[6:0] ? phv_data_60 : _GEN_641; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_643 = 7'h3d == total_offset_6[6:0] ? phv_data_61 : _GEN_642; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_644 = 7'h3e == total_offset_6[6:0] ? phv_data_62 : _GEN_643; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_645 = 7'h3f == total_offset_6[6:0] ? phv_data_63 : _GEN_644; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_646 = 7'h40 == total_offset_6[6:0] ? phv_data_64 : _GEN_645; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_647 = 7'h41 == total_offset_6[6:0] ? phv_data_65 : _GEN_646; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_648 = 7'h42 == total_offset_6[6:0] ? phv_data_66 : _GEN_647; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_649 = 7'h43 == total_offset_6[6:0] ? phv_data_67 : _GEN_648; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_650 = 7'h44 == total_offset_6[6:0] ? phv_data_68 : _GEN_649; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_651 = 7'h45 == total_offset_6[6:0] ? phv_data_69 : _GEN_650; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_652 = 7'h46 == total_offset_6[6:0] ? phv_data_70 : _GEN_651; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_653 = 7'h47 == total_offset_6[6:0] ? phv_data_71 : _GEN_652; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_654 = 7'h48 == total_offset_6[6:0] ? phv_data_72 : _GEN_653; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_655 = 7'h49 == total_offset_6[6:0] ? phv_data_73 : _GEN_654; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_656 = 7'h4a == total_offset_6[6:0] ? phv_data_74 : _GEN_655; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_657 = 7'h4b == total_offset_6[6:0] ? phv_data_75 : _GEN_656; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_658 = 7'h4c == total_offset_6[6:0] ? phv_data_76 : _GEN_657; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_659 = 7'h4d == total_offset_6[6:0] ? phv_data_77 : _GEN_658; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_660 = 7'h4e == total_offset_6[6:0] ? phv_data_78 : _GEN_659; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_661 = 7'h4f == total_offset_6[6:0] ? phv_data_79 : _GEN_660; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_662 = 7'h50 == total_offset_6[6:0] ? phv_data_80 : _GEN_661; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_663 = 7'h51 == total_offset_6[6:0] ? phv_data_81 : _GEN_662; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_664 = 7'h52 == total_offset_6[6:0] ? phv_data_82 : _GEN_663; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_665 = 7'h53 == total_offset_6[6:0] ? phv_data_83 : _GEN_664; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_666 = 7'h54 == total_offset_6[6:0] ? phv_data_84 : _GEN_665; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_667 = 7'h55 == total_offset_6[6:0] ? phv_data_85 : _GEN_666; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_668 = 7'h56 == total_offset_6[6:0] ? phv_data_86 : _GEN_667; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_669 = 7'h57 == total_offset_6[6:0] ? phv_data_87 : _GEN_668; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_670 = 7'h58 == total_offset_6[6:0] ? phv_data_88 : _GEN_669; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_671 = 7'h59 == total_offset_6[6:0] ? phv_data_89 : _GEN_670; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_672 = 7'h5a == total_offset_6[6:0] ? phv_data_90 : _GEN_671; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_673 = 7'h5b == total_offset_6[6:0] ? phv_data_91 : _GEN_672; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_674 = 7'h5c == total_offset_6[6:0] ? phv_data_92 : _GEN_673; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_675 = 7'h5d == total_offset_6[6:0] ? phv_data_93 : _GEN_674; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_676 = 7'h5e == total_offset_6[6:0] ? phv_data_94 : _GEN_675; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_677 = 7'h5f == total_offset_6[6:0] ? phv_data_95 : _GEN_676; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes__6 = 8'h6 < length_0 ? _GEN_677 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_7 = offset_0 + 8'h7; // @[executor.scala 158:57]
  wire [7:0] _GEN_680 = 7'h1 == total_offset_7[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_681 = 7'h2 == total_offset_7[6:0] ? phv_data_2 : _GEN_680; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_682 = 7'h3 == total_offset_7[6:0] ? phv_data_3 : _GEN_681; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_683 = 7'h4 == total_offset_7[6:0] ? phv_data_4 : _GEN_682; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_684 = 7'h5 == total_offset_7[6:0] ? phv_data_5 : _GEN_683; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_685 = 7'h6 == total_offset_7[6:0] ? phv_data_6 : _GEN_684; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_686 = 7'h7 == total_offset_7[6:0] ? phv_data_7 : _GEN_685; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_687 = 7'h8 == total_offset_7[6:0] ? phv_data_8 : _GEN_686; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_688 = 7'h9 == total_offset_7[6:0] ? phv_data_9 : _GEN_687; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_689 = 7'ha == total_offset_7[6:0] ? phv_data_10 : _GEN_688; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_690 = 7'hb == total_offset_7[6:0] ? phv_data_11 : _GEN_689; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_691 = 7'hc == total_offset_7[6:0] ? phv_data_12 : _GEN_690; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_692 = 7'hd == total_offset_7[6:0] ? phv_data_13 : _GEN_691; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_693 = 7'he == total_offset_7[6:0] ? phv_data_14 : _GEN_692; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_694 = 7'hf == total_offset_7[6:0] ? phv_data_15 : _GEN_693; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_695 = 7'h10 == total_offset_7[6:0] ? phv_data_16 : _GEN_694; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_696 = 7'h11 == total_offset_7[6:0] ? phv_data_17 : _GEN_695; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_697 = 7'h12 == total_offset_7[6:0] ? phv_data_18 : _GEN_696; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_698 = 7'h13 == total_offset_7[6:0] ? phv_data_19 : _GEN_697; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_699 = 7'h14 == total_offset_7[6:0] ? phv_data_20 : _GEN_698; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_700 = 7'h15 == total_offset_7[6:0] ? phv_data_21 : _GEN_699; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_701 = 7'h16 == total_offset_7[6:0] ? phv_data_22 : _GEN_700; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_702 = 7'h17 == total_offset_7[6:0] ? phv_data_23 : _GEN_701; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_703 = 7'h18 == total_offset_7[6:0] ? phv_data_24 : _GEN_702; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_704 = 7'h19 == total_offset_7[6:0] ? phv_data_25 : _GEN_703; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_705 = 7'h1a == total_offset_7[6:0] ? phv_data_26 : _GEN_704; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_706 = 7'h1b == total_offset_7[6:0] ? phv_data_27 : _GEN_705; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_707 = 7'h1c == total_offset_7[6:0] ? phv_data_28 : _GEN_706; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_708 = 7'h1d == total_offset_7[6:0] ? phv_data_29 : _GEN_707; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_709 = 7'h1e == total_offset_7[6:0] ? phv_data_30 : _GEN_708; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_710 = 7'h1f == total_offset_7[6:0] ? phv_data_31 : _GEN_709; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_711 = 7'h20 == total_offset_7[6:0] ? phv_data_32 : _GEN_710; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_712 = 7'h21 == total_offset_7[6:0] ? phv_data_33 : _GEN_711; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_713 = 7'h22 == total_offset_7[6:0] ? phv_data_34 : _GEN_712; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_714 = 7'h23 == total_offset_7[6:0] ? phv_data_35 : _GEN_713; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_715 = 7'h24 == total_offset_7[6:0] ? phv_data_36 : _GEN_714; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_716 = 7'h25 == total_offset_7[6:0] ? phv_data_37 : _GEN_715; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_717 = 7'h26 == total_offset_7[6:0] ? phv_data_38 : _GEN_716; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_718 = 7'h27 == total_offset_7[6:0] ? phv_data_39 : _GEN_717; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_719 = 7'h28 == total_offset_7[6:0] ? phv_data_40 : _GEN_718; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_720 = 7'h29 == total_offset_7[6:0] ? phv_data_41 : _GEN_719; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_721 = 7'h2a == total_offset_7[6:0] ? phv_data_42 : _GEN_720; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_722 = 7'h2b == total_offset_7[6:0] ? phv_data_43 : _GEN_721; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_723 = 7'h2c == total_offset_7[6:0] ? phv_data_44 : _GEN_722; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_724 = 7'h2d == total_offset_7[6:0] ? phv_data_45 : _GEN_723; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_725 = 7'h2e == total_offset_7[6:0] ? phv_data_46 : _GEN_724; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_726 = 7'h2f == total_offset_7[6:0] ? phv_data_47 : _GEN_725; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_727 = 7'h30 == total_offset_7[6:0] ? phv_data_48 : _GEN_726; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_728 = 7'h31 == total_offset_7[6:0] ? phv_data_49 : _GEN_727; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_729 = 7'h32 == total_offset_7[6:0] ? phv_data_50 : _GEN_728; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_730 = 7'h33 == total_offset_7[6:0] ? phv_data_51 : _GEN_729; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_731 = 7'h34 == total_offset_7[6:0] ? phv_data_52 : _GEN_730; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_732 = 7'h35 == total_offset_7[6:0] ? phv_data_53 : _GEN_731; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_733 = 7'h36 == total_offset_7[6:0] ? phv_data_54 : _GEN_732; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_734 = 7'h37 == total_offset_7[6:0] ? phv_data_55 : _GEN_733; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_735 = 7'h38 == total_offset_7[6:0] ? phv_data_56 : _GEN_734; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_736 = 7'h39 == total_offset_7[6:0] ? phv_data_57 : _GEN_735; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_737 = 7'h3a == total_offset_7[6:0] ? phv_data_58 : _GEN_736; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_738 = 7'h3b == total_offset_7[6:0] ? phv_data_59 : _GEN_737; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_739 = 7'h3c == total_offset_7[6:0] ? phv_data_60 : _GEN_738; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_740 = 7'h3d == total_offset_7[6:0] ? phv_data_61 : _GEN_739; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_741 = 7'h3e == total_offset_7[6:0] ? phv_data_62 : _GEN_740; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_742 = 7'h3f == total_offset_7[6:0] ? phv_data_63 : _GEN_741; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_743 = 7'h40 == total_offset_7[6:0] ? phv_data_64 : _GEN_742; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_744 = 7'h41 == total_offset_7[6:0] ? phv_data_65 : _GEN_743; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_745 = 7'h42 == total_offset_7[6:0] ? phv_data_66 : _GEN_744; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_746 = 7'h43 == total_offset_7[6:0] ? phv_data_67 : _GEN_745; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_747 = 7'h44 == total_offset_7[6:0] ? phv_data_68 : _GEN_746; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_748 = 7'h45 == total_offset_7[6:0] ? phv_data_69 : _GEN_747; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_749 = 7'h46 == total_offset_7[6:0] ? phv_data_70 : _GEN_748; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_750 = 7'h47 == total_offset_7[6:0] ? phv_data_71 : _GEN_749; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_751 = 7'h48 == total_offset_7[6:0] ? phv_data_72 : _GEN_750; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_752 = 7'h49 == total_offset_7[6:0] ? phv_data_73 : _GEN_751; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_753 = 7'h4a == total_offset_7[6:0] ? phv_data_74 : _GEN_752; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_754 = 7'h4b == total_offset_7[6:0] ? phv_data_75 : _GEN_753; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_755 = 7'h4c == total_offset_7[6:0] ? phv_data_76 : _GEN_754; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_756 = 7'h4d == total_offset_7[6:0] ? phv_data_77 : _GEN_755; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_757 = 7'h4e == total_offset_7[6:0] ? phv_data_78 : _GEN_756; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_758 = 7'h4f == total_offset_7[6:0] ? phv_data_79 : _GEN_757; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_759 = 7'h50 == total_offset_7[6:0] ? phv_data_80 : _GEN_758; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_760 = 7'h51 == total_offset_7[6:0] ? phv_data_81 : _GEN_759; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_761 = 7'h52 == total_offset_7[6:0] ? phv_data_82 : _GEN_760; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_762 = 7'h53 == total_offset_7[6:0] ? phv_data_83 : _GEN_761; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_763 = 7'h54 == total_offset_7[6:0] ? phv_data_84 : _GEN_762; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_764 = 7'h55 == total_offset_7[6:0] ? phv_data_85 : _GEN_763; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_765 = 7'h56 == total_offset_7[6:0] ? phv_data_86 : _GEN_764; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_766 = 7'h57 == total_offset_7[6:0] ? phv_data_87 : _GEN_765; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_767 = 7'h58 == total_offset_7[6:0] ? phv_data_88 : _GEN_766; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_768 = 7'h59 == total_offset_7[6:0] ? phv_data_89 : _GEN_767; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_769 = 7'h5a == total_offset_7[6:0] ? phv_data_90 : _GEN_768; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_770 = 7'h5b == total_offset_7[6:0] ? phv_data_91 : _GEN_769; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_771 = 7'h5c == total_offset_7[6:0] ? phv_data_92 : _GEN_770; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_772 = 7'h5d == total_offset_7[6:0] ? phv_data_93 : _GEN_771; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_773 = 7'h5e == total_offset_7[6:0] ? phv_data_94 : _GEN_772; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_774 = 7'h5f == total_offset_7[6:0] ? phv_data_95 : _GEN_773; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes__7 = 8'h7 < length_0 ? _GEN_774 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [63:0] _io_field_out_0_T = {bytes__0,bytes__1,bytes__2,bytes__3,bytes__4,bytes__5,bytes__6,bytes__7}; // @[Cat.scala 30:58]
  wire [2:0] args_offset = io_field_out_0_lo[13:11]; // @[primitive.scala 34:52]
  wire [2:0] args_length = io_field_out_0_lo[10:8]; // @[primitive.scala 35:52]
  wire [8:0] _total_offset_T_8 = {{6'd0}, args_offset}; // @[executor.scala 173:60]
  wire [7:0] total_offset_8 = _total_offset_T_8[7:0]; // @[executor.scala 173:60]
  wire [7:0] _GEN_3372 = {{5'd0}, args_length}; // @[executor.scala 174:48]
  wire [7:0] _GEN_777 = 3'h1 == total_offset_8[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_778 = 3'h2 == total_offset_8[2:0] ? args_2 : _GEN_777; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_779 = 3'h3 == total_offset_8[2:0] ? args_3 : _GEN_778; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_780 = 3'h4 == total_offset_8[2:0] ? args_4 : _GEN_779; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_781 = 3'h5 == total_offset_8[2:0] ? args_5 : _GEN_780; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_782 = 3'h6 == total_offset_8[2:0] ? args_6 : _GEN_781; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_1_0 = 8'h0 < _GEN_3372 ? _GEN_782 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [7:0] _GEN_3373 = {{5'd0}, args_offset}; // @[executor.scala 173:60]
  wire [7:0] total_offset_9 = _GEN_3373 + 8'h1; // @[executor.scala 173:60]
  wire [7:0] _GEN_785 = 3'h1 == total_offset_9[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_786 = 3'h2 == total_offset_9[2:0] ? args_2 : _GEN_785; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_787 = 3'h3 == total_offset_9[2:0] ? args_3 : _GEN_786; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_788 = 3'h4 == total_offset_9[2:0] ? args_4 : _GEN_787; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_789 = 3'h5 == total_offset_9[2:0] ? args_5 : _GEN_788; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_790 = 3'h6 == total_offset_9[2:0] ? args_6 : _GEN_789; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_1_1 = 8'h1 < _GEN_3372 ? _GEN_790 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [7:0] total_offset_10 = _GEN_3373 + 8'h2; // @[executor.scala 173:60]
  wire [7:0] _GEN_793 = 3'h1 == total_offset_10[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_794 = 3'h2 == total_offset_10[2:0] ? args_2 : _GEN_793; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_795 = 3'h3 == total_offset_10[2:0] ? args_3 : _GEN_794; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_796 = 3'h4 == total_offset_10[2:0] ? args_4 : _GEN_795; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_797 = 3'h5 == total_offset_10[2:0] ? args_5 : _GEN_796; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_798 = 3'h6 == total_offset_10[2:0] ? args_6 : _GEN_797; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_1_2 = 8'h2 < _GEN_3372 ? _GEN_798 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [7:0] total_offset_11 = _GEN_3373 + 8'h3; // @[executor.scala 173:60]
  wire [7:0] _GEN_801 = 3'h1 == total_offset_11[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_802 = 3'h2 == total_offset_11[2:0] ? args_2 : _GEN_801; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_803 = 3'h3 == total_offset_11[2:0] ? args_3 : _GEN_802; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_804 = 3'h4 == total_offset_11[2:0] ? args_4 : _GEN_803; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_805 = 3'h5 == total_offset_11[2:0] ? args_5 : _GEN_804; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_806 = 3'h6 == total_offset_11[2:0] ? args_6 : _GEN_805; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_1_3 = 8'h3 < _GEN_3372 ? _GEN_806 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [7:0] total_offset_12 = _GEN_3373 + 8'h4; // @[executor.scala 173:60]
  wire [7:0] _GEN_809 = 3'h1 == total_offset_12[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_810 = 3'h2 == total_offset_12[2:0] ? args_2 : _GEN_809; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_811 = 3'h3 == total_offset_12[2:0] ? args_3 : _GEN_810; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_812 = 3'h4 == total_offset_12[2:0] ? args_4 : _GEN_811; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_813 = 3'h5 == total_offset_12[2:0] ? args_5 : _GEN_812; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_814 = 3'h6 == total_offset_12[2:0] ? args_6 : _GEN_813; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_1_4 = 8'h4 < _GEN_3372 ? _GEN_814 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [7:0] total_offset_13 = _GEN_3373 + 8'h5; // @[executor.scala 173:60]
  wire [7:0] _GEN_817 = 3'h1 == total_offset_13[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_818 = 3'h2 == total_offset_13[2:0] ? args_2 : _GEN_817; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_819 = 3'h3 == total_offset_13[2:0] ? args_3 : _GEN_818; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_820 = 3'h4 == total_offset_13[2:0] ? args_4 : _GEN_819; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_821 = 3'h5 == total_offset_13[2:0] ? args_5 : _GEN_820; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_822 = 3'h6 == total_offset_13[2:0] ? args_6 : _GEN_821; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_1_5 = 8'h5 < _GEN_3372 ? _GEN_822 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [7:0] total_offset_14 = _GEN_3373 + 8'h6; // @[executor.scala 173:60]
  wire [7:0] _GEN_825 = 3'h1 == total_offset_14[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_826 = 3'h2 == total_offset_14[2:0] ? args_2 : _GEN_825; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_827 = 3'h3 == total_offset_14[2:0] ? args_3 : _GEN_826; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_828 = 3'h4 == total_offset_14[2:0] ? args_4 : _GEN_827; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_829 = 3'h5 == total_offset_14[2:0] ? args_5 : _GEN_828; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_830 = 3'h6 == total_offset_14[2:0] ? args_6 : _GEN_829; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_1_6 = 8'h6 < _GEN_3372 ? _GEN_830 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [63:0] _io_field_out_0_T_1 = {bytes_1_0,bytes_1_1,bytes_1_2,bytes_1_3,bytes_1_4,bytes_1_5,bytes_1_6,8'h0}; // @[Cat.scala 30:58]
  wire [49:0] io_field_out_0_hi_12 = io_field_out_0_lo[13] ? 50'h3ffffffffffff : 50'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _io_field_out_0_T_4 = {io_field_out_0_hi_12,io_field_out_0_lo}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_840 = 4'ha == opcode ? _io_field_out_0_T_1 : _io_field_out_0_T_4; // @[executor.scala 167:55 executor.scala 180:41 executor.scala 183:41]
  wire [63:0] _GEN_841 = from_header ? _io_field_out_0_T : _GEN_840; // @[executor.scala 152:36 executor.scala 165:37]
  wire [3:0] opcode_1 = vliw_1[31:28]; // @[primitive.scala 9:44]
  wire [13:0] io_field_out_1_lo = vliw_1[13:0]; // @[primitive.scala 11:44]
  wire  from_header_1 = length_1 != 8'h0; // @[executor.scala 151:45]
  wire [8:0] _total_offset_T_16 = {{1'd0}, offset_1}; // @[executor.scala 158:57]
  wire [7:0] total_offset_16 = _total_offset_T_16[7:0]; // @[executor.scala 158:57]
  wire [7:0] _GEN_844 = 7'h1 == total_offset_16[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_845 = 7'h2 == total_offset_16[6:0] ? phv_data_2 : _GEN_844; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_846 = 7'h3 == total_offset_16[6:0] ? phv_data_3 : _GEN_845; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_847 = 7'h4 == total_offset_16[6:0] ? phv_data_4 : _GEN_846; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_848 = 7'h5 == total_offset_16[6:0] ? phv_data_5 : _GEN_847; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_849 = 7'h6 == total_offset_16[6:0] ? phv_data_6 : _GEN_848; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_850 = 7'h7 == total_offset_16[6:0] ? phv_data_7 : _GEN_849; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_851 = 7'h8 == total_offset_16[6:0] ? phv_data_8 : _GEN_850; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_852 = 7'h9 == total_offset_16[6:0] ? phv_data_9 : _GEN_851; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_853 = 7'ha == total_offset_16[6:0] ? phv_data_10 : _GEN_852; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_854 = 7'hb == total_offset_16[6:0] ? phv_data_11 : _GEN_853; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_855 = 7'hc == total_offset_16[6:0] ? phv_data_12 : _GEN_854; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_856 = 7'hd == total_offset_16[6:0] ? phv_data_13 : _GEN_855; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_857 = 7'he == total_offset_16[6:0] ? phv_data_14 : _GEN_856; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_858 = 7'hf == total_offset_16[6:0] ? phv_data_15 : _GEN_857; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_859 = 7'h10 == total_offset_16[6:0] ? phv_data_16 : _GEN_858; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_860 = 7'h11 == total_offset_16[6:0] ? phv_data_17 : _GEN_859; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_861 = 7'h12 == total_offset_16[6:0] ? phv_data_18 : _GEN_860; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_862 = 7'h13 == total_offset_16[6:0] ? phv_data_19 : _GEN_861; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_863 = 7'h14 == total_offset_16[6:0] ? phv_data_20 : _GEN_862; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_864 = 7'h15 == total_offset_16[6:0] ? phv_data_21 : _GEN_863; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_865 = 7'h16 == total_offset_16[6:0] ? phv_data_22 : _GEN_864; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_866 = 7'h17 == total_offset_16[6:0] ? phv_data_23 : _GEN_865; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_867 = 7'h18 == total_offset_16[6:0] ? phv_data_24 : _GEN_866; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_868 = 7'h19 == total_offset_16[6:0] ? phv_data_25 : _GEN_867; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_869 = 7'h1a == total_offset_16[6:0] ? phv_data_26 : _GEN_868; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_870 = 7'h1b == total_offset_16[6:0] ? phv_data_27 : _GEN_869; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_871 = 7'h1c == total_offset_16[6:0] ? phv_data_28 : _GEN_870; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_872 = 7'h1d == total_offset_16[6:0] ? phv_data_29 : _GEN_871; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_873 = 7'h1e == total_offset_16[6:0] ? phv_data_30 : _GEN_872; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_874 = 7'h1f == total_offset_16[6:0] ? phv_data_31 : _GEN_873; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_875 = 7'h20 == total_offset_16[6:0] ? phv_data_32 : _GEN_874; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_876 = 7'h21 == total_offset_16[6:0] ? phv_data_33 : _GEN_875; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_877 = 7'h22 == total_offset_16[6:0] ? phv_data_34 : _GEN_876; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_878 = 7'h23 == total_offset_16[6:0] ? phv_data_35 : _GEN_877; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_879 = 7'h24 == total_offset_16[6:0] ? phv_data_36 : _GEN_878; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_880 = 7'h25 == total_offset_16[6:0] ? phv_data_37 : _GEN_879; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_881 = 7'h26 == total_offset_16[6:0] ? phv_data_38 : _GEN_880; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_882 = 7'h27 == total_offset_16[6:0] ? phv_data_39 : _GEN_881; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_883 = 7'h28 == total_offset_16[6:0] ? phv_data_40 : _GEN_882; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_884 = 7'h29 == total_offset_16[6:0] ? phv_data_41 : _GEN_883; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_885 = 7'h2a == total_offset_16[6:0] ? phv_data_42 : _GEN_884; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_886 = 7'h2b == total_offset_16[6:0] ? phv_data_43 : _GEN_885; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_887 = 7'h2c == total_offset_16[6:0] ? phv_data_44 : _GEN_886; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_888 = 7'h2d == total_offset_16[6:0] ? phv_data_45 : _GEN_887; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_889 = 7'h2e == total_offset_16[6:0] ? phv_data_46 : _GEN_888; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_890 = 7'h2f == total_offset_16[6:0] ? phv_data_47 : _GEN_889; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_891 = 7'h30 == total_offset_16[6:0] ? phv_data_48 : _GEN_890; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_892 = 7'h31 == total_offset_16[6:0] ? phv_data_49 : _GEN_891; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_893 = 7'h32 == total_offset_16[6:0] ? phv_data_50 : _GEN_892; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_894 = 7'h33 == total_offset_16[6:0] ? phv_data_51 : _GEN_893; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_895 = 7'h34 == total_offset_16[6:0] ? phv_data_52 : _GEN_894; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_896 = 7'h35 == total_offset_16[6:0] ? phv_data_53 : _GEN_895; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_897 = 7'h36 == total_offset_16[6:0] ? phv_data_54 : _GEN_896; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_898 = 7'h37 == total_offset_16[6:0] ? phv_data_55 : _GEN_897; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_899 = 7'h38 == total_offset_16[6:0] ? phv_data_56 : _GEN_898; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_900 = 7'h39 == total_offset_16[6:0] ? phv_data_57 : _GEN_899; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_901 = 7'h3a == total_offset_16[6:0] ? phv_data_58 : _GEN_900; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_902 = 7'h3b == total_offset_16[6:0] ? phv_data_59 : _GEN_901; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_903 = 7'h3c == total_offset_16[6:0] ? phv_data_60 : _GEN_902; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_904 = 7'h3d == total_offset_16[6:0] ? phv_data_61 : _GEN_903; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_905 = 7'h3e == total_offset_16[6:0] ? phv_data_62 : _GEN_904; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_906 = 7'h3f == total_offset_16[6:0] ? phv_data_63 : _GEN_905; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_907 = 7'h40 == total_offset_16[6:0] ? phv_data_64 : _GEN_906; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_908 = 7'h41 == total_offset_16[6:0] ? phv_data_65 : _GEN_907; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_909 = 7'h42 == total_offset_16[6:0] ? phv_data_66 : _GEN_908; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_910 = 7'h43 == total_offset_16[6:0] ? phv_data_67 : _GEN_909; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_911 = 7'h44 == total_offset_16[6:0] ? phv_data_68 : _GEN_910; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_912 = 7'h45 == total_offset_16[6:0] ? phv_data_69 : _GEN_911; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_913 = 7'h46 == total_offset_16[6:0] ? phv_data_70 : _GEN_912; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_914 = 7'h47 == total_offset_16[6:0] ? phv_data_71 : _GEN_913; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_915 = 7'h48 == total_offset_16[6:0] ? phv_data_72 : _GEN_914; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_916 = 7'h49 == total_offset_16[6:0] ? phv_data_73 : _GEN_915; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_917 = 7'h4a == total_offset_16[6:0] ? phv_data_74 : _GEN_916; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_918 = 7'h4b == total_offset_16[6:0] ? phv_data_75 : _GEN_917; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_919 = 7'h4c == total_offset_16[6:0] ? phv_data_76 : _GEN_918; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_920 = 7'h4d == total_offset_16[6:0] ? phv_data_77 : _GEN_919; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_921 = 7'h4e == total_offset_16[6:0] ? phv_data_78 : _GEN_920; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_922 = 7'h4f == total_offset_16[6:0] ? phv_data_79 : _GEN_921; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_923 = 7'h50 == total_offset_16[6:0] ? phv_data_80 : _GEN_922; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_924 = 7'h51 == total_offset_16[6:0] ? phv_data_81 : _GEN_923; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_925 = 7'h52 == total_offset_16[6:0] ? phv_data_82 : _GEN_924; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_926 = 7'h53 == total_offset_16[6:0] ? phv_data_83 : _GEN_925; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_927 = 7'h54 == total_offset_16[6:0] ? phv_data_84 : _GEN_926; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_928 = 7'h55 == total_offset_16[6:0] ? phv_data_85 : _GEN_927; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_929 = 7'h56 == total_offset_16[6:0] ? phv_data_86 : _GEN_928; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_930 = 7'h57 == total_offset_16[6:0] ? phv_data_87 : _GEN_929; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_931 = 7'h58 == total_offset_16[6:0] ? phv_data_88 : _GEN_930; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_932 = 7'h59 == total_offset_16[6:0] ? phv_data_89 : _GEN_931; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_933 = 7'h5a == total_offset_16[6:0] ? phv_data_90 : _GEN_932; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_934 = 7'h5b == total_offset_16[6:0] ? phv_data_91 : _GEN_933; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_935 = 7'h5c == total_offset_16[6:0] ? phv_data_92 : _GEN_934; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_936 = 7'h5d == total_offset_16[6:0] ? phv_data_93 : _GEN_935; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_937 = 7'h5e == total_offset_16[6:0] ? phv_data_94 : _GEN_936; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_938 = 7'h5f == total_offset_16[6:0] ? phv_data_95 : _GEN_937; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes_2_0 = 8'h0 < length_1 ? _GEN_938 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_17 = offset_1 + 8'h1; // @[executor.scala 158:57]
  wire [7:0] _GEN_941 = 7'h1 == total_offset_17[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_942 = 7'h2 == total_offset_17[6:0] ? phv_data_2 : _GEN_941; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_943 = 7'h3 == total_offset_17[6:0] ? phv_data_3 : _GEN_942; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_944 = 7'h4 == total_offset_17[6:0] ? phv_data_4 : _GEN_943; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_945 = 7'h5 == total_offset_17[6:0] ? phv_data_5 : _GEN_944; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_946 = 7'h6 == total_offset_17[6:0] ? phv_data_6 : _GEN_945; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_947 = 7'h7 == total_offset_17[6:0] ? phv_data_7 : _GEN_946; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_948 = 7'h8 == total_offset_17[6:0] ? phv_data_8 : _GEN_947; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_949 = 7'h9 == total_offset_17[6:0] ? phv_data_9 : _GEN_948; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_950 = 7'ha == total_offset_17[6:0] ? phv_data_10 : _GEN_949; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_951 = 7'hb == total_offset_17[6:0] ? phv_data_11 : _GEN_950; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_952 = 7'hc == total_offset_17[6:0] ? phv_data_12 : _GEN_951; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_953 = 7'hd == total_offset_17[6:0] ? phv_data_13 : _GEN_952; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_954 = 7'he == total_offset_17[6:0] ? phv_data_14 : _GEN_953; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_955 = 7'hf == total_offset_17[6:0] ? phv_data_15 : _GEN_954; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_956 = 7'h10 == total_offset_17[6:0] ? phv_data_16 : _GEN_955; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_957 = 7'h11 == total_offset_17[6:0] ? phv_data_17 : _GEN_956; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_958 = 7'h12 == total_offset_17[6:0] ? phv_data_18 : _GEN_957; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_959 = 7'h13 == total_offset_17[6:0] ? phv_data_19 : _GEN_958; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_960 = 7'h14 == total_offset_17[6:0] ? phv_data_20 : _GEN_959; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_961 = 7'h15 == total_offset_17[6:0] ? phv_data_21 : _GEN_960; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_962 = 7'h16 == total_offset_17[6:0] ? phv_data_22 : _GEN_961; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_963 = 7'h17 == total_offset_17[6:0] ? phv_data_23 : _GEN_962; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_964 = 7'h18 == total_offset_17[6:0] ? phv_data_24 : _GEN_963; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_965 = 7'h19 == total_offset_17[6:0] ? phv_data_25 : _GEN_964; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_966 = 7'h1a == total_offset_17[6:0] ? phv_data_26 : _GEN_965; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_967 = 7'h1b == total_offset_17[6:0] ? phv_data_27 : _GEN_966; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_968 = 7'h1c == total_offset_17[6:0] ? phv_data_28 : _GEN_967; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_969 = 7'h1d == total_offset_17[6:0] ? phv_data_29 : _GEN_968; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_970 = 7'h1e == total_offset_17[6:0] ? phv_data_30 : _GEN_969; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_971 = 7'h1f == total_offset_17[6:0] ? phv_data_31 : _GEN_970; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_972 = 7'h20 == total_offset_17[6:0] ? phv_data_32 : _GEN_971; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_973 = 7'h21 == total_offset_17[6:0] ? phv_data_33 : _GEN_972; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_974 = 7'h22 == total_offset_17[6:0] ? phv_data_34 : _GEN_973; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_975 = 7'h23 == total_offset_17[6:0] ? phv_data_35 : _GEN_974; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_976 = 7'h24 == total_offset_17[6:0] ? phv_data_36 : _GEN_975; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_977 = 7'h25 == total_offset_17[6:0] ? phv_data_37 : _GEN_976; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_978 = 7'h26 == total_offset_17[6:0] ? phv_data_38 : _GEN_977; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_979 = 7'h27 == total_offset_17[6:0] ? phv_data_39 : _GEN_978; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_980 = 7'h28 == total_offset_17[6:0] ? phv_data_40 : _GEN_979; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_981 = 7'h29 == total_offset_17[6:0] ? phv_data_41 : _GEN_980; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_982 = 7'h2a == total_offset_17[6:0] ? phv_data_42 : _GEN_981; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_983 = 7'h2b == total_offset_17[6:0] ? phv_data_43 : _GEN_982; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_984 = 7'h2c == total_offset_17[6:0] ? phv_data_44 : _GEN_983; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_985 = 7'h2d == total_offset_17[6:0] ? phv_data_45 : _GEN_984; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_986 = 7'h2e == total_offset_17[6:0] ? phv_data_46 : _GEN_985; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_987 = 7'h2f == total_offset_17[6:0] ? phv_data_47 : _GEN_986; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_988 = 7'h30 == total_offset_17[6:0] ? phv_data_48 : _GEN_987; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_989 = 7'h31 == total_offset_17[6:0] ? phv_data_49 : _GEN_988; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_990 = 7'h32 == total_offset_17[6:0] ? phv_data_50 : _GEN_989; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_991 = 7'h33 == total_offset_17[6:0] ? phv_data_51 : _GEN_990; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_992 = 7'h34 == total_offset_17[6:0] ? phv_data_52 : _GEN_991; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_993 = 7'h35 == total_offset_17[6:0] ? phv_data_53 : _GEN_992; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_994 = 7'h36 == total_offset_17[6:0] ? phv_data_54 : _GEN_993; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_995 = 7'h37 == total_offset_17[6:0] ? phv_data_55 : _GEN_994; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_996 = 7'h38 == total_offset_17[6:0] ? phv_data_56 : _GEN_995; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_997 = 7'h39 == total_offset_17[6:0] ? phv_data_57 : _GEN_996; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_998 = 7'h3a == total_offset_17[6:0] ? phv_data_58 : _GEN_997; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_999 = 7'h3b == total_offset_17[6:0] ? phv_data_59 : _GEN_998; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1000 = 7'h3c == total_offset_17[6:0] ? phv_data_60 : _GEN_999; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1001 = 7'h3d == total_offset_17[6:0] ? phv_data_61 : _GEN_1000; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1002 = 7'h3e == total_offset_17[6:0] ? phv_data_62 : _GEN_1001; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1003 = 7'h3f == total_offset_17[6:0] ? phv_data_63 : _GEN_1002; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1004 = 7'h40 == total_offset_17[6:0] ? phv_data_64 : _GEN_1003; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1005 = 7'h41 == total_offset_17[6:0] ? phv_data_65 : _GEN_1004; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1006 = 7'h42 == total_offset_17[6:0] ? phv_data_66 : _GEN_1005; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1007 = 7'h43 == total_offset_17[6:0] ? phv_data_67 : _GEN_1006; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1008 = 7'h44 == total_offset_17[6:0] ? phv_data_68 : _GEN_1007; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1009 = 7'h45 == total_offset_17[6:0] ? phv_data_69 : _GEN_1008; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1010 = 7'h46 == total_offset_17[6:0] ? phv_data_70 : _GEN_1009; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1011 = 7'h47 == total_offset_17[6:0] ? phv_data_71 : _GEN_1010; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1012 = 7'h48 == total_offset_17[6:0] ? phv_data_72 : _GEN_1011; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1013 = 7'h49 == total_offset_17[6:0] ? phv_data_73 : _GEN_1012; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1014 = 7'h4a == total_offset_17[6:0] ? phv_data_74 : _GEN_1013; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1015 = 7'h4b == total_offset_17[6:0] ? phv_data_75 : _GEN_1014; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1016 = 7'h4c == total_offset_17[6:0] ? phv_data_76 : _GEN_1015; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1017 = 7'h4d == total_offset_17[6:0] ? phv_data_77 : _GEN_1016; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1018 = 7'h4e == total_offset_17[6:0] ? phv_data_78 : _GEN_1017; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1019 = 7'h4f == total_offset_17[6:0] ? phv_data_79 : _GEN_1018; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1020 = 7'h50 == total_offset_17[6:0] ? phv_data_80 : _GEN_1019; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1021 = 7'h51 == total_offset_17[6:0] ? phv_data_81 : _GEN_1020; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1022 = 7'h52 == total_offset_17[6:0] ? phv_data_82 : _GEN_1021; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1023 = 7'h53 == total_offset_17[6:0] ? phv_data_83 : _GEN_1022; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1024 = 7'h54 == total_offset_17[6:0] ? phv_data_84 : _GEN_1023; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1025 = 7'h55 == total_offset_17[6:0] ? phv_data_85 : _GEN_1024; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1026 = 7'h56 == total_offset_17[6:0] ? phv_data_86 : _GEN_1025; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1027 = 7'h57 == total_offset_17[6:0] ? phv_data_87 : _GEN_1026; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1028 = 7'h58 == total_offset_17[6:0] ? phv_data_88 : _GEN_1027; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1029 = 7'h59 == total_offset_17[6:0] ? phv_data_89 : _GEN_1028; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1030 = 7'h5a == total_offset_17[6:0] ? phv_data_90 : _GEN_1029; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1031 = 7'h5b == total_offset_17[6:0] ? phv_data_91 : _GEN_1030; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1032 = 7'h5c == total_offset_17[6:0] ? phv_data_92 : _GEN_1031; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1033 = 7'h5d == total_offset_17[6:0] ? phv_data_93 : _GEN_1032; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1034 = 7'h5e == total_offset_17[6:0] ? phv_data_94 : _GEN_1033; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1035 = 7'h5f == total_offset_17[6:0] ? phv_data_95 : _GEN_1034; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes_2_1 = 8'h1 < length_1 ? _GEN_1035 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_18 = offset_1 + 8'h2; // @[executor.scala 158:57]
  wire [7:0] _GEN_1038 = 7'h1 == total_offset_18[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1039 = 7'h2 == total_offset_18[6:0] ? phv_data_2 : _GEN_1038; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1040 = 7'h3 == total_offset_18[6:0] ? phv_data_3 : _GEN_1039; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1041 = 7'h4 == total_offset_18[6:0] ? phv_data_4 : _GEN_1040; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1042 = 7'h5 == total_offset_18[6:0] ? phv_data_5 : _GEN_1041; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1043 = 7'h6 == total_offset_18[6:0] ? phv_data_6 : _GEN_1042; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1044 = 7'h7 == total_offset_18[6:0] ? phv_data_7 : _GEN_1043; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1045 = 7'h8 == total_offset_18[6:0] ? phv_data_8 : _GEN_1044; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1046 = 7'h9 == total_offset_18[6:0] ? phv_data_9 : _GEN_1045; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1047 = 7'ha == total_offset_18[6:0] ? phv_data_10 : _GEN_1046; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1048 = 7'hb == total_offset_18[6:0] ? phv_data_11 : _GEN_1047; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1049 = 7'hc == total_offset_18[6:0] ? phv_data_12 : _GEN_1048; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1050 = 7'hd == total_offset_18[6:0] ? phv_data_13 : _GEN_1049; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1051 = 7'he == total_offset_18[6:0] ? phv_data_14 : _GEN_1050; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1052 = 7'hf == total_offset_18[6:0] ? phv_data_15 : _GEN_1051; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1053 = 7'h10 == total_offset_18[6:0] ? phv_data_16 : _GEN_1052; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1054 = 7'h11 == total_offset_18[6:0] ? phv_data_17 : _GEN_1053; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1055 = 7'h12 == total_offset_18[6:0] ? phv_data_18 : _GEN_1054; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1056 = 7'h13 == total_offset_18[6:0] ? phv_data_19 : _GEN_1055; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1057 = 7'h14 == total_offset_18[6:0] ? phv_data_20 : _GEN_1056; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1058 = 7'h15 == total_offset_18[6:0] ? phv_data_21 : _GEN_1057; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1059 = 7'h16 == total_offset_18[6:0] ? phv_data_22 : _GEN_1058; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1060 = 7'h17 == total_offset_18[6:0] ? phv_data_23 : _GEN_1059; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1061 = 7'h18 == total_offset_18[6:0] ? phv_data_24 : _GEN_1060; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1062 = 7'h19 == total_offset_18[6:0] ? phv_data_25 : _GEN_1061; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1063 = 7'h1a == total_offset_18[6:0] ? phv_data_26 : _GEN_1062; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1064 = 7'h1b == total_offset_18[6:0] ? phv_data_27 : _GEN_1063; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1065 = 7'h1c == total_offset_18[6:0] ? phv_data_28 : _GEN_1064; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1066 = 7'h1d == total_offset_18[6:0] ? phv_data_29 : _GEN_1065; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1067 = 7'h1e == total_offset_18[6:0] ? phv_data_30 : _GEN_1066; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1068 = 7'h1f == total_offset_18[6:0] ? phv_data_31 : _GEN_1067; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1069 = 7'h20 == total_offset_18[6:0] ? phv_data_32 : _GEN_1068; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1070 = 7'h21 == total_offset_18[6:0] ? phv_data_33 : _GEN_1069; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1071 = 7'h22 == total_offset_18[6:0] ? phv_data_34 : _GEN_1070; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1072 = 7'h23 == total_offset_18[6:0] ? phv_data_35 : _GEN_1071; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1073 = 7'h24 == total_offset_18[6:0] ? phv_data_36 : _GEN_1072; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1074 = 7'h25 == total_offset_18[6:0] ? phv_data_37 : _GEN_1073; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1075 = 7'h26 == total_offset_18[6:0] ? phv_data_38 : _GEN_1074; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1076 = 7'h27 == total_offset_18[6:0] ? phv_data_39 : _GEN_1075; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1077 = 7'h28 == total_offset_18[6:0] ? phv_data_40 : _GEN_1076; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1078 = 7'h29 == total_offset_18[6:0] ? phv_data_41 : _GEN_1077; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1079 = 7'h2a == total_offset_18[6:0] ? phv_data_42 : _GEN_1078; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1080 = 7'h2b == total_offset_18[6:0] ? phv_data_43 : _GEN_1079; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1081 = 7'h2c == total_offset_18[6:0] ? phv_data_44 : _GEN_1080; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1082 = 7'h2d == total_offset_18[6:0] ? phv_data_45 : _GEN_1081; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1083 = 7'h2e == total_offset_18[6:0] ? phv_data_46 : _GEN_1082; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1084 = 7'h2f == total_offset_18[6:0] ? phv_data_47 : _GEN_1083; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1085 = 7'h30 == total_offset_18[6:0] ? phv_data_48 : _GEN_1084; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1086 = 7'h31 == total_offset_18[6:0] ? phv_data_49 : _GEN_1085; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1087 = 7'h32 == total_offset_18[6:0] ? phv_data_50 : _GEN_1086; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1088 = 7'h33 == total_offset_18[6:0] ? phv_data_51 : _GEN_1087; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1089 = 7'h34 == total_offset_18[6:0] ? phv_data_52 : _GEN_1088; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1090 = 7'h35 == total_offset_18[6:0] ? phv_data_53 : _GEN_1089; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1091 = 7'h36 == total_offset_18[6:0] ? phv_data_54 : _GEN_1090; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1092 = 7'h37 == total_offset_18[6:0] ? phv_data_55 : _GEN_1091; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1093 = 7'h38 == total_offset_18[6:0] ? phv_data_56 : _GEN_1092; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1094 = 7'h39 == total_offset_18[6:0] ? phv_data_57 : _GEN_1093; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1095 = 7'h3a == total_offset_18[6:0] ? phv_data_58 : _GEN_1094; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1096 = 7'h3b == total_offset_18[6:0] ? phv_data_59 : _GEN_1095; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1097 = 7'h3c == total_offset_18[6:0] ? phv_data_60 : _GEN_1096; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1098 = 7'h3d == total_offset_18[6:0] ? phv_data_61 : _GEN_1097; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1099 = 7'h3e == total_offset_18[6:0] ? phv_data_62 : _GEN_1098; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1100 = 7'h3f == total_offset_18[6:0] ? phv_data_63 : _GEN_1099; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1101 = 7'h40 == total_offset_18[6:0] ? phv_data_64 : _GEN_1100; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1102 = 7'h41 == total_offset_18[6:0] ? phv_data_65 : _GEN_1101; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1103 = 7'h42 == total_offset_18[6:0] ? phv_data_66 : _GEN_1102; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1104 = 7'h43 == total_offset_18[6:0] ? phv_data_67 : _GEN_1103; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1105 = 7'h44 == total_offset_18[6:0] ? phv_data_68 : _GEN_1104; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1106 = 7'h45 == total_offset_18[6:0] ? phv_data_69 : _GEN_1105; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1107 = 7'h46 == total_offset_18[6:0] ? phv_data_70 : _GEN_1106; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1108 = 7'h47 == total_offset_18[6:0] ? phv_data_71 : _GEN_1107; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1109 = 7'h48 == total_offset_18[6:0] ? phv_data_72 : _GEN_1108; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1110 = 7'h49 == total_offset_18[6:0] ? phv_data_73 : _GEN_1109; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1111 = 7'h4a == total_offset_18[6:0] ? phv_data_74 : _GEN_1110; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1112 = 7'h4b == total_offset_18[6:0] ? phv_data_75 : _GEN_1111; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1113 = 7'h4c == total_offset_18[6:0] ? phv_data_76 : _GEN_1112; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1114 = 7'h4d == total_offset_18[6:0] ? phv_data_77 : _GEN_1113; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1115 = 7'h4e == total_offset_18[6:0] ? phv_data_78 : _GEN_1114; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1116 = 7'h4f == total_offset_18[6:0] ? phv_data_79 : _GEN_1115; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1117 = 7'h50 == total_offset_18[6:0] ? phv_data_80 : _GEN_1116; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1118 = 7'h51 == total_offset_18[6:0] ? phv_data_81 : _GEN_1117; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1119 = 7'h52 == total_offset_18[6:0] ? phv_data_82 : _GEN_1118; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1120 = 7'h53 == total_offset_18[6:0] ? phv_data_83 : _GEN_1119; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1121 = 7'h54 == total_offset_18[6:0] ? phv_data_84 : _GEN_1120; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1122 = 7'h55 == total_offset_18[6:0] ? phv_data_85 : _GEN_1121; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1123 = 7'h56 == total_offset_18[6:0] ? phv_data_86 : _GEN_1122; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1124 = 7'h57 == total_offset_18[6:0] ? phv_data_87 : _GEN_1123; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1125 = 7'h58 == total_offset_18[6:0] ? phv_data_88 : _GEN_1124; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1126 = 7'h59 == total_offset_18[6:0] ? phv_data_89 : _GEN_1125; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1127 = 7'h5a == total_offset_18[6:0] ? phv_data_90 : _GEN_1126; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1128 = 7'h5b == total_offset_18[6:0] ? phv_data_91 : _GEN_1127; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1129 = 7'h5c == total_offset_18[6:0] ? phv_data_92 : _GEN_1128; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1130 = 7'h5d == total_offset_18[6:0] ? phv_data_93 : _GEN_1129; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1131 = 7'h5e == total_offset_18[6:0] ? phv_data_94 : _GEN_1130; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1132 = 7'h5f == total_offset_18[6:0] ? phv_data_95 : _GEN_1131; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes_2_2 = 8'h2 < length_1 ? _GEN_1132 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_19 = offset_1 + 8'h3; // @[executor.scala 158:57]
  wire [7:0] _GEN_1135 = 7'h1 == total_offset_19[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1136 = 7'h2 == total_offset_19[6:0] ? phv_data_2 : _GEN_1135; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1137 = 7'h3 == total_offset_19[6:0] ? phv_data_3 : _GEN_1136; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1138 = 7'h4 == total_offset_19[6:0] ? phv_data_4 : _GEN_1137; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1139 = 7'h5 == total_offset_19[6:0] ? phv_data_5 : _GEN_1138; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1140 = 7'h6 == total_offset_19[6:0] ? phv_data_6 : _GEN_1139; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1141 = 7'h7 == total_offset_19[6:0] ? phv_data_7 : _GEN_1140; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1142 = 7'h8 == total_offset_19[6:0] ? phv_data_8 : _GEN_1141; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1143 = 7'h9 == total_offset_19[6:0] ? phv_data_9 : _GEN_1142; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1144 = 7'ha == total_offset_19[6:0] ? phv_data_10 : _GEN_1143; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1145 = 7'hb == total_offset_19[6:0] ? phv_data_11 : _GEN_1144; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1146 = 7'hc == total_offset_19[6:0] ? phv_data_12 : _GEN_1145; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1147 = 7'hd == total_offset_19[6:0] ? phv_data_13 : _GEN_1146; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1148 = 7'he == total_offset_19[6:0] ? phv_data_14 : _GEN_1147; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1149 = 7'hf == total_offset_19[6:0] ? phv_data_15 : _GEN_1148; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1150 = 7'h10 == total_offset_19[6:0] ? phv_data_16 : _GEN_1149; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1151 = 7'h11 == total_offset_19[6:0] ? phv_data_17 : _GEN_1150; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1152 = 7'h12 == total_offset_19[6:0] ? phv_data_18 : _GEN_1151; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1153 = 7'h13 == total_offset_19[6:0] ? phv_data_19 : _GEN_1152; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1154 = 7'h14 == total_offset_19[6:0] ? phv_data_20 : _GEN_1153; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1155 = 7'h15 == total_offset_19[6:0] ? phv_data_21 : _GEN_1154; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1156 = 7'h16 == total_offset_19[6:0] ? phv_data_22 : _GEN_1155; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1157 = 7'h17 == total_offset_19[6:0] ? phv_data_23 : _GEN_1156; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1158 = 7'h18 == total_offset_19[6:0] ? phv_data_24 : _GEN_1157; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1159 = 7'h19 == total_offset_19[6:0] ? phv_data_25 : _GEN_1158; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1160 = 7'h1a == total_offset_19[6:0] ? phv_data_26 : _GEN_1159; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1161 = 7'h1b == total_offset_19[6:0] ? phv_data_27 : _GEN_1160; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1162 = 7'h1c == total_offset_19[6:0] ? phv_data_28 : _GEN_1161; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1163 = 7'h1d == total_offset_19[6:0] ? phv_data_29 : _GEN_1162; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1164 = 7'h1e == total_offset_19[6:0] ? phv_data_30 : _GEN_1163; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1165 = 7'h1f == total_offset_19[6:0] ? phv_data_31 : _GEN_1164; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1166 = 7'h20 == total_offset_19[6:0] ? phv_data_32 : _GEN_1165; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1167 = 7'h21 == total_offset_19[6:0] ? phv_data_33 : _GEN_1166; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1168 = 7'h22 == total_offset_19[6:0] ? phv_data_34 : _GEN_1167; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1169 = 7'h23 == total_offset_19[6:0] ? phv_data_35 : _GEN_1168; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1170 = 7'h24 == total_offset_19[6:0] ? phv_data_36 : _GEN_1169; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1171 = 7'h25 == total_offset_19[6:0] ? phv_data_37 : _GEN_1170; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1172 = 7'h26 == total_offset_19[6:0] ? phv_data_38 : _GEN_1171; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1173 = 7'h27 == total_offset_19[6:0] ? phv_data_39 : _GEN_1172; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1174 = 7'h28 == total_offset_19[6:0] ? phv_data_40 : _GEN_1173; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1175 = 7'h29 == total_offset_19[6:0] ? phv_data_41 : _GEN_1174; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1176 = 7'h2a == total_offset_19[6:0] ? phv_data_42 : _GEN_1175; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1177 = 7'h2b == total_offset_19[6:0] ? phv_data_43 : _GEN_1176; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1178 = 7'h2c == total_offset_19[6:0] ? phv_data_44 : _GEN_1177; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1179 = 7'h2d == total_offset_19[6:0] ? phv_data_45 : _GEN_1178; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1180 = 7'h2e == total_offset_19[6:0] ? phv_data_46 : _GEN_1179; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1181 = 7'h2f == total_offset_19[6:0] ? phv_data_47 : _GEN_1180; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1182 = 7'h30 == total_offset_19[6:0] ? phv_data_48 : _GEN_1181; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1183 = 7'h31 == total_offset_19[6:0] ? phv_data_49 : _GEN_1182; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1184 = 7'h32 == total_offset_19[6:0] ? phv_data_50 : _GEN_1183; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1185 = 7'h33 == total_offset_19[6:0] ? phv_data_51 : _GEN_1184; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1186 = 7'h34 == total_offset_19[6:0] ? phv_data_52 : _GEN_1185; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1187 = 7'h35 == total_offset_19[6:0] ? phv_data_53 : _GEN_1186; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1188 = 7'h36 == total_offset_19[6:0] ? phv_data_54 : _GEN_1187; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1189 = 7'h37 == total_offset_19[6:0] ? phv_data_55 : _GEN_1188; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1190 = 7'h38 == total_offset_19[6:0] ? phv_data_56 : _GEN_1189; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1191 = 7'h39 == total_offset_19[6:0] ? phv_data_57 : _GEN_1190; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1192 = 7'h3a == total_offset_19[6:0] ? phv_data_58 : _GEN_1191; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1193 = 7'h3b == total_offset_19[6:0] ? phv_data_59 : _GEN_1192; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1194 = 7'h3c == total_offset_19[6:0] ? phv_data_60 : _GEN_1193; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1195 = 7'h3d == total_offset_19[6:0] ? phv_data_61 : _GEN_1194; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1196 = 7'h3e == total_offset_19[6:0] ? phv_data_62 : _GEN_1195; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1197 = 7'h3f == total_offset_19[6:0] ? phv_data_63 : _GEN_1196; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1198 = 7'h40 == total_offset_19[6:0] ? phv_data_64 : _GEN_1197; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1199 = 7'h41 == total_offset_19[6:0] ? phv_data_65 : _GEN_1198; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1200 = 7'h42 == total_offset_19[6:0] ? phv_data_66 : _GEN_1199; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1201 = 7'h43 == total_offset_19[6:0] ? phv_data_67 : _GEN_1200; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1202 = 7'h44 == total_offset_19[6:0] ? phv_data_68 : _GEN_1201; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1203 = 7'h45 == total_offset_19[6:0] ? phv_data_69 : _GEN_1202; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1204 = 7'h46 == total_offset_19[6:0] ? phv_data_70 : _GEN_1203; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1205 = 7'h47 == total_offset_19[6:0] ? phv_data_71 : _GEN_1204; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1206 = 7'h48 == total_offset_19[6:0] ? phv_data_72 : _GEN_1205; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1207 = 7'h49 == total_offset_19[6:0] ? phv_data_73 : _GEN_1206; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1208 = 7'h4a == total_offset_19[6:0] ? phv_data_74 : _GEN_1207; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1209 = 7'h4b == total_offset_19[6:0] ? phv_data_75 : _GEN_1208; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1210 = 7'h4c == total_offset_19[6:0] ? phv_data_76 : _GEN_1209; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1211 = 7'h4d == total_offset_19[6:0] ? phv_data_77 : _GEN_1210; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1212 = 7'h4e == total_offset_19[6:0] ? phv_data_78 : _GEN_1211; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1213 = 7'h4f == total_offset_19[6:0] ? phv_data_79 : _GEN_1212; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1214 = 7'h50 == total_offset_19[6:0] ? phv_data_80 : _GEN_1213; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1215 = 7'h51 == total_offset_19[6:0] ? phv_data_81 : _GEN_1214; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1216 = 7'h52 == total_offset_19[6:0] ? phv_data_82 : _GEN_1215; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1217 = 7'h53 == total_offset_19[6:0] ? phv_data_83 : _GEN_1216; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1218 = 7'h54 == total_offset_19[6:0] ? phv_data_84 : _GEN_1217; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1219 = 7'h55 == total_offset_19[6:0] ? phv_data_85 : _GEN_1218; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1220 = 7'h56 == total_offset_19[6:0] ? phv_data_86 : _GEN_1219; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1221 = 7'h57 == total_offset_19[6:0] ? phv_data_87 : _GEN_1220; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1222 = 7'h58 == total_offset_19[6:0] ? phv_data_88 : _GEN_1221; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1223 = 7'h59 == total_offset_19[6:0] ? phv_data_89 : _GEN_1222; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1224 = 7'h5a == total_offset_19[6:0] ? phv_data_90 : _GEN_1223; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1225 = 7'h5b == total_offset_19[6:0] ? phv_data_91 : _GEN_1224; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1226 = 7'h5c == total_offset_19[6:0] ? phv_data_92 : _GEN_1225; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1227 = 7'h5d == total_offset_19[6:0] ? phv_data_93 : _GEN_1226; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1228 = 7'h5e == total_offset_19[6:0] ? phv_data_94 : _GEN_1227; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1229 = 7'h5f == total_offset_19[6:0] ? phv_data_95 : _GEN_1228; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes_2_3 = 8'h3 < length_1 ? _GEN_1229 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_20 = offset_1 + 8'h4; // @[executor.scala 158:57]
  wire [7:0] _GEN_1232 = 7'h1 == total_offset_20[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1233 = 7'h2 == total_offset_20[6:0] ? phv_data_2 : _GEN_1232; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1234 = 7'h3 == total_offset_20[6:0] ? phv_data_3 : _GEN_1233; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1235 = 7'h4 == total_offset_20[6:0] ? phv_data_4 : _GEN_1234; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1236 = 7'h5 == total_offset_20[6:0] ? phv_data_5 : _GEN_1235; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1237 = 7'h6 == total_offset_20[6:0] ? phv_data_6 : _GEN_1236; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1238 = 7'h7 == total_offset_20[6:0] ? phv_data_7 : _GEN_1237; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1239 = 7'h8 == total_offset_20[6:0] ? phv_data_8 : _GEN_1238; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1240 = 7'h9 == total_offset_20[6:0] ? phv_data_9 : _GEN_1239; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1241 = 7'ha == total_offset_20[6:0] ? phv_data_10 : _GEN_1240; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1242 = 7'hb == total_offset_20[6:0] ? phv_data_11 : _GEN_1241; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1243 = 7'hc == total_offset_20[6:0] ? phv_data_12 : _GEN_1242; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1244 = 7'hd == total_offset_20[6:0] ? phv_data_13 : _GEN_1243; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1245 = 7'he == total_offset_20[6:0] ? phv_data_14 : _GEN_1244; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1246 = 7'hf == total_offset_20[6:0] ? phv_data_15 : _GEN_1245; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1247 = 7'h10 == total_offset_20[6:0] ? phv_data_16 : _GEN_1246; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1248 = 7'h11 == total_offset_20[6:0] ? phv_data_17 : _GEN_1247; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1249 = 7'h12 == total_offset_20[6:0] ? phv_data_18 : _GEN_1248; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1250 = 7'h13 == total_offset_20[6:0] ? phv_data_19 : _GEN_1249; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1251 = 7'h14 == total_offset_20[6:0] ? phv_data_20 : _GEN_1250; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1252 = 7'h15 == total_offset_20[6:0] ? phv_data_21 : _GEN_1251; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1253 = 7'h16 == total_offset_20[6:0] ? phv_data_22 : _GEN_1252; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1254 = 7'h17 == total_offset_20[6:0] ? phv_data_23 : _GEN_1253; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1255 = 7'h18 == total_offset_20[6:0] ? phv_data_24 : _GEN_1254; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1256 = 7'h19 == total_offset_20[6:0] ? phv_data_25 : _GEN_1255; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1257 = 7'h1a == total_offset_20[6:0] ? phv_data_26 : _GEN_1256; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1258 = 7'h1b == total_offset_20[6:0] ? phv_data_27 : _GEN_1257; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1259 = 7'h1c == total_offset_20[6:0] ? phv_data_28 : _GEN_1258; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1260 = 7'h1d == total_offset_20[6:0] ? phv_data_29 : _GEN_1259; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1261 = 7'h1e == total_offset_20[6:0] ? phv_data_30 : _GEN_1260; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1262 = 7'h1f == total_offset_20[6:0] ? phv_data_31 : _GEN_1261; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1263 = 7'h20 == total_offset_20[6:0] ? phv_data_32 : _GEN_1262; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1264 = 7'h21 == total_offset_20[6:0] ? phv_data_33 : _GEN_1263; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1265 = 7'h22 == total_offset_20[6:0] ? phv_data_34 : _GEN_1264; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1266 = 7'h23 == total_offset_20[6:0] ? phv_data_35 : _GEN_1265; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1267 = 7'h24 == total_offset_20[6:0] ? phv_data_36 : _GEN_1266; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1268 = 7'h25 == total_offset_20[6:0] ? phv_data_37 : _GEN_1267; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1269 = 7'h26 == total_offset_20[6:0] ? phv_data_38 : _GEN_1268; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1270 = 7'h27 == total_offset_20[6:0] ? phv_data_39 : _GEN_1269; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1271 = 7'h28 == total_offset_20[6:0] ? phv_data_40 : _GEN_1270; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1272 = 7'h29 == total_offset_20[6:0] ? phv_data_41 : _GEN_1271; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1273 = 7'h2a == total_offset_20[6:0] ? phv_data_42 : _GEN_1272; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1274 = 7'h2b == total_offset_20[6:0] ? phv_data_43 : _GEN_1273; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1275 = 7'h2c == total_offset_20[6:0] ? phv_data_44 : _GEN_1274; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1276 = 7'h2d == total_offset_20[6:0] ? phv_data_45 : _GEN_1275; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1277 = 7'h2e == total_offset_20[6:0] ? phv_data_46 : _GEN_1276; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1278 = 7'h2f == total_offset_20[6:0] ? phv_data_47 : _GEN_1277; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1279 = 7'h30 == total_offset_20[6:0] ? phv_data_48 : _GEN_1278; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1280 = 7'h31 == total_offset_20[6:0] ? phv_data_49 : _GEN_1279; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1281 = 7'h32 == total_offset_20[6:0] ? phv_data_50 : _GEN_1280; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1282 = 7'h33 == total_offset_20[6:0] ? phv_data_51 : _GEN_1281; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1283 = 7'h34 == total_offset_20[6:0] ? phv_data_52 : _GEN_1282; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1284 = 7'h35 == total_offset_20[6:0] ? phv_data_53 : _GEN_1283; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1285 = 7'h36 == total_offset_20[6:0] ? phv_data_54 : _GEN_1284; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1286 = 7'h37 == total_offset_20[6:0] ? phv_data_55 : _GEN_1285; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1287 = 7'h38 == total_offset_20[6:0] ? phv_data_56 : _GEN_1286; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1288 = 7'h39 == total_offset_20[6:0] ? phv_data_57 : _GEN_1287; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1289 = 7'h3a == total_offset_20[6:0] ? phv_data_58 : _GEN_1288; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1290 = 7'h3b == total_offset_20[6:0] ? phv_data_59 : _GEN_1289; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1291 = 7'h3c == total_offset_20[6:0] ? phv_data_60 : _GEN_1290; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1292 = 7'h3d == total_offset_20[6:0] ? phv_data_61 : _GEN_1291; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1293 = 7'h3e == total_offset_20[6:0] ? phv_data_62 : _GEN_1292; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1294 = 7'h3f == total_offset_20[6:0] ? phv_data_63 : _GEN_1293; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1295 = 7'h40 == total_offset_20[6:0] ? phv_data_64 : _GEN_1294; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1296 = 7'h41 == total_offset_20[6:0] ? phv_data_65 : _GEN_1295; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1297 = 7'h42 == total_offset_20[6:0] ? phv_data_66 : _GEN_1296; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1298 = 7'h43 == total_offset_20[6:0] ? phv_data_67 : _GEN_1297; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1299 = 7'h44 == total_offset_20[6:0] ? phv_data_68 : _GEN_1298; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1300 = 7'h45 == total_offset_20[6:0] ? phv_data_69 : _GEN_1299; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1301 = 7'h46 == total_offset_20[6:0] ? phv_data_70 : _GEN_1300; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1302 = 7'h47 == total_offset_20[6:0] ? phv_data_71 : _GEN_1301; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1303 = 7'h48 == total_offset_20[6:0] ? phv_data_72 : _GEN_1302; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1304 = 7'h49 == total_offset_20[6:0] ? phv_data_73 : _GEN_1303; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1305 = 7'h4a == total_offset_20[6:0] ? phv_data_74 : _GEN_1304; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1306 = 7'h4b == total_offset_20[6:0] ? phv_data_75 : _GEN_1305; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1307 = 7'h4c == total_offset_20[6:0] ? phv_data_76 : _GEN_1306; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1308 = 7'h4d == total_offset_20[6:0] ? phv_data_77 : _GEN_1307; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1309 = 7'h4e == total_offset_20[6:0] ? phv_data_78 : _GEN_1308; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1310 = 7'h4f == total_offset_20[6:0] ? phv_data_79 : _GEN_1309; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1311 = 7'h50 == total_offset_20[6:0] ? phv_data_80 : _GEN_1310; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1312 = 7'h51 == total_offset_20[6:0] ? phv_data_81 : _GEN_1311; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1313 = 7'h52 == total_offset_20[6:0] ? phv_data_82 : _GEN_1312; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1314 = 7'h53 == total_offset_20[6:0] ? phv_data_83 : _GEN_1313; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1315 = 7'h54 == total_offset_20[6:0] ? phv_data_84 : _GEN_1314; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1316 = 7'h55 == total_offset_20[6:0] ? phv_data_85 : _GEN_1315; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1317 = 7'h56 == total_offset_20[6:0] ? phv_data_86 : _GEN_1316; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1318 = 7'h57 == total_offset_20[6:0] ? phv_data_87 : _GEN_1317; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1319 = 7'h58 == total_offset_20[6:0] ? phv_data_88 : _GEN_1318; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1320 = 7'h59 == total_offset_20[6:0] ? phv_data_89 : _GEN_1319; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1321 = 7'h5a == total_offset_20[6:0] ? phv_data_90 : _GEN_1320; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1322 = 7'h5b == total_offset_20[6:0] ? phv_data_91 : _GEN_1321; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1323 = 7'h5c == total_offset_20[6:0] ? phv_data_92 : _GEN_1322; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1324 = 7'h5d == total_offset_20[6:0] ? phv_data_93 : _GEN_1323; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1325 = 7'h5e == total_offset_20[6:0] ? phv_data_94 : _GEN_1324; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1326 = 7'h5f == total_offset_20[6:0] ? phv_data_95 : _GEN_1325; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes_2_4 = 8'h4 < length_1 ? _GEN_1326 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_21 = offset_1 + 8'h5; // @[executor.scala 158:57]
  wire [7:0] _GEN_1329 = 7'h1 == total_offset_21[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1330 = 7'h2 == total_offset_21[6:0] ? phv_data_2 : _GEN_1329; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1331 = 7'h3 == total_offset_21[6:0] ? phv_data_3 : _GEN_1330; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1332 = 7'h4 == total_offset_21[6:0] ? phv_data_4 : _GEN_1331; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1333 = 7'h5 == total_offset_21[6:0] ? phv_data_5 : _GEN_1332; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1334 = 7'h6 == total_offset_21[6:0] ? phv_data_6 : _GEN_1333; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1335 = 7'h7 == total_offset_21[6:0] ? phv_data_7 : _GEN_1334; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1336 = 7'h8 == total_offset_21[6:0] ? phv_data_8 : _GEN_1335; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1337 = 7'h9 == total_offset_21[6:0] ? phv_data_9 : _GEN_1336; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1338 = 7'ha == total_offset_21[6:0] ? phv_data_10 : _GEN_1337; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1339 = 7'hb == total_offset_21[6:0] ? phv_data_11 : _GEN_1338; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1340 = 7'hc == total_offset_21[6:0] ? phv_data_12 : _GEN_1339; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1341 = 7'hd == total_offset_21[6:0] ? phv_data_13 : _GEN_1340; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1342 = 7'he == total_offset_21[6:0] ? phv_data_14 : _GEN_1341; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1343 = 7'hf == total_offset_21[6:0] ? phv_data_15 : _GEN_1342; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1344 = 7'h10 == total_offset_21[6:0] ? phv_data_16 : _GEN_1343; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1345 = 7'h11 == total_offset_21[6:0] ? phv_data_17 : _GEN_1344; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1346 = 7'h12 == total_offset_21[6:0] ? phv_data_18 : _GEN_1345; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1347 = 7'h13 == total_offset_21[6:0] ? phv_data_19 : _GEN_1346; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1348 = 7'h14 == total_offset_21[6:0] ? phv_data_20 : _GEN_1347; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1349 = 7'h15 == total_offset_21[6:0] ? phv_data_21 : _GEN_1348; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1350 = 7'h16 == total_offset_21[6:0] ? phv_data_22 : _GEN_1349; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1351 = 7'h17 == total_offset_21[6:0] ? phv_data_23 : _GEN_1350; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1352 = 7'h18 == total_offset_21[6:0] ? phv_data_24 : _GEN_1351; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1353 = 7'h19 == total_offset_21[6:0] ? phv_data_25 : _GEN_1352; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1354 = 7'h1a == total_offset_21[6:0] ? phv_data_26 : _GEN_1353; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1355 = 7'h1b == total_offset_21[6:0] ? phv_data_27 : _GEN_1354; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1356 = 7'h1c == total_offset_21[6:0] ? phv_data_28 : _GEN_1355; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1357 = 7'h1d == total_offset_21[6:0] ? phv_data_29 : _GEN_1356; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1358 = 7'h1e == total_offset_21[6:0] ? phv_data_30 : _GEN_1357; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1359 = 7'h1f == total_offset_21[6:0] ? phv_data_31 : _GEN_1358; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1360 = 7'h20 == total_offset_21[6:0] ? phv_data_32 : _GEN_1359; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1361 = 7'h21 == total_offset_21[6:0] ? phv_data_33 : _GEN_1360; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1362 = 7'h22 == total_offset_21[6:0] ? phv_data_34 : _GEN_1361; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1363 = 7'h23 == total_offset_21[6:0] ? phv_data_35 : _GEN_1362; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1364 = 7'h24 == total_offset_21[6:0] ? phv_data_36 : _GEN_1363; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1365 = 7'h25 == total_offset_21[6:0] ? phv_data_37 : _GEN_1364; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1366 = 7'h26 == total_offset_21[6:0] ? phv_data_38 : _GEN_1365; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1367 = 7'h27 == total_offset_21[6:0] ? phv_data_39 : _GEN_1366; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1368 = 7'h28 == total_offset_21[6:0] ? phv_data_40 : _GEN_1367; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1369 = 7'h29 == total_offset_21[6:0] ? phv_data_41 : _GEN_1368; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1370 = 7'h2a == total_offset_21[6:0] ? phv_data_42 : _GEN_1369; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1371 = 7'h2b == total_offset_21[6:0] ? phv_data_43 : _GEN_1370; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1372 = 7'h2c == total_offset_21[6:0] ? phv_data_44 : _GEN_1371; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1373 = 7'h2d == total_offset_21[6:0] ? phv_data_45 : _GEN_1372; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1374 = 7'h2e == total_offset_21[6:0] ? phv_data_46 : _GEN_1373; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1375 = 7'h2f == total_offset_21[6:0] ? phv_data_47 : _GEN_1374; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1376 = 7'h30 == total_offset_21[6:0] ? phv_data_48 : _GEN_1375; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1377 = 7'h31 == total_offset_21[6:0] ? phv_data_49 : _GEN_1376; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1378 = 7'h32 == total_offset_21[6:0] ? phv_data_50 : _GEN_1377; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1379 = 7'h33 == total_offset_21[6:0] ? phv_data_51 : _GEN_1378; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1380 = 7'h34 == total_offset_21[6:0] ? phv_data_52 : _GEN_1379; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1381 = 7'h35 == total_offset_21[6:0] ? phv_data_53 : _GEN_1380; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1382 = 7'h36 == total_offset_21[6:0] ? phv_data_54 : _GEN_1381; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1383 = 7'h37 == total_offset_21[6:0] ? phv_data_55 : _GEN_1382; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1384 = 7'h38 == total_offset_21[6:0] ? phv_data_56 : _GEN_1383; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1385 = 7'h39 == total_offset_21[6:0] ? phv_data_57 : _GEN_1384; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1386 = 7'h3a == total_offset_21[6:0] ? phv_data_58 : _GEN_1385; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1387 = 7'h3b == total_offset_21[6:0] ? phv_data_59 : _GEN_1386; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1388 = 7'h3c == total_offset_21[6:0] ? phv_data_60 : _GEN_1387; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1389 = 7'h3d == total_offset_21[6:0] ? phv_data_61 : _GEN_1388; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1390 = 7'h3e == total_offset_21[6:0] ? phv_data_62 : _GEN_1389; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1391 = 7'h3f == total_offset_21[6:0] ? phv_data_63 : _GEN_1390; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1392 = 7'h40 == total_offset_21[6:0] ? phv_data_64 : _GEN_1391; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1393 = 7'h41 == total_offset_21[6:0] ? phv_data_65 : _GEN_1392; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1394 = 7'h42 == total_offset_21[6:0] ? phv_data_66 : _GEN_1393; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1395 = 7'h43 == total_offset_21[6:0] ? phv_data_67 : _GEN_1394; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1396 = 7'h44 == total_offset_21[6:0] ? phv_data_68 : _GEN_1395; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1397 = 7'h45 == total_offset_21[6:0] ? phv_data_69 : _GEN_1396; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1398 = 7'h46 == total_offset_21[6:0] ? phv_data_70 : _GEN_1397; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1399 = 7'h47 == total_offset_21[6:0] ? phv_data_71 : _GEN_1398; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1400 = 7'h48 == total_offset_21[6:0] ? phv_data_72 : _GEN_1399; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1401 = 7'h49 == total_offset_21[6:0] ? phv_data_73 : _GEN_1400; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1402 = 7'h4a == total_offset_21[6:0] ? phv_data_74 : _GEN_1401; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1403 = 7'h4b == total_offset_21[6:0] ? phv_data_75 : _GEN_1402; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1404 = 7'h4c == total_offset_21[6:0] ? phv_data_76 : _GEN_1403; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1405 = 7'h4d == total_offset_21[6:0] ? phv_data_77 : _GEN_1404; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1406 = 7'h4e == total_offset_21[6:0] ? phv_data_78 : _GEN_1405; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1407 = 7'h4f == total_offset_21[6:0] ? phv_data_79 : _GEN_1406; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1408 = 7'h50 == total_offset_21[6:0] ? phv_data_80 : _GEN_1407; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1409 = 7'h51 == total_offset_21[6:0] ? phv_data_81 : _GEN_1408; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1410 = 7'h52 == total_offset_21[6:0] ? phv_data_82 : _GEN_1409; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1411 = 7'h53 == total_offset_21[6:0] ? phv_data_83 : _GEN_1410; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1412 = 7'h54 == total_offset_21[6:0] ? phv_data_84 : _GEN_1411; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1413 = 7'h55 == total_offset_21[6:0] ? phv_data_85 : _GEN_1412; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1414 = 7'h56 == total_offset_21[6:0] ? phv_data_86 : _GEN_1413; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1415 = 7'h57 == total_offset_21[6:0] ? phv_data_87 : _GEN_1414; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1416 = 7'h58 == total_offset_21[6:0] ? phv_data_88 : _GEN_1415; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1417 = 7'h59 == total_offset_21[6:0] ? phv_data_89 : _GEN_1416; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1418 = 7'h5a == total_offset_21[6:0] ? phv_data_90 : _GEN_1417; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1419 = 7'h5b == total_offset_21[6:0] ? phv_data_91 : _GEN_1418; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1420 = 7'h5c == total_offset_21[6:0] ? phv_data_92 : _GEN_1419; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1421 = 7'h5d == total_offset_21[6:0] ? phv_data_93 : _GEN_1420; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1422 = 7'h5e == total_offset_21[6:0] ? phv_data_94 : _GEN_1421; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1423 = 7'h5f == total_offset_21[6:0] ? phv_data_95 : _GEN_1422; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes_2_5 = 8'h5 < length_1 ? _GEN_1423 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_22 = offset_1 + 8'h6; // @[executor.scala 158:57]
  wire [7:0] _GEN_1426 = 7'h1 == total_offset_22[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1427 = 7'h2 == total_offset_22[6:0] ? phv_data_2 : _GEN_1426; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1428 = 7'h3 == total_offset_22[6:0] ? phv_data_3 : _GEN_1427; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1429 = 7'h4 == total_offset_22[6:0] ? phv_data_4 : _GEN_1428; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1430 = 7'h5 == total_offset_22[6:0] ? phv_data_5 : _GEN_1429; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1431 = 7'h6 == total_offset_22[6:0] ? phv_data_6 : _GEN_1430; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1432 = 7'h7 == total_offset_22[6:0] ? phv_data_7 : _GEN_1431; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1433 = 7'h8 == total_offset_22[6:0] ? phv_data_8 : _GEN_1432; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1434 = 7'h9 == total_offset_22[6:0] ? phv_data_9 : _GEN_1433; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1435 = 7'ha == total_offset_22[6:0] ? phv_data_10 : _GEN_1434; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1436 = 7'hb == total_offset_22[6:0] ? phv_data_11 : _GEN_1435; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1437 = 7'hc == total_offset_22[6:0] ? phv_data_12 : _GEN_1436; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1438 = 7'hd == total_offset_22[6:0] ? phv_data_13 : _GEN_1437; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1439 = 7'he == total_offset_22[6:0] ? phv_data_14 : _GEN_1438; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1440 = 7'hf == total_offset_22[6:0] ? phv_data_15 : _GEN_1439; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1441 = 7'h10 == total_offset_22[6:0] ? phv_data_16 : _GEN_1440; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1442 = 7'h11 == total_offset_22[6:0] ? phv_data_17 : _GEN_1441; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1443 = 7'h12 == total_offset_22[6:0] ? phv_data_18 : _GEN_1442; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1444 = 7'h13 == total_offset_22[6:0] ? phv_data_19 : _GEN_1443; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1445 = 7'h14 == total_offset_22[6:0] ? phv_data_20 : _GEN_1444; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1446 = 7'h15 == total_offset_22[6:0] ? phv_data_21 : _GEN_1445; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1447 = 7'h16 == total_offset_22[6:0] ? phv_data_22 : _GEN_1446; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1448 = 7'h17 == total_offset_22[6:0] ? phv_data_23 : _GEN_1447; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1449 = 7'h18 == total_offset_22[6:0] ? phv_data_24 : _GEN_1448; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1450 = 7'h19 == total_offset_22[6:0] ? phv_data_25 : _GEN_1449; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1451 = 7'h1a == total_offset_22[6:0] ? phv_data_26 : _GEN_1450; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1452 = 7'h1b == total_offset_22[6:0] ? phv_data_27 : _GEN_1451; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1453 = 7'h1c == total_offset_22[6:0] ? phv_data_28 : _GEN_1452; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1454 = 7'h1d == total_offset_22[6:0] ? phv_data_29 : _GEN_1453; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1455 = 7'h1e == total_offset_22[6:0] ? phv_data_30 : _GEN_1454; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1456 = 7'h1f == total_offset_22[6:0] ? phv_data_31 : _GEN_1455; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1457 = 7'h20 == total_offset_22[6:0] ? phv_data_32 : _GEN_1456; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1458 = 7'h21 == total_offset_22[6:0] ? phv_data_33 : _GEN_1457; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1459 = 7'h22 == total_offset_22[6:0] ? phv_data_34 : _GEN_1458; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1460 = 7'h23 == total_offset_22[6:0] ? phv_data_35 : _GEN_1459; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1461 = 7'h24 == total_offset_22[6:0] ? phv_data_36 : _GEN_1460; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1462 = 7'h25 == total_offset_22[6:0] ? phv_data_37 : _GEN_1461; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1463 = 7'h26 == total_offset_22[6:0] ? phv_data_38 : _GEN_1462; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1464 = 7'h27 == total_offset_22[6:0] ? phv_data_39 : _GEN_1463; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1465 = 7'h28 == total_offset_22[6:0] ? phv_data_40 : _GEN_1464; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1466 = 7'h29 == total_offset_22[6:0] ? phv_data_41 : _GEN_1465; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1467 = 7'h2a == total_offset_22[6:0] ? phv_data_42 : _GEN_1466; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1468 = 7'h2b == total_offset_22[6:0] ? phv_data_43 : _GEN_1467; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1469 = 7'h2c == total_offset_22[6:0] ? phv_data_44 : _GEN_1468; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1470 = 7'h2d == total_offset_22[6:0] ? phv_data_45 : _GEN_1469; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1471 = 7'h2e == total_offset_22[6:0] ? phv_data_46 : _GEN_1470; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1472 = 7'h2f == total_offset_22[6:0] ? phv_data_47 : _GEN_1471; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1473 = 7'h30 == total_offset_22[6:0] ? phv_data_48 : _GEN_1472; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1474 = 7'h31 == total_offset_22[6:0] ? phv_data_49 : _GEN_1473; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1475 = 7'h32 == total_offset_22[6:0] ? phv_data_50 : _GEN_1474; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1476 = 7'h33 == total_offset_22[6:0] ? phv_data_51 : _GEN_1475; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1477 = 7'h34 == total_offset_22[6:0] ? phv_data_52 : _GEN_1476; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1478 = 7'h35 == total_offset_22[6:0] ? phv_data_53 : _GEN_1477; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1479 = 7'h36 == total_offset_22[6:0] ? phv_data_54 : _GEN_1478; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1480 = 7'h37 == total_offset_22[6:0] ? phv_data_55 : _GEN_1479; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1481 = 7'h38 == total_offset_22[6:0] ? phv_data_56 : _GEN_1480; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1482 = 7'h39 == total_offset_22[6:0] ? phv_data_57 : _GEN_1481; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1483 = 7'h3a == total_offset_22[6:0] ? phv_data_58 : _GEN_1482; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1484 = 7'h3b == total_offset_22[6:0] ? phv_data_59 : _GEN_1483; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1485 = 7'h3c == total_offset_22[6:0] ? phv_data_60 : _GEN_1484; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1486 = 7'h3d == total_offset_22[6:0] ? phv_data_61 : _GEN_1485; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1487 = 7'h3e == total_offset_22[6:0] ? phv_data_62 : _GEN_1486; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1488 = 7'h3f == total_offset_22[6:0] ? phv_data_63 : _GEN_1487; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1489 = 7'h40 == total_offset_22[6:0] ? phv_data_64 : _GEN_1488; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1490 = 7'h41 == total_offset_22[6:0] ? phv_data_65 : _GEN_1489; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1491 = 7'h42 == total_offset_22[6:0] ? phv_data_66 : _GEN_1490; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1492 = 7'h43 == total_offset_22[6:0] ? phv_data_67 : _GEN_1491; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1493 = 7'h44 == total_offset_22[6:0] ? phv_data_68 : _GEN_1492; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1494 = 7'h45 == total_offset_22[6:0] ? phv_data_69 : _GEN_1493; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1495 = 7'h46 == total_offset_22[6:0] ? phv_data_70 : _GEN_1494; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1496 = 7'h47 == total_offset_22[6:0] ? phv_data_71 : _GEN_1495; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1497 = 7'h48 == total_offset_22[6:0] ? phv_data_72 : _GEN_1496; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1498 = 7'h49 == total_offset_22[6:0] ? phv_data_73 : _GEN_1497; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1499 = 7'h4a == total_offset_22[6:0] ? phv_data_74 : _GEN_1498; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1500 = 7'h4b == total_offset_22[6:0] ? phv_data_75 : _GEN_1499; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1501 = 7'h4c == total_offset_22[6:0] ? phv_data_76 : _GEN_1500; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1502 = 7'h4d == total_offset_22[6:0] ? phv_data_77 : _GEN_1501; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1503 = 7'h4e == total_offset_22[6:0] ? phv_data_78 : _GEN_1502; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1504 = 7'h4f == total_offset_22[6:0] ? phv_data_79 : _GEN_1503; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1505 = 7'h50 == total_offset_22[6:0] ? phv_data_80 : _GEN_1504; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1506 = 7'h51 == total_offset_22[6:0] ? phv_data_81 : _GEN_1505; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1507 = 7'h52 == total_offset_22[6:0] ? phv_data_82 : _GEN_1506; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1508 = 7'h53 == total_offset_22[6:0] ? phv_data_83 : _GEN_1507; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1509 = 7'h54 == total_offset_22[6:0] ? phv_data_84 : _GEN_1508; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1510 = 7'h55 == total_offset_22[6:0] ? phv_data_85 : _GEN_1509; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1511 = 7'h56 == total_offset_22[6:0] ? phv_data_86 : _GEN_1510; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1512 = 7'h57 == total_offset_22[6:0] ? phv_data_87 : _GEN_1511; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1513 = 7'h58 == total_offset_22[6:0] ? phv_data_88 : _GEN_1512; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1514 = 7'h59 == total_offset_22[6:0] ? phv_data_89 : _GEN_1513; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1515 = 7'h5a == total_offset_22[6:0] ? phv_data_90 : _GEN_1514; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1516 = 7'h5b == total_offset_22[6:0] ? phv_data_91 : _GEN_1515; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1517 = 7'h5c == total_offset_22[6:0] ? phv_data_92 : _GEN_1516; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1518 = 7'h5d == total_offset_22[6:0] ? phv_data_93 : _GEN_1517; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1519 = 7'h5e == total_offset_22[6:0] ? phv_data_94 : _GEN_1518; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1520 = 7'h5f == total_offset_22[6:0] ? phv_data_95 : _GEN_1519; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes_2_6 = 8'h6 < length_1 ? _GEN_1520 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_23 = offset_1 + 8'h7; // @[executor.scala 158:57]
  wire [7:0] _GEN_1523 = 7'h1 == total_offset_23[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1524 = 7'h2 == total_offset_23[6:0] ? phv_data_2 : _GEN_1523; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1525 = 7'h3 == total_offset_23[6:0] ? phv_data_3 : _GEN_1524; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1526 = 7'h4 == total_offset_23[6:0] ? phv_data_4 : _GEN_1525; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1527 = 7'h5 == total_offset_23[6:0] ? phv_data_5 : _GEN_1526; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1528 = 7'h6 == total_offset_23[6:0] ? phv_data_6 : _GEN_1527; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1529 = 7'h7 == total_offset_23[6:0] ? phv_data_7 : _GEN_1528; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1530 = 7'h8 == total_offset_23[6:0] ? phv_data_8 : _GEN_1529; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1531 = 7'h9 == total_offset_23[6:0] ? phv_data_9 : _GEN_1530; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1532 = 7'ha == total_offset_23[6:0] ? phv_data_10 : _GEN_1531; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1533 = 7'hb == total_offset_23[6:0] ? phv_data_11 : _GEN_1532; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1534 = 7'hc == total_offset_23[6:0] ? phv_data_12 : _GEN_1533; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1535 = 7'hd == total_offset_23[6:0] ? phv_data_13 : _GEN_1534; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1536 = 7'he == total_offset_23[6:0] ? phv_data_14 : _GEN_1535; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1537 = 7'hf == total_offset_23[6:0] ? phv_data_15 : _GEN_1536; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1538 = 7'h10 == total_offset_23[6:0] ? phv_data_16 : _GEN_1537; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1539 = 7'h11 == total_offset_23[6:0] ? phv_data_17 : _GEN_1538; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1540 = 7'h12 == total_offset_23[6:0] ? phv_data_18 : _GEN_1539; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1541 = 7'h13 == total_offset_23[6:0] ? phv_data_19 : _GEN_1540; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1542 = 7'h14 == total_offset_23[6:0] ? phv_data_20 : _GEN_1541; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1543 = 7'h15 == total_offset_23[6:0] ? phv_data_21 : _GEN_1542; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1544 = 7'h16 == total_offset_23[6:0] ? phv_data_22 : _GEN_1543; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1545 = 7'h17 == total_offset_23[6:0] ? phv_data_23 : _GEN_1544; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1546 = 7'h18 == total_offset_23[6:0] ? phv_data_24 : _GEN_1545; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1547 = 7'h19 == total_offset_23[6:0] ? phv_data_25 : _GEN_1546; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1548 = 7'h1a == total_offset_23[6:0] ? phv_data_26 : _GEN_1547; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1549 = 7'h1b == total_offset_23[6:0] ? phv_data_27 : _GEN_1548; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1550 = 7'h1c == total_offset_23[6:0] ? phv_data_28 : _GEN_1549; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1551 = 7'h1d == total_offset_23[6:0] ? phv_data_29 : _GEN_1550; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1552 = 7'h1e == total_offset_23[6:0] ? phv_data_30 : _GEN_1551; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1553 = 7'h1f == total_offset_23[6:0] ? phv_data_31 : _GEN_1552; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1554 = 7'h20 == total_offset_23[6:0] ? phv_data_32 : _GEN_1553; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1555 = 7'h21 == total_offset_23[6:0] ? phv_data_33 : _GEN_1554; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1556 = 7'h22 == total_offset_23[6:0] ? phv_data_34 : _GEN_1555; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1557 = 7'h23 == total_offset_23[6:0] ? phv_data_35 : _GEN_1556; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1558 = 7'h24 == total_offset_23[6:0] ? phv_data_36 : _GEN_1557; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1559 = 7'h25 == total_offset_23[6:0] ? phv_data_37 : _GEN_1558; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1560 = 7'h26 == total_offset_23[6:0] ? phv_data_38 : _GEN_1559; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1561 = 7'h27 == total_offset_23[6:0] ? phv_data_39 : _GEN_1560; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1562 = 7'h28 == total_offset_23[6:0] ? phv_data_40 : _GEN_1561; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1563 = 7'h29 == total_offset_23[6:0] ? phv_data_41 : _GEN_1562; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1564 = 7'h2a == total_offset_23[6:0] ? phv_data_42 : _GEN_1563; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1565 = 7'h2b == total_offset_23[6:0] ? phv_data_43 : _GEN_1564; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1566 = 7'h2c == total_offset_23[6:0] ? phv_data_44 : _GEN_1565; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1567 = 7'h2d == total_offset_23[6:0] ? phv_data_45 : _GEN_1566; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1568 = 7'h2e == total_offset_23[6:0] ? phv_data_46 : _GEN_1567; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1569 = 7'h2f == total_offset_23[6:0] ? phv_data_47 : _GEN_1568; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1570 = 7'h30 == total_offset_23[6:0] ? phv_data_48 : _GEN_1569; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1571 = 7'h31 == total_offset_23[6:0] ? phv_data_49 : _GEN_1570; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1572 = 7'h32 == total_offset_23[6:0] ? phv_data_50 : _GEN_1571; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1573 = 7'h33 == total_offset_23[6:0] ? phv_data_51 : _GEN_1572; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1574 = 7'h34 == total_offset_23[6:0] ? phv_data_52 : _GEN_1573; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1575 = 7'h35 == total_offset_23[6:0] ? phv_data_53 : _GEN_1574; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1576 = 7'h36 == total_offset_23[6:0] ? phv_data_54 : _GEN_1575; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1577 = 7'h37 == total_offset_23[6:0] ? phv_data_55 : _GEN_1576; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1578 = 7'h38 == total_offset_23[6:0] ? phv_data_56 : _GEN_1577; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1579 = 7'h39 == total_offset_23[6:0] ? phv_data_57 : _GEN_1578; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1580 = 7'h3a == total_offset_23[6:0] ? phv_data_58 : _GEN_1579; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1581 = 7'h3b == total_offset_23[6:0] ? phv_data_59 : _GEN_1580; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1582 = 7'h3c == total_offset_23[6:0] ? phv_data_60 : _GEN_1581; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1583 = 7'h3d == total_offset_23[6:0] ? phv_data_61 : _GEN_1582; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1584 = 7'h3e == total_offset_23[6:0] ? phv_data_62 : _GEN_1583; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1585 = 7'h3f == total_offset_23[6:0] ? phv_data_63 : _GEN_1584; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1586 = 7'h40 == total_offset_23[6:0] ? phv_data_64 : _GEN_1585; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1587 = 7'h41 == total_offset_23[6:0] ? phv_data_65 : _GEN_1586; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1588 = 7'h42 == total_offset_23[6:0] ? phv_data_66 : _GEN_1587; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1589 = 7'h43 == total_offset_23[6:0] ? phv_data_67 : _GEN_1588; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1590 = 7'h44 == total_offset_23[6:0] ? phv_data_68 : _GEN_1589; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1591 = 7'h45 == total_offset_23[6:0] ? phv_data_69 : _GEN_1590; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1592 = 7'h46 == total_offset_23[6:0] ? phv_data_70 : _GEN_1591; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1593 = 7'h47 == total_offset_23[6:0] ? phv_data_71 : _GEN_1592; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1594 = 7'h48 == total_offset_23[6:0] ? phv_data_72 : _GEN_1593; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1595 = 7'h49 == total_offset_23[6:0] ? phv_data_73 : _GEN_1594; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1596 = 7'h4a == total_offset_23[6:0] ? phv_data_74 : _GEN_1595; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1597 = 7'h4b == total_offset_23[6:0] ? phv_data_75 : _GEN_1596; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1598 = 7'h4c == total_offset_23[6:0] ? phv_data_76 : _GEN_1597; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1599 = 7'h4d == total_offset_23[6:0] ? phv_data_77 : _GEN_1598; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1600 = 7'h4e == total_offset_23[6:0] ? phv_data_78 : _GEN_1599; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1601 = 7'h4f == total_offset_23[6:0] ? phv_data_79 : _GEN_1600; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1602 = 7'h50 == total_offset_23[6:0] ? phv_data_80 : _GEN_1601; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1603 = 7'h51 == total_offset_23[6:0] ? phv_data_81 : _GEN_1602; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1604 = 7'h52 == total_offset_23[6:0] ? phv_data_82 : _GEN_1603; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1605 = 7'h53 == total_offset_23[6:0] ? phv_data_83 : _GEN_1604; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1606 = 7'h54 == total_offset_23[6:0] ? phv_data_84 : _GEN_1605; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1607 = 7'h55 == total_offset_23[6:0] ? phv_data_85 : _GEN_1606; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1608 = 7'h56 == total_offset_23[6:0] ? phv_data_86 : _GEN_1607; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1609 = 7'h57 == total_offset_23[6:0] ? phv_data_87 : _GEN_1608; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1610 = 7'h58 == total_offset_23[6:0] ? phv_data_88 : _GEN_1609; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1611 = 7'h59 == total_offset_23[6:0] ? phv_data_89 : _GEN_1610; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1612 = 7'h5a == total_offset_23[6:0] ? phv_data_90 : _GEN_1611; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1613 = 7'h5b == total_offset_23[6:0] ? phv_data_91 : _GEN_1612; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1614 = 7'h5c == total_offset_23[6:0] ? phv_data_92 : _GEN_1613; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1615 = 7'h5d == total_offset_23[6:0] ? phv_data_93 : _GEN_1614; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1616 = 7'h5e == total_offset_23[6:0] ? phv_data_94 : _GEN_1615; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1617 = 7'h5f == total_offset_23[6:0] ? phv_data_95 : _GEN_1616; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes_2_7 = 8'h7 < length_1 ? _GEN_1617 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [63:0] _io_field_out_1_T = {bytes_2_0,bytes_2_1,bytes_2_2,bytes_2_3,bytes_2_4,bytes_2_5,bytes_2_6,bytes_2_7}; // @[Cat.scala 30:58]
  wire [2:0] args_offset_1 = io_field_out_1_lo[13:11]; // @[primitive.scala 34:52]
  wire [2:0] args_length_1 = io_field_out_1_lo[10:8]; // @[primitive.scala 35:52]
  wire [8:0] _total_offset_T_24 = {{6'd0}, args_offset_1}; // @[executor.scala 173:60]
  wire [7:0] total_offset_24 = _total_offset_T_24[7:0]; // @[executor.scala 173:60]
  wire [7:0] _GEN_3386 = {{5'd0}, args_length_1}; // @[executor.scala 174:48]
  wire [7:0] _GEN_1620 = 3'h1 == total_offset_24[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1621 = 3'h2 == total_offset_24[2:0] ? args_2 : _GEN_1620; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1622 = 3'h3 == total_offset_24[2:0] ? args_3 : _GEN_1621; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1623 = 3'h4 == total_offset_24[2:0] ? args_4 : _GEN_1622; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1624 = 3'h5 == total_offset_24[2:0] ? args_5 : _GEN_1623; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1625 = 3'h6 == total_offset_24[2:0] ? args_6 : _GEN_1624; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_3_0 = 8'h0 < _GEN_3386 ? _GEN_1625 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [7:0] _GEN_3387 = {{5'd0}, args_offset_1}; // @[executor.scala 173:60]
  wire [7:0] total_offset_25 = _GEN_3387 + 8'h1; // @[executor.scala 173:60]
  wire [7:0] _GEN_1628 = 3'h1 == total_offset_25[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1629 = 3'h2 == total_offset_25[2:0] ? args_2 : _GEN_1628; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1630 = 3'h3 == total_offset_25[2:0] ? args_3 : _GEN_1629; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1631 = 3'h4 == total_offset_25[2:0] ? args_4 : _GEN_1630; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1632 = 3'h5 == total_offset_25[2:0] ? args_5 : _GEN_1631; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1633 = 3'h6 == total_offset_25[2:0] ? args_6 : _GEN_1632; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_3_1 = 8'h1 < _GEN_3386 ? _GEN_1633 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [7:0] total_offset_26 = _GEN_3387 + 8'h2; // @[executor.scala 173:60]
  wire [7:0] _GEN_1636 = 3'h1 == total_offset_26[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1637 = 3'h2 == total_offset_26[2:0] ? args_2 : _GEN_1636; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1638 = 3'h3 == total_offset_26[2:0] ? args_3 : _GEN_1637; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1639 = 3'h4 == total_offset_26[2:0] ? args_4 : _GEN_1638; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1640 = 3'h5 == total_offset_26[2:0] ? args_5 : _GEN_1639; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1641 = 3'h6 == total_offset_26[2:0] ? args_6 : _GEN_1640; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_3_2 = 8'h2 < _GEN_3386 ? _GEN_1641 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [7:0] total_offset_27 = _GEN_3387 + 8'h3; // @[executor.scala 173:60]
  wire [7:0] _GEN_1644 = 3'h1 == total_offset_27[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1645 = 3'h2 == total_offset_27[2:0] ? args_2 : _GEN_1644; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1646 = 3'h3 == total_offset_27[2:0] ? args_3 : _GEN_1645; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1647 = 3'h4 == total_offset_27[2:0] ? args_4 : _GEN_1646; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1648 = 3'h5 == total_offset_27[2:0] ? args_5 : _GEN_1647; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1649 = 3'h6 == total_offset_27[2:0] ? args_6 : _GEN_1648; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_3_3 = 8'h3 < _GEN_3386 ? _GEN_1649 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [7:0] total_offset_28 = _GEN_3387 + 8'h4; // @[executor.scala 173:60]
  wire [7:0] _GEN_1652 = 3'h1 == total_offset_28[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1653 = 3'h2 == total_offset_28[2:0] ? args_2 : _GEN_1652; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1654 = 3'h3 == total_offset_28[2:0] ? args_3 : _GEN_1653; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1655 = 3'h4 == total_offset_28[2:0] ? args_4 : _GEN_1654; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1656 = 3'h5 == total_offset_28[2:0] ? args_5 : _GEN_1655; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1657 = 3'h6 == total_offset_28[2:0] ? args_6 : _GEN_1656; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_3_4 = 8'h4 < _GEN_3386 ? _GEN_1657 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [7:0] total_offset_29 = _GEN_3387 + 8'h5; // @[executor.scala 173:60]
  wire [7:0] _GEN_1660 = 3'h1 == total_offset_29[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1661 = 3'h2 == total_offset_29[2:0] ? args_2 : _GEN_1660; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1662 = 3'h3 == total_offset_29[2:0] ? args_3 : _GEN_1661; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1663 = 3'h4 == total_offset_29[2:0] ? args_4 : _GEN_1662; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1664 = 3'h5 == total_offset_29[2:0] ? args_5 : _GEN_1663; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1665 = 3'h6 == total_offset_29[2:0] ? args_6 : _GEN_1664; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_3_5 = 8'h5 < _GEN_3386 ? _GEN_1665 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [7:0] total_offset_30 = _GEN_3387 + 8'h6; // @[executor.scala 173:60]
  wire [7:0] _GEN_1668 = 3'h1 == total_offset_30[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1669 = 3'h2 == total_offset_30[2:0] ? args_2 : _GEN_1668; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1670 = 3'h3 == total_offset_30[2:0] ? args_3 : _GEN_1669; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1671 = 3'h4 == total_offset_30[2:0] ? args_4 : _GEN_1670; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1672 = 3'h5 == total_offset_30[2:0] ? args_5 : _GEN_1671; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_1673 = 3'h6 == total_offset_30[2:0] ? args_6 : _GEN_1672; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_3_6 = 8'h6 < _GEN_3386 ? _GEN_1673 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [63:0] _io_field_out_1_T_1 = {bytes_3_0,bytes_3_1,bytes_3_2,bytes_3_3,bytes_3_4,bytes_3_5,bytes_3_6,8'h0}; // @[Cat.scala 30:58]
  wire [49:0] io_field_out_1_hi_12 = io_field_out_1_lo[13] ? 50'h3ffffffffffff : 50'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _io_field_out_1_T_4 = {io_field_out_1_hi_12,io_field_out_1_lo}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_1683 = 4'ha == opcode_1 ? _io_field_out_1_T_1 : _io_field_out_1_T_4; // @[executor.scala 167:55 executor.scala 180:41 executor.scala 183:41]
  wire [63:0] _GEN_1684 = from_header_1 ? _io_field_out_1_T : _GEN_1683; // @[executor.scala 152:36 executor.scala 165:37]
  wire [3:0] opcode_2 = vliw_2[31:28]; // @[primitive.scala 9:44]
  wire [13:0] io_field_out_2_lo = vliw_2[13:0]; // @[primitive.scala 11:44]
  wire  from_header_2 = length_2 != 8'h0; // @[executor.scala 151:45]
  wire [8:0] _total_offset_T_32 = {{1'd0}, offset_2}; // @[executor.scala 158:57]
  wire [7:0] total_offset_32 = _total_offset_T_32[7:0]; // @[executor.scala 158:57]
  wire [7:0] _GEN_1687 = 7'h1 == total_offset_32[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1688 = 7'h2 == total_offset_32[6:0] ? phv_data_2 : _GEN_1687; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1689 = 7'h3 == total_offset_32[6:0] ? phv_data_3 : _GEN_1688; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1690 = 7'h4 == total_offset_32[6:0] ? phv_data_4 : _GEN_1689; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1691 = 7'h5 == total_offset_32[6:0] ? phv_data_5 : _GEN_1690; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1692 = 7'h6 == total_offset_32[6:0] ? phv_data_6 : _GEN_1691; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1693 = 7'h7 == total_offset_32[6:0] ? phv_data_7 : _GEN_1692; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1694 = 7'h8 == total_offset_32[6:0] ? phv_data_8 : _GEN_1693; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1695 = 7'h9 == total_offset_32[6:0] ? phv_data_9 : _GEN_1694; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1696 = 7'ha == total_offset_32[6:0] ? phv_data_10 : _GEN_1695; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1697 = 7'hb == total_offset_32[6:0] ? phv_data_11 : _GEN_1696; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1698 = 7'hc == total_offset_32[6:0] ? phv_data_12 : _GEN_1697; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1699 = 7'hd == total_offset_32[6:0] ? phv_data_13 : _GEN_1698; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1700 = 7'he == total_offset_32[6:0] ? phv_data_14 : _GEN_1699; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1701 = 7'hf == total_offset_32[6:0] ? phv_data_15 : _GEN_1700; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1702 = 7'h10 == total_offset_32[6:0] ? phv_data_16 : _GEN_1701; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1703 = 7'h11 == total_offset_32[6:0] ? phv_data_17 : _GEN_1702; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1704 = 7'h12 == total_offset_32[6:0] ? phv_data_18 : _GEN_1703; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1705 = 7'h13 == total_offset_32[6:0] ? phv_data_19 : _GEN_1704; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1706 = 7'h14 == total_offset_32[6:0] ? phv_data_20 : _GEN_1705; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1707 = 7'h15 == total_offset_32[6:0] ? phv_data_21 : _GEN_1706; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1708 = 7'h16 == total_offset_32[6:0] ? phv_data_22 : _GEN_1707; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1709 = 7'h17 == total_offset_32[6:0] ? phv_data_23 : _GEN_1708; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1710 = 7'h18 == total_offset_32[6:0] ? phv_data_24 : _GEN_1709; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1711 = 7'h19 == total_offset_32[6:0] ? phv_data_25 : _GEN_1710; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1712 = 7'h1a == total_offset_32[6:0] ? phv_data_26 : _GEN_1711; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1713 = 7'h1b == total_offset_32[6:0] ? phv_data_27 : _GEN_1712; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1714 = 7'h1c == total_offset_32[6:0] ? phv_data_28 : _GEN_1713; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1715 = 7'h1d == total_offset_32[6:0] ? phv_data_29 : _GEN_1714; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1716 = 7'h1e == total_offset_32[6:0] ? phv_data_30 : _GEN_1715; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1717 = 7'h1f == total_offset_32[6:0] ? phv_data_31 : _GEN_1716; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1718 = 7'h20 == total_offset_32[6:0] ? phv_data_32 : _GEN_1717; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1719 = 7'h21 == total_offset_32[6:0] ? phv_data_33 : _GEN_1718; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1720 = 7'h22 == total_offset_32[6:0] ? phv_data_34 : _GEN_1719; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1721 = 7'h23 == total_offset_32[6:0] ? phv_data_35 : _GEN_1720; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1722 = 7'h24 == total_offset_32[6:0] ? phv_data_36 : _GEN_1721; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1723 = 7'h25 == total_offset_32[6:0] ? phv_data_37 : _GEN_1722; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1724 = 7'h26 == total_offset_32[6:0] ? phv_data_38 : _GEN_1723; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1725 = 7'h27 == total_offset_32[6:0] ? phv_data_39 : _GEN_1724; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1726 = 7'h28 == total_offset_32[6:0] ? phv_data_40 : _GEN_1725; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1727 = 7'h29 == total_offset_32[6:0] ? phv_data_41 : _GEN_1726; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1728 = 7'h2a == total_offset_32[6:0] ? phv_data_42 : _GEN_1727; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1729 = 7'h2b == total_offset_32[6:0] ? phv_data_43 : _GEN_1728; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1730 = 7'h2c == total_offset_32[6:0] ? phv_data_44 : _GEN_1729; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1731 = 7'h2d == total_offset_32[6:0] ? phv_data_45 : _GEN_1730; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1732 = 7'h2e == total_offset_32[6:0] ? phv_data_46 : _GEN_1731; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1733 = 7'h2f == total_offset_32[6:0] ? phv_data_47 : _GEN_1732; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1734 = 7'h30 == total_offset_32[6:0] ? phv_data_48 : _GEN_1733; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1735 = 7'h31 == total_offset_32[6:0] ? phv_data_49 : _GEN_1734; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1736 = 7'h32 == total_offset_32[6:0] ? phv_data_50 : _GEN_1735; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1737 = 7'h33 == total_offset_32[6:0] ? phv_data_51 : _GEN_1736; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1738 = 7'h34 == total_offset_32[6:0] ? phv_data_52 : _GEN_1737; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1739 = 7'h35 == total_offset_32[6:0] ? phv_data_53 : _GEN_1738; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1740 = 7'h36 == total_offset_32[6:0] ? phv_data_54 : _GEN_1739; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1741 = 7'h37 == total_offset_32[6:0] ? phv_data_55 : _GEN_1740; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1742 = 7'h38 == total_offset_32[6:0] ? phv_data_56 : _GEN_1741; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1743 = 7'h39 == total_offset_32[6:0] ? phv_data_57 : _GEN_1742; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1744 = 7'h3a == total_offset_32[6:0] ? phv_data_58 : _GEN_1743; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1745 = 7'h3b == total_offset_32[6:0] ? phv_data_59 : _GEN_1744; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1746 = 7'h3c == total_offset_32[6:0] ? phv_data_60 : _GEN_1745; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1747 = 7'h3d == total_offset_32[6:0] ? phv_data_61 : _GEN_1746; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1748 = 7'h3e == total_offset_32[6:0] ? phv_data_62 : _GEN_1747; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1749 = 7'h3f == total_offset_32[6:0] ? phv_data_63 : _GEN_1748; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1750 = 7'h40 == total_offset_32[6:0] ? phv_data_64 : _GEN_1749; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1751 = 7'h41 == total_offset_32[6:0] ? phv_data_65 : _GEN_1750; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1752 = 7'h42 == total_offset_32[6:0] ? phv_data_66 : _GEN_1751; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1753 = 7'h43 == total_offset_32[6:0] ? phv_data_67 : _GEN_1752; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1754 = 7'h44 == total_offset_32[6:0] ? phv_data_68 : _GEN_1753; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1755 = 7'h45 == total_offset_32[6:0] ? phv_data_69 : _GEN_1754; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1756 = 7'h46 == total_offset_32[6:0] ? phv_data_70 : _GEN_1755; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1757 = 7'h47 == total_offset_32[6:0] ? phv_data_71 : _GEN_1756; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1758 = 7'h48 == total_offset_32[6:0] ? phv_data_72 : _GEN_1757; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1759 = 7'h49 == total_offset_32[6:0] ? phv_data_73 : _GEN_1758; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1760 = 7'h4a == total_offset_32[6:0] ? phv_data_74 : _GEN_1759; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1761 = 7'h4b == total_offset_32[6:0] ? phv_data_75 : _GEN_1760; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1762 = 7'h4c == total_offset_32[6:0] ? phv_data_76 : _GEN_1761; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1763 = 7'h4d == total_offset_32[6:0] ? phv_data_77 : _GEN_1762; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1764 = 7'h4e == total_offset_32[6:0] ? phv_data_78 : _GEN_1763; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1765 = 7'h4f == total_offset_32[6:0] ? phv_data_79 : _GEN_1764; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1766 = 7'h50 == total_offset_32[6:0] ? phv_data_80 : _GEN_1765; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1767 = 7'h51 == total_offset_32[6:0] ? phv_data_81 : _GEN_1766; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1768 = 7'h52 == total_offset_32[6:0] ? phv_data_82 : _GEN_1767; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1769 = 7'h53 == total_offset_32[6:0] ? phv_data_83 : _GEN_1768; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1770 = 7'h54 == total_offset_32[6:0] ? phv_data_84 : _GEN_1769; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1771 = 7'h55 == total_offset_32[6:0] ? phv_data_85 : _GEN_1770; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1772 = 7'h56 == total_offset_32[6:0] ? phv_data_86 : _GEN_1771; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1773 = 7'h57 == total_offset_32[6:0] ? phv_data_87 : _GEN_1772; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1774 = 7'h58 == total_offset_32[6:0] ? phv_data_88 : _GEN_1773; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1775 = 7'h59 == total_offset_32[6:0] ? phv_data_89 : _GEN_1774; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1776 = 7'h5a == total_offset_32[6:0] ? phv_data_90 : _GEN_1775; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1777 = 7'h5b == total_offset_32[6:0] ? phv_data_91 : _GEN_1776; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1778 = 7'h5c == total_offset_32[6:0] ? phv_data_92 : _GEN_1777; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1779 = 7'h5d == total_offset_32[6:0] ? phv_data_93 : _GEN_1778; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1780 = 7'h5e == total_offset_32[6:0] ? phv_data_94 : _GEN_1779; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1781 = 7'h5f == total_offset_32[6:0] ? phv_data_95 : _GEN_1780; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes_4_0 = 8'h0 < length_2 ? _GEN_1781 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_33 = offset_2 + 8'h1; // @[executor.scala 158:57]
  wire [7:0] _GEN_1784 = 7'h1 == total_offset_33[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1785 = 7'h2 == total_offset_33[6:0] ? phv_data_2 : _GEN_1784; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1786 = 7'h3 == total_offset_33[6:0] ? phv_data_3 : _GEN_1785; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1787 = 7'h4 == total_offset_33[6:0] ? phv_data_4 : _GEN_1786; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1788 = 7'h5 == total_offset_33[6:0] ? phv_data_5 : _GEN_1787; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1789 = 7'h6 == total_offset_33[6:0] ? phv_data_6 : _GEN_1788; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1790 = 7'h7 == total_offset_33[6:0] ? phv_data_7 : _GEN_1789; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1791 = 7'h8 == total_offset_33[6:0] ? phv_data_8 : _GEN_1790; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1792 = 7'h9 == total_offset_33[6:0] ? phv_data_9 : _GEN_1791; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1793 = 7'ha == total_offset_33[6:0] ? phv_data_10 : _GEN_1792; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1794 = 7'hb == total_offset_33[6:0] ? phv_data_11 : _GEN_1793; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1795 = 7'hc == total_offset_33[6:0] ? phv_data_12 : _GEN_1794; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1796 = 7'hd == total_offset_33[6:0] ? phv_data_13 : _GEN_1795; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1797 = 7'he == total_offset_33[6:0] ? phv_data_14 : _GEN_1796; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1798 = 7'hf == total_offset_33[6:0] ? phv_data_15 : _GEN_1797; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1799 = 7'h10 == total_offset_33[6:0] ? phv_data_16 : _GEN_1798; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1800 = 7'h11 == total_offset_33[6:0] ? phv_data_17 : _GEN_1799; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1801 = 7'h12 == total_offset_33[6:0] ? phv_data_18 : _GEN_1800; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1802 = 7'h13 == total_offset_33[6:0] ? phv_data_19 : _GEN_1801; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1803 = 7'h14 == total_offset_33[6:0] ? phv_data_20 : _GEN_1802; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1804 = 7'h15 == total_offset_33[6:0] ? phv_data_21 : _GEN_1803; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1805 = 7'h16 == total_offset_33[6:0] ? phv_data_22 : _GEN_1804; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1806 = 7'h17 == total_offset_33[6:0] ? phv_data_23 : _GEN_1805; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1807 = 7'h18 == total_offset_33[6:0] ? phv_data_24 : _GEN_1806; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1808 = 7'h19 == total_offset_33[6:0] ? phv_data_25 : _GEN_1807; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1809 = 7'h1a == total_offset_33[6:0] ? phv_data_26 : _GEN_1808; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1810 = 7'h1b == total_offset_33[6:0] ? phv_data_27 : _GEN_1809; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1811 = 7'h1c == total_offset_33[6:0] ? phv_data_28 : _GEN_1810; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1812 = 7'h1d == total_offset_33[6:0] ? phv_data_29 : _GEN_1811; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1813 = 7'h1e == total_offset_33[6:0] ? phv_data_30 : _GEN_1812; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1814 = 7'h1f == total_offset_33[6:0] ? phv_data_31 : _GEN_1813; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1815 = 7'h20 == total_offset_33[6:0] ? phv_data_32 : _GEN_1814; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1816 = 7'h21 == total_offset_33[6:0] ? phv_data_33 : _GEN_1815; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1817 = 7'h22 == total_offset_33[6:0] ? phv_data_34 : _GEN_1816; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1818 = 7'h23 == total_offset_33[6:0] ? phv_data_35 : _GEN_1817; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1819 = 7'h24 == total_offset_33[6:0] ? phv_data_36 : _GEN_1818; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1820 = 7'h25 == total_offset_33[6:0] ? phv_data_37 : _GEN_1819; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1821 = 7'h26 == total_offset_33[6:0] ? phv_data_38 : _GEN_1820; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1822 = 7'h27 == total_offset_33[6:0] ? phv_data_39 : _GEN_1821; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1823 = 7'h28 == total_offset_33[6:0] ? phv_data_40 : _GEN_1822; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1824 = 7'h29 == total_offset_33[6:0] ? phv_data_41 : _GEN_1823; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1825 = 7'h2a == total_offset_33[6:0] ? phv_data_42 : _GEN_1824; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1826 = 7'h2b == total_offset_33[6:0] ? phv_data_43 : _GEN_1825; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1827 = 7'h2c == total_offset_33[6:0] ? phv_data_44 : _GEN_1826; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1828 = 7'h2d == total_offset_33[6:0] ? phv_data_45 : _GEN_1827; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1829 = 7'h2e == total_offset_33[6:0] ? phv_data_46 : _GEN_1828; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1830 = 7'h2f == total_offset_33[6:0] ? phv_data_47 : _GEN_1829; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1831 = 7'h30 == total_offset_33[6:0] ? phv_data_48 : _GEN_1830; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1832 = 7'h31 == total_offset_33[6:0] ? phv_data_49 : _GEN_1831; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1833 = 7'h32 == total_offset_33[6:0] ? phv_data_50 : _GEN_1832; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1834 = 7'h33 == total_offset_33[6:0] ? phv_data_51 : _GEN_1833; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1835 = 7'h34 == total_offset_33[6:0] ? phv_data_52 : _GEN_1834; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1836 = 7'h35 == total_offset_33[6:0] ? phv_data_53 : _GEN_1835; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1837 = 7'h36 == total_offset_33[6:0] ? phv_data_54 : _GEN_1836; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1838 = 7'h37 == total_offset_33[6:0] ? phv_data_55 : _GEN_1837; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1839 = 7'h38 == total_offset_33[6:0] ? phv_data_56 : _GEN_1838; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1840 = 7'h39 == total_offset_33[6:0] ? phv_data_57 : _GEN_1839; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1841 = 7'h3a == total_offset_33[6:0] ? phv_data_58 : _GEN_1840; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1842 = 7'h3b == total_offset_33[6:0] ? phv_data_59 : _GEN_1841; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1843 = 7'h3c == total_offset_33[6:0] ? phv_data_60 : _GEN_1842; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1844 = 7'h3d == total_offset_33[6:0] ? phv_data_61 : _GEN_1843; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1845 = 7'h3e == total_offset_33[6:0] ? phv_data_62 : _GEN_1844; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1846 = 7'h3f == total_offset_33[6:0] ? phv_data_63 : _GEN_1845; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1847 = 7'h40 == total_offset_33[6:0] ? phv_data_64 : _GEN_1846; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1848 = 7'h41 == total_offset_33[6:0] ? phv_data_65 : _GEN_1847; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1849 = 7'h42 == total_offset_33[6:0] ? phv_data_66 : _GEN_1848; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1850 = 7'h43 == total_offset_33[6:0] ? phv_data_67 : _GEN_1849; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1851 = 7'h44 == total_offset_33[6:0] ? phv_data_68 : _GEN_1850; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1852 = 7'h45 == total_offset_33[6:0] ? phv_data_69 : _GEN_1851; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1853 = 7'h46 == total_offset_33[6:0] ? phv_data_70 : _GEN_1852; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1854 = 7'h47 == total_offset_33[6:0] ? phv_data_71 : _GEN_1853; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1855 = 7'h48 == total_offset_33[6:0] ? phv_data_72 : _GEN_1854; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1856 = 7'h49 == total_offset_33[6:0] ? phv_data_73 : _GEN_1855; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1857 = 7'h4a == total_offset_33[6:0] ? phv_data_74 : _GEN_1856; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1858 = 7'h4b == total_offset_33[6:0] ? phv_data_75 : _GEN_1857; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1859 = 7'h4c == total_offset_33[6:0] ? phv_data_76 : _GEN_1858; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1860 = 7'h4d == total_offset_33[6:0] ? phv_data_77 : _GEN_1859; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1861 = 7'h4e == total_offset_33[6:0] ? phv_data_78 : _GEN_1860; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1862 = 7'h4f == total_offset_33[6:0] ? phv_data_79 : _GEN_1861; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1863 = 7'h50 == total_offset_33[6:0] ? phv_data_80 : _GEN_1862; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1864 = 7'h51 == total_offset_33[6:0] ? phv_data_81 : _GEN_1863; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1865 = 7'h52 == total_offset_33[6:0] ? phv_data_82 : _GEN_1864; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1866 = 7'h53 == total_offset_33[6:0] ? phv_data_83 : _GEN_1865; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1867 = 7'h54 == total_offset_33[6:0] ? phv_data_84 : _GEN_1866; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1868 = 7'h55 == total_offset_33[6:0] ? phv_data_85 : _GEN_1867; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1869 = 7'h56 == total_offset_33[6:0] ? phv_data_86 : _GEN_1868; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1870 = 7'h57 == total_offset_33[6:0] ? phv_data_87 : _GEN_1869; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1871 = 7'h58 == total_offset_33[6:0] ? phv_data_88 : _GEN_1870; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1872 = 7'h59 == total_offset_33[6:0] ? phv_data_89 : _GEN_1871; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1873 = 7'h5a == total_offset_33[6:0] ? phv_data_90 : _GEN_1872; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1874 = 7'h5b == total_offset_33[6:0] ? phv_data_91 : _GEN_1873; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1875 = 7'h5c == total_offset_33[6:0] ? phv_data_92 : _GEN_1874; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1876 = 7'h5d == total_offset_33[6:0] ? phv_data_93 : _GEN_1875; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1877 = 7'h5e == total_offset_33[6:0] ? phv_data_94 : _GEN_1876; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1878 = 7'h5f == total_offset_33[6:0] ? phv_data_95 : _GEN_1877; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes_4_1 = 8'h1 < length_2 ? _GEN_1878 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_34 = offset_2 + 8'h2; // @[executor.scala 158:57]
  wire [7:0] _GEN_1881 = 7'h1 == total_offset_34[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1882 = 7'h2 == total_offset_34[6:0] ? phv_data_2 : _GEN_1881; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1883 = 7'h3 == total_offset_34[6:0] ? phv_data_3 : _GEN_1882; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1884 = 7'h4 == total_offset_34[6:0] ? phv_data_4 : _GEN_1883; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1885 = 7'h5 == total_offset_34[6:0] ? phv_data_5 : _GEN_1884; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1886 = 7'h6 == total_offset_34[6:0] ? phv_data_6 : _GEN_1885; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1887 = 7'h7 == total_offset_34[6:0] ? phv_data_7 : _GEN_1886; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1888 = 7'h8 == total_offset_34[6:0] ? phv_data_8 : _GEN_1887; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1889 = 7'h9 == total_offset_34[6:0] ? phv_data_9 : _GEN_1888; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1890 = 7'ha == total_offset_34[6:0] ? phv_data_10 : _GEN_1889; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1891 = 7'hb == total_offset_34[6:0] ? phv_data_11 : _GEN_1890; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1892 = 7'hc == total_offset_34[6:0] ? phv_data_12 : _GEN_1891; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1893 = 7'hd == total_offset_34[6:0] ? phv_data_13 : _GEN_1892; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1894 = 7'he == total_offset_34[6:0] ? phv_data_14 : _GEN_1893; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1895 = 7'hf == total_offset_34[6:0] ? phv_data_15 : _GEN_1894; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1896 = 7'h10 == total_offset_34[6:0] ? phv_data_16 : _GEN_1895; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1897 = 7'h11 == total_offset_34[6:0] ? phv_data_17 : _GEN_1896; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1898 = 7'h12 == total_offset_34[6:0] ? phv_data_18 : _GEN_1897; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1899 = 7'h13 == total_offset_34[6:0] ? phv_data_19 : _GEN_1898; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1900 = 7'h14 == total_offset_34[6:0] ? phv_data_20 : _GEN_1899; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1901 = 7'h15 == total_offset_34[6:0] ? phv_data_21 : _GEN_1900; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1902 = 7'h16 == total_offset_34[6:0] ? phv_data_22 : _GEN_1901; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1903 = 7'h17 == total_offset_34[6:0] ? phv_data_23 : _GEN_1902; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1904 = 7'h18 == total_offset_34[6:0] ? phv_data_24 : _GEN_1903; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1905 = 7'h19 == total_offset_34[6:0] ? phv_data_25 : _GEN_1904; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1906 = 7'h1a == total_offset_34[6:0] ? phv_data_26 : _GEN_1905; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1907 = 7'h1b == total_offset_34[6:0] ? phv_data_27 : _GEN_1906; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1908 = 7'h1c == total_offset_34[6:0] ? phv_data_28 : _GEN_1907; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1909 = 7'h1d == total_offset_34[6:0] ? phv_data_29 : _GEN_1908; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1910 = 7'h1e == total_offset_34[6:0] ? phv_data_30 : _GEN_1909; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1911 = 7'h1f == total_offset_34[6:0] ? phv_data_31 : _GEN_1910; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1912 = 7'h20 == total_offset_34[6:0] ? phv_data_32 : _GEN_1911; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1913 = 7'h21 == total_offset_34[6:0] ? phv_data_33 : _GEN_1912; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1914 = 7'h22 == total_offset_34[6:0] ? phv_data_34 : _GEN_1913; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1915 = 7'h23 == total_offset_34[6:0] ? phv_data_35 : _GEN_1914; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1916 = 7'h24 == total_offset_34[6:0] ? phv_data_36 : _GEN_1915; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1917 = 7'h25 == total_offset_34[6:0] ? phv_data_37 : _GEN_1916; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1918 = 7'h26 == total_offset_34[6:0] ? phv_data_38 : _GEN_1917; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1919 = 7'h27 == total_offset_34[6:0] ? phv_data_39 : _GEN_1918; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1920 = 7'h28 == total_offset_34[6:0] ? phv_data_40 : _GEN_1919; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1921 = 7'h29 == total_offset_34[6:0] ? phv_data_41 : _GEN_1920; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1922 = 7'h2a == total_offset_34[6:0] ? phv_data_42 : _GEN_1921; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1923 = 7'h2b == total_offset_34[6:0] ? phv_data_43 : _GEN_1922; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1924 = 7'h2c == total_offset_34[6:0] ? phv_data_44 : _GEN_1923; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1925 = 7'h2d == total_offset_34[6:0] ? phv_data_45 : _GEN_1924; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1926 = 7'h2e == total_offset_34[6:0] ? phv_data_46 : _GEN_1925; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1927 = 7'h2f == total_offset_34[6:0] ? phv_data_47 : _GEN_1926; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1928 = 7'h30 == total_offset_34[6:0] ? phv_data_48 : _GEN_1927; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1929 = 7'h31 == total_offset_34[6:0] ? phv_data_49 : _GEN_1928; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1930 = 7'h32 == total_offset_34[6:0] ? phv_data_50 : _GEN_1929; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1931 = 7'h33 == total_offset_34[6:0] ? phv_data_51 : _GEN_1930; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1932 = 7'h34 == total_offset_34[6:0] ? phv_data_52 : _GEN_1931; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1933 = 7'h35 == total_offset_34[6:0] ? phv_data_53 : _GEN_1932; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1934 = 7'h36 == total_offset_34[6:0] ? phv_data_54 : _GEN_1933; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1935 = 7'h37 == total_offset_34[6:0] ? phv_data_55 : _GEN_1934; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1936 = 7'h38 == total_offset_34[6:0] ? phv_data_56 : _GEN_1935; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1937 = 7'h39 == total_offset_34[6:0] ? phv_data_57 : _GEN_1936; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1938 = 7'h3a == total_offset_34[6:0] ? phv_data_58 : _GEN_1937; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1939 = 7'h3b == total_offset_34[6:0] ? phv_data_59 : _GEN_1938; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1940 = 7'h3c == total_offset_34[6:0] ? phv_data_60 : _GEN_1939; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1941 = 7'h3d == total_offset_34[6:0] ? phv_data_61 : _GEN_1940; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1942 = 7'h3e == total_offset_34[6:0] ? phv_data_62 : _GEN_1941; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1943 = 7'h3f == total_offset_34[6:0] ? phv_data_63 : _GEN_1942; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1944 = 7'h40 == total_offset_34[6:0] ? phv_data_64 : _GEN_1943; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1945 = 7'h41 == total_offset_34[6:0] ? phv_data_65 : _GEN_1944; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1946 = 7'h42 == total_offset_34[6:0] ? phv_data_66 : _GEN_1945; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1947 = 7'h43 == total_offset_34[6:0] ? phv_data_67 : _GEN_1946; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1948 = 7'h44 == total_offset_34[6:0] ? phv_data_68 : _GEN_1947; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1949 = 7'h45 == total_offset_34[6:0] ? phv_data_69 : _GEN_1948; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1950 = 7'h46 == total_offset_34[6:0] ? phv_data_70 : _GEN_1949; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1951 = 7'h47 == total_offset_34[6:0] ? phv_data_71 : _GEN_1950; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1952 = 7'h48 == total_offset_34[6:0] ? phv_data_72 : _GEN_1951; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1953 = 7'h49 == total_offset_34[6:0] ? phv_data_73 : _GEN_1952; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1954 = 7'h4a == total_offset_34[6:0] ? phv_data_74 : _GEN_1953; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1955 = 7'h4b == total_offset_34[6:0] ? phv_data_75 : _GEN_1954; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1956 = 7'h4c == total_offset_34[6:0] ? phv_data_76 : _GEN_1955; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1957 = 7'h4d == total_offset_34[6:0] ? phv_data_77 : _GEN_1956; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1958 = 7'h4e == total_offset_34[6:0] ? phv_data_78 : _GEN_1957; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1959 = 7'h4f == total_offset_34[6:0] ? phv_data_79 : _GEN_1958; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1960 = 7'h50 == total_offset_34[6:0] ? phv_data_80 : _GEN_1959; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1961 = 7'h51 == total_offset_34[6:0] ? phv_data_81 : _GEN_1960; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1962 = 7'h52 == total_offset_34[6:0] ? phv_data_82 : _GEN_1961; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1963 = 7'h53 == total_offset_34[6:0] ? phv_data_83 : _GEN_1962; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1964 = 7'h54 == total_offset_34[6:0] ? phv_data_84 : _GEN_1963; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1965 = 7'h55 == total_offset_34[6:0] ? phv_data_85 : _GEN_1964; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1966 = 7'h56 == total_offset_34[6:0] ? phv_data_86 : _GEN_1965; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1967 = 7'h57 == total_offset_34[6:0] ? phv_data_87 : _GEN_1966; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1968 = 7'h58 == total_offset_34[6:0] ? phv_data_88 : _GEN_1967; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1969 = 7'h59 == total_offset_34[6:0] ? phv_data_89 : _GEN_1968; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1970 = 7'h5a == total_offset_34[6:0] ? phv_data_90 : _GEN_1969; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1971 = 7'h5b == total_offset_34[6:0] ? phv_data_91 : _GEN_1970; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1972 = 7'h5c == total_offset_34[6:0] ? phv_data_92 : _GEN_1971; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1973 = 7'h5d == total_offset_34[6:0] ? phv_data_93 : _GEN_1972; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1974 = 7'h5e == total_offset_34[6:0] ? phv_data_94 : _GEN_1973; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1975 = 7'h5f == total_offset_34[6:0] ? phv_data_95 : _GEN_1974; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes_4_2 = 8'h2 < length_2 ? _GEN_1975 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_35 = offset_2 + 8'h3; // @[executor.scala 158:57]
  wire [7:0] _GEN_1978 = 7'h1 == total_offset_35[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1979 = 7'h2 == total_offset_35[6:0] ? phv_data_2 : _GEN_1978; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1980 = 7'h3 == total_offset_35[6:0] ? phv_data_3 : _GEN_1979; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1981 = 7'h4 == total_offset_35[6:0] ? phv_data_4 : _GEN_1980; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1982 = 7'h5 == total_offset_35[6:0] ? phv_data_5 : _GEN_1981; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1983 = 7'h6 == total_offset_35[6:0] ? phv_data_6 : _GEN_1982; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1984 = 7'h7 == total_offset_35[6:0] ? phv_data_7 : _GEN_1983; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1985 = 7'h8 == total_offset_35[6:0] ? phv_data_8 : _GEN_1984; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1986 = 7'h9 == total_offset_35[6:0] ? phv_data_9 : _GEN_1985; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1987 = 7'ha == total_offset_35[6:0] ? phv_data_10 : _GEN_1986; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1988 = 7'hb == total_offset_35[6:0] ? phv_data_11 : _GEN_1987; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1989 = 7'hc == total_offset_35[6:0] ? phv_data_12 : _GEN_1988; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1990 = 7'hd == total_offset_35[6:0] ? phv_data_13 : _GEN_1989; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1991 = 7'he == total_offset_35[6:0] ? phv_data_14 : _GEN_1990; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1992 = 7'hf == total_offset_35[6:0] ? phv_data_15 : _GEN_1991; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1993 = 7'h10 == total_offset_35[6:0] ? phv_data_16 : _GEN_1992; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1994 = 7'h11 == total_offset_35[6:0] ? phv_data_17 : _GEN_1993; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1995 = 7'h12 == total_offset_35[6:0] ? phv_data_18 : _GEN_1994; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1996 = 7'h13 == total_offset_35[6:0] ? phv_data_19 : _GEN_1995; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1997 = 7'h14 == total_offset_35[6:0] ? phv_data_20 : _GEN_1996; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1998 = 7'h15 == total_offset_35[6:0] ? phv_data_21 : _GEN_1997; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_1999 = 7'h16 == total_offset_35[6:0] ? phv_data_22 : _GEN_1998; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2000 = 7'h17 == total_offset_35[6:0] ? phv_data_23 : _GEN_1999; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2001 = 7'h18 == total_offset_35[6:0] ? phv_data_24 : _GEN_2000; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2002 = 7'h19 == total_offset_35[6:0] ? phv_data_25 : _GEN_2001; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2003 = 7'h1a == total_offset_35[6:0] ? phv_data_26 : _GEN_2002; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2004 = 7'h1b == total_offset_35[6:0] ? phv_data_27 : _GEN_2003; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2005 = 7'h1c == total_offset_35[6:0] ? phv_data_28 : _GEN_2004; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2006 = 7'h1d == total_offset_35[6:0] ? phv_data_29 : _GEN_2005; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2007 = 7'h1e == total_offset_35[6:0] ? phv_data_30 : _GEN_2006; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2008 = 7'h1f == total_offset_35[6:0] ? phv_data_31 : _GEN_2007; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2009 = 7'h20 == total_offset_35[6:0] ? phv_data_32 : _GEN_2008; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2010 = 7'h21 == total_offset_35[6:0] ? phv_data_33 : _GEN_2009; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2011 = 7'h22 == total_offset_35[6:0] ? phv_data_34 : _GEN_2010; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2012 = 7'h23 == total_offset_35[6:0] ? phv_data_35 : _GEN_2011; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2013 = 7'h24 == total_offset_35[6:0] ? phv_data_36 : _GEN_2012; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2014 = 7'h25 == total_offset_35[6:0] ? phv_data_37 : _GEN_2013; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2015 = 7'h26 == total_offset_35[6:0] ? phv_data_38 : _GEN_2014; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2016 = 7'h27 == total_offset_35[6:0] ? phv_data_39 : _GEN_2015; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2017 = 7'h28 == total_offset_35[6:0] ? phv_data_40 : _GEN_2016; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2018 = 7'h29 == total_offset_35[6:0] ? phv_data_41 : _GEN_2017; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2019 = 7'h2a == total_offset_35[6:0] ? phv_data_42 : _GEN_2018; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2020 = 7'h2b == total_offset_35[6:0] ? phv_data_43 : _GEN_2019; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2021 = 7'h2c == total_offset_35[6:0] ? phv_data_44 : _GEN_2020; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2022 = 7'h2d == total_offset_35[6:0] ? phv_data_45 : _GEN_2021; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2023 = 7'h2e == total_offset_35[6:0] ? phv_data_46 : _GEN_2022; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2024 = 7'h2f == total_offset_35[6:0] ? phv_data_47 : _GEN_2023; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2025 = 7'h30 == total_offset_35[6:0] ? phv_data_48 : _GEN_2024; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2026 = 7'h31 == total_offset_35[6:0] ? phv_data_49 : _GEN_2025; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2027 = 7'h32 == total_offset_35[6:0] ? phv_data_50 : _GEN_2026; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2028 = 7'h33 == total_offset_35[6:0] ? phv_data_51 : _GEN_2027; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2029 = 7'h34 == total_offset_35[6:0] ? phv_data_52 : _GEN_2028; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2030 = 7'h35 == total_offset_35[6:0] ? phv_data_53 : _GEN_2029; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2031 = 7'h36 == total_offset_35[6:0] ? phv_data_54 : _GEN_2030; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2032 = 7'h37 == total_offset_35[6:0] ? phv_data_55 : _GEN_2031; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2033 = 7'h38 == total_offset_35[6:0] ? phv_data_56 : _GEN_2032; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2034 = 7'h39 == total_offset_35[6:0] ? phv_data_57 : _GEN_2033; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2035 = 7'h3a == total_offset_35[6:0] ? phv_data_58 : _GEN_2034; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2036 = 7'h3b == total_offset_35[6:0] ? phv_data_59 : _GEN_2035; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2037 = 7'h3c == total_offset_35[6:0] ? phv_data_60 : _GEN_2036; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2038 = 7'h3d == total_offset_35[6:0] ? phv_data_61 : _GEN_2037; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2039 = 7'h3e == total_offset_35[6:0] ? phv_data_62 : _GEN_2038; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2040 = 7'h3f == total_offset_35[6:0] ? phv_data_63 : _GEN_2039; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2041 = 7'h40 == total_offset_35[6:0] ? phv_data_64 : _GEN_2040; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2042 = 7'h41 == total_offset_35[6:0] ? phv_data_65 : _GEN_2041; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2043 = 7'h42 == total_offset_35[6:0] ? phv_data_66 : _GEN_2042; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2044 = 7'h43 == total_offset_35[6:0] ? phv_data_67 : _GEN_2043; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2045 = 7'h44 == total_offset_35[6:0] ? phv_data_68 : _GEN_2044; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2046 = 7'h45 == total_offset_35[6:0] ? phv_data_69 : _GEN_2045; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2047 = 7'h46 == total_offset_35[6:0] ? phv_data_70 : _GEN_2046; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2048 = 7'h47 == total_offset_35[6:0] ? phv_data_71 : _GEN_2047; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2049 = 7'h48 == total_offset_35[6:0] ? phv_data_72 : _GEN_2048; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2050 = 7'h49 == total_offset_35[6:0] ? phv_data_73 : _GEN_2049; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2051 = 7'h4a == total_offset_35[6:0] ? phv_data_74 : _GEN_2050; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2052 = 7'h4b == total_offset_35[6:0] ? phv_data_75 : _GEN_2051; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2053 = 7'h4c == total_offset_35[6:0] ? phv_data_76 : _GEN_2052; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2054 = 7'h4d == total_offset_35[6:0] ? phv_data_77 : _GEN_2053; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2055 = 7'h4e == total_offset_35[6:0] ? phv_data_78 : _GEN_2054; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2056 = 7'h4f == total_offset_35[6:0] ? phv_data_79 : _GEN_2055; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2057 = 7'h50 == total_offset_35[6:0] ? phv_data_80 : _GEN_2056; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2058 = 7'h51 == total_offset_35[6:0] ? phv_data_81 : _GEN_2057; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2059 = 7'h52 == total_offset_35[6:0] ? phv_data_82 : _GEN_2058; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2060 = 7'h53 == total_offset_35[6:0] ? phv_data_83 : _GEN_2059; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2061 = 7'h54 == total_offset_35[6:0] ? phv_data_84 : _GEN_2060; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2062 = 7'h55 == total_offset_35[6:0] ? phv_data_85 : _GEN_2061; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2063 = 7'h56 == total_offset_35[6:0] ? phv_data_86 : _GEN_2062; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2064 = 7'h57 == total_offset_35[6:0] ? phv_data_87 : _GEN_2063; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2065 = 7'h58 == total_offset_35[6:0] ? phv_data_88 : _GEN_2064; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2066 = 7'h59 == total_offset_35[6:0] ? phv_data_89 : _GEN_2065; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2067 = 7'h5a == total_offset_35[6:0] ? phv_data_90 : _GEN_2066; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2068 = 7'h5b == total_offset_35[6:0] ? phv_data_91 : _GEN_2067; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2069 = 7'h5c == total_offset_35[6:0] ? phv_data_92 : _GEN_2068; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2070 = 7'h5d == total_offset_35[6:0] ? phv_data_93 : _GEN_2069; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2071 = 7'h5e == total_offset_35[6:0] ? phv_data_94 : _GEN_2070; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2072 = 7'h5f == total_offset_35[6:0] ? phv_data_95 : _GEN_2071; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes_4_3 = 8'h3 < length_2 ? _GEN_2072 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_36 = offset_2 + 8'h4; // @[executor.scala 158:57]
  wire [7:0] _GEN_2075 = 7'h1 == total_offset_36[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2076 = 7'h2 == total_offset_36[6:0] ? phv_data_2 : _GEN_2075; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2077 = 7'h3 == total_offset_36[6:0] ? phv_data_3 : _GEN_2076; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2078 = 7'h4 == total_offset_36[6:0] ? phv_data_4 : _GEN_2077; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2079 = 7'h5 == total_offset_36[6:0] ? phv_data_5 : _GEN_2078; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2080 = 7'h6 == total_offset_36[6:0] ? phv_data_6 : _GEN_2079; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2081 = 7'h7 == total_offset_36[6:0] ? phv_data_7 : _GEN_2080; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2082 = 7'h8 == total_offset_36[6:0] ? phv_data_8 : _GEN_2081; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2083 = 7'h9 == total_offset_36[6:0] ? phv_data_9 : _GEN_2082; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2084 = 7'ha == total_offset_36[6:0] ? phv_data_10 : _GEN_2083; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2085 = 7'hb == total_offset_36[6:0] ? phv_data_11 : _GEN_2084; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2086 = 7'hc == total_offset_36[6:0] ? phv_data_12 : _GEN_2085; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2087 = 7'hd == total_offset_36[6:0] ? phv_data_13 : _GEN_2086; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2088 = 7'he == total_offset_36[6:0] ? phv_data_14 : _GEN_2087; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2089 = 7'hf == total_offset_36[6:0] ? phv_data_15 : _GEN_2088; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2090 = 7'h10 == total_offset_36[6:0] ? phv_data_16 : _GEN_2089; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2091 = 7'h11 == total_offset_36[6:0] ? phv_data_17 : _GEN_2090; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2092 = 7'h12 == total_offset_36[6:0] ? phv_data_18 : _GEN_2091; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2093 = 7'h13 == total_offset_36[6:0] ? phv_data_19 : _GEN_2092; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2094 = 7'h14 == total_offset_36[6:0] ? phv_data_20 : _GEN_2093; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2095 = 7'h15 == total_offset_36[6:0] ? phv_data_21 : _GEN_2094; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2096 = 7'h16 == total_offset_36[6:0] ? phv_data_22 : _GEN_2095; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2097 = 7'h17 == total_offset_36[6:0] ? phv_data_23 : _GEN_2096; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2098 = 7'h18 == total_offset_36[6:0] ? phv_data_24 : _GEN_2097; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2099 = 7'h19 == total_offset_36[6:0] ? phv_data_25 : _GEN_2098; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2100 = 7'h1a == total_offset_36[6:0] ? phv_data_26 : _GEN_2099; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2101 = 7'h1b == total_offset_36[6:0] ? phv_data_27 : _GEN_2100; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2102 = 7'h1c == total_offset_36[6:0] ? phv_data_28 : _GEN_2101; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2103 = 7'h1d == total_offset_36[6:0] ? phv_data_29 : _GEN_2102; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2104 = 7'h1e == total_offset_36[6:0] ? phv_data_30 : _GEN_2103; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2105 = 7'h1f == total_offset_36[6:0] ? phv_data_31 : _GEN_2104; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2106 = 7'h20 == total_offset_36[6:0] ? phv_data_32 : _GEN_2105; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2107 = 7'h21 == total_offset_36[6:0] ? phv_data_33 : _GEN_2106; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2108 = 7'h22 == total_offset_36[6:0] ? phv_data_34 : _GEN_2107; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2109 = 7'h23 == total_offset_36[6:0] ? phv_data_35 : _GEN_2108; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2110 = 7'h24 == total_offset_36[6:0] ? phv_data_36 : _GEN_2109; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2111 = 7'h25 == total_offset_36[6:0] ? phv_data_37 : _GEN_2110; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2112 = 7'h26 == total_offset_36[6:0] ? phv_data_38 : _GEN_2111; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2113 = 7'h27 == total_offset_36[6:0] ? phv_data_39 : _GEN_2112; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2114 = 7'h28 == total_offset_36[6:0] ? phv_data_40 : _GEN_2113; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2115 = 7'h29 == total_offset_36[6:0] ? phv_data_41 : _GEN_2114; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2116 = 7'h2a == total_offset_36[6:0] ? phv_data_42 : _GEN_2115; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2117 = 7'h2b == total_offset_36[6:0] ? phv_data_43 : _GEN_2116; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2118 = 7'h2c == total_offset_36[6:0] ? phv_data_44 : _GEN_2117; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2119 = 7'h2d == total_offset_36[6:0] ? phv_data_45 : _GEN_2118; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2120 = 7'h2e == total_offset_36[6:0] ? phv_data_46 : _GEN_2119; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2121 = 7'h2f == total_offset_36[6:0] ? phv_data_47 : _GEN_2120; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2122 = 7'h30 == total_offset_36[6:0] ? phv_data_48 : _GEN_2121; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2123 = 7'h31 == total_offset_36[6:0] ? phv_data_49 : _GEN_2122; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2124 = 7'h32 == total_offset_36[6:0] ? phv_data_50 : _GEN_2123; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2125 = 7'h33 == total_offset_36[6:0] ? phv_data_51 : _GEN_2124; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2126 = 7'h34 == total_offset_36[6:0] ? phv_data_52 : _GEN_2125; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2127 = 7'h35 == total_offset_36[6:0] ? phv_data_53 : _GEN_2126; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2128 = 7'h36 == total_offset_36[6:0] ? phv_data_54 : _GEN_2127; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2129 = 7'h37 == total_offset_36[6:0] ? phv_data_55 : _GEN_2128; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2130 = 7'h38 == total_offset_36[6:0] ? phv_data_56 : _GEN_2129; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2131 = 7'h39 == total_offset_36[6:0] ? phv_data_57 : _GEN_2130; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2132 = 7'h3a == total_offset_36[6:0] ? phv_data_58 : _GEN_2131; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2133 = 7'h3b == total_offset_36[6:0] ? phv_data_59 : _GEN_2132; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2134 = 7'h3c == total_offset_36[6:0] ? phv_data_60 : _GEN_2133; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2135 = 7'h3d == total_offset_36[6:0] ? phv_data_61 : _GEN_2134; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2136 = 7'h3e == total_offset_36[6:0] ? phv_data_62 : _GEN_2135; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2137 = 7'h3f == total_offset_36[6:0] ? phv_data_63 : _GEN_2136; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2138 = 7'h40 == total_offset_36[6:0] ? phv_data_64 : _GEN_2137; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2139 = 7'h41 == total_offset_36[6:0] ? phv_data_65 : _GEN_2138; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2140 = 7'h42 == total_offset_36[6:0] ? phv_data_66 : _GEN_2139; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2141 = 7'h43 == total_offset_36[6:0] ? phv_data_67 : _GEN_2140; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2142 = 7'h44 == total_offset_36[6:0] ? phv_data_68 : _GEN_2141; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2143 = 7'h45 == total_offset_36[6:0] ? phv_data_69 : _GEN_2142; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2144 = 7'h46 == total_offset_36[6:0] ? phv_data_70 : _GEN_2143; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2145 = 7'h47 == total_offset_36[6:0] ? phv_data_71 : _GEN_2144; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2146 = 7'h48 == total_offset_36[6:0] ? phv_data_72 : _GEN_2145; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2147 = 7'h49 == total_offset_36[6:0] ? phv_data_73 : _GEN_2146; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2148 = 7'h4a == total_offset_36[6:0] ? phv_data_74 : _GEN_2147; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2149 = 7'h4b == total_offset_36[6:0] ? phv_data_75 : _GEN_2148; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2150 = 7'h4c == total_offset_36[6:0] ? phv_data_76 : _GEN_2149; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2151 = 7'h4d == total_offset_36[6:0] ? phv_data_77 : _GEN_2150; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2152 = 7'h4e == total_offset_36[6:0] ? phv_data_78 : _GEN_2151; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2153 = 7'h4f == total_offset_36[6:0] ? phv_data_79 : _GEN_2152; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2154 = 7'h50 == total_offset_36[6:0] ? phv_data_80 : _GEN_2153; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2155 = 7'h51 == total_offset_36[6:0] ? phv_data_81 : _GEN_2154; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2156 = 7'h52 == total_offset_36[6:0] ? phv_data_82 : _GEN_2155; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2157 = 7'h53 == total_offset_36[6:0] ? phv_data_83 : _GEN_2156; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2158 = 7'h54 == total_offset_36[6:0] ? phv_data_84 : _GEN_2157; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2159 = 7'h55 == total_offset_36[6:0] ? phv_data_85 : _GEN_2158; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2160 = 7'h56 == total_offset_36[6:0] ? phv_data_86 : _GEN_2159; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2161 = 7'h57 == total_offset_36[6:0] ? phv_data_87 : _GEN_2160; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2162 = 7'h58 == total_offset_36[6:0] ? phv_data_88 : _GEN_2161; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2163 = 7'h59 == total_offset_36[6:0] ? phv_data_89 : _GEN_2162; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2164 = 7'h5a == total_offset_36[6:0] ? phv_data_90 : _GEN_2163; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2165 = 7'h5b == total_offset_36[6:0] ? phv_data_91 : _GEN_2164; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2166 = 7'h5c == total_offset_36[6:0] ? phv_data_92 : _GEN_2165; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2167 = 7'h5d == total_offset_36[6:0] ? phv_data_93 : _GEN_2166; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2168 = 7'h5e == total_offset_36[6:0] ? phv_data_94 : _GEN_2167; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2169 = 7'h5f == total_offset_36[6:0] ? phv_data_95 : _GEN_2168; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes_4_4 = 8'h4 < length_2 ? _GEN_2169 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_37 = offset_2 + 8'h5; // @[executor.scala 158:57]
  wire [7:0] _GEN_2172 = 7'h1 == total_offset_37[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2173 = 7'h2 == total_offset_37[6:0] ? phv_data_2 : _GEN_2172; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2174 = 7'h3 == total_offset_37[6:0] ? phv_data_3 : _GEN_2173; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2175 = 7'h4 == total_offset_37[6:0] ? phv_data_4 : _GEN_2174; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2176 = 7'h5 == total_offset_37[6:0] ? phv_data_5 : _GEN_2175; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2177 = 7'h6 == total_offset_37[6:0] ? phv_data_6 : _GEN_2176; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2178 = 7'h7 == total_offset_37[6:0] ? phv_data_7 : _GEN_2177; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2179 = 7'h8 == total_offset_37[6:0] ? phv_data_8 : _GEN_2178; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2180 = 7'h9 == total_offset_37[6:0] ? phv_data_9 : _GEN_2179; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2181 = 7'ha == total_offset_37[6:0] ? phv_data_10 : _GEN_2180; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2182 = 7'hb == total_offset_37[6:0] ? phv_data_11 : _GEN_2181; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2183 = 7'hc == total_offset_37[6:0] ? phv_data_12 : _GEN_2182; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2184 = 7'hd == total_offset_37[6:0] ? phv_data_13 : _GEN_2183; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2185 = 7'he == total_offset_37[6:0] ? phv_data_14 : _GEN_2184; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2186 = 7'hf == total_offset_37[6:0] ? phv_data_15 : _GEN_2185; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2187 = 7'h10 == total_offset_37[6:0] ? phv_data_16 : _GEN_2186; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2188 = 7'h11 == total_offset_37[6:0] ? phv_data_17 : _GEN_2187; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2189 = 7'h12 == total_offset_37[6:0] ? phv_data_18 : _GEN_2188; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2190 = 7'h13 == total_offset_37[6:0] ? phv_data_19 : _GEN_2189; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2191 = 7'h14 == total_offset_37[6:0] ? phv_data_20 : _GEN_2190; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2192 = 7'h15 == total_offset_37[6:0] ? phv_data_21 : _GEN_2191; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2193 = 7'h16 == total_offset_37[6:0] ? phv_data_22 : _GEN_2192; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2194 = 7'h17 == total_offset_37[6:0] ? phv_data_23 : _GEN_2193; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2195 = 7'h18 == total_offset_37[6:0] ? phv_data_24 : _GEN_2194; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2196 = 7'h19 == total_offset_37[6:0] ? phv_data_25 : _GEN_2195; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2197 = 7'h1a == total_offset_37[6:0] ? phv_data_26 : _GEN_2196; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2198 = 7'h1b == total_offset_37[6:0] ? phv_data_27 : _GEN_2197; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2199 = 7'h1c == total_offset_37[6:0] ? phv_data_28 : _GEN_2198; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2200 = 7'h1d == total_offset_37[6:0] ? phv_data_29 : _GEN_2199; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2201 = 7'h1e == total_offset_37[6:0] ? phv_data_30 : _GEN_2200; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2202 = 7'h1f == total_offset_37[6:0] ? phv_data_31 : _GEN_2201; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2203 = 7'h20 == total_offset_37[6:0] ? phv_data_32 : _GEN_2202; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2204 = 7'h21 == total_offset_37[6:0] ? phv_data_33 : _GEN_2203; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2205 = 7'h22 == total_offset_37[6:0] ? phv_data_34 : _GEN_2204; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2206 = 7'h23 == total_offset_37[6:0] ? phv_data_35 : _GEN_2205; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2207 = 7'h24 == total_offset_37[6:0] ? phv_data_36 : _GEN_2206; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2208 = 7'h25 == total_offset_37[6:0] ? phv_data_37 : _GEN_2207; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2209 = 7'h26 == total_offset_37[6:0] ? phv_data_38 : _GEN_2208; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2210 = 7'h27 == total_offset_37[6:0] ? phv_data_39 : _GEN_2209; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2211 = 7'h28 == total_offset_37[6:0] ? phv_data_40 : _GEN_2210; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2212 = 7'h29 == total_offset_37[6:0] ? phv_data_41 : _GEN_2211; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2213 = 7'h2a == total_offset_37[6:0] ? phv_data_42 : _GEN_2212; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2214 = 7'h2b == total_offset_37[6:0] ? phv_data_43 : _GEN_2213; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2215 = 7'h2c == total_offset_37[6:0] ? phv_data_44 : _GEN_2214; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2216 = 7'h2d == total_offset_37[6:0] ? phv_data_45 : _GEN_2215; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2217 = 7'h2e == total_offset_37[6:0] ? phv_data_46 : _GEN_2216; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2218 = 7'h2f == total_offset_37[6:0] ? phv_data_47 : _GEN_2217; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2219 = 7'h30 == total_offset_37[6:0] ? phv_data_48 : _GEN_2218; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2220 = 7'h31 == total_offset_37[6:0] ? phv_data_49 : _GEN_2219; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2221 = 7'h32 == total_offset_37[6:0] ? phv_data_50 : _GEN_2220; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2222 = 7'h33 == total_offset_37[6:0] ? phv_data_51 : _GEN_2221; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2223 = 7'h34 == total_offset_37[6:0] ? phv_data_52 : _GEN_2222; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2224 = 7'h35 == total_offset_37[6:0] ? phv_data_53 : _GEN_2223; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2225 = 7'h36 == total_offset_37[6:0] ? phv_data_54 : _GEN_2224; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2226 = 7'h37 == total_offset_37[6:0] ? phv_data_55 : _GEN_2225; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2227 = 7'h38 == total_offset_37[6:0] ? phv_data_56 : _GEN_2226; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2228 = 7'h39 == total_offset_37[6:0] ? phv_data_57 : _GEN_2227; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2229 = 7'h3a == total_offset_37[6:0] ? phv_data_58 : _GEN_2228; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2230 = 7'h3b == total_offset_37[6:0] ? phv_data_59 : _GEN_2229; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2231 = 7'h3c == total_offset_37[6:0] ? phv_data_60 : _GEN_2230; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2232 = 7'h3d == total_offset_37[6:0] ? phv_data_61 : _GEN_2231; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2233 = 7'h3e == total_offset_37[6:0] ? phv_data_62 : _GEN_2232; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2234 = 7'h3f == total_offset_37[6:0] ? phv_data_63 : _GEN_2233; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2235 = 7'h40 == total_offset_37[6:0] ? phv_data_64 : _GEN_2234; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2236 = 7'h41 == total_offset_37[6:0] ? phv_data_65 : _GEN_2235; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2237 = 7'h42 == total_offset_37[6:0] ? phv_data_66 : _GEN_2236; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2238 = 7'h43 == total_offset_37[6:0] ? phv_data_67 : _GEN_2237; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2239 = 7'h44 == total_offset_37[6:0] ? phv_data_68 : _GEN_2238; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2240 = 7'h45 == total_offset_37[6:0] ? phv_data_69 : _GEN_2239; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2241 = 7'h46 == total_offset_37[6:0] ? phv_data_70 : _GEN_2240; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2242 = 7'h47 == total_offset_37[6:0] ? phv_data_71 : _GEN_2241; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2243 = 7'h48 == total_offset_37[6:0] ? phv_data_72 : _GEN_2242; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2244 = 7'h49 == total_offset_37[6:0] ? phv_data_73 : _GEN_2243; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2245 = 7'h4a == total_offset_37[6:0] ? phv_data_74 : _GEN_2244; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2246 = 7'h4b == total_offset_37[6:0] ? phv_data_75 : _GEN_2245; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2247 = 7'h4c == total_offset_37[6:0] ? phv_data_76 : _GEN_2246; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2248 = 7'h4d == total_offset_37[6:0] ? phv_data_77 : _GEN_2247; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2249 = 7'h4e == total_offset_37[6:0] ? phv_data_78 : _GEN_2248; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2250 = 7'h4f == total_offset_37[6:0] ? phv_data_79 : _GEN_2249; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2251 = 7'h50 == total_offset_37[6:0] ? phv_data_80 : _GEN_2250; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2252 = 7'h51 == total_offset_37[6:0] ? phv_data_81 : _GEN_2251; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2253 = 7'h52 == total_offset_37[6:0] ? phv_data_82 : _GEN_2252; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2254 = 7'h53 == total_offset_37[6:0] ? phv_data_83 : _GEN_2253; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2255 = 7'h54 == total_offset_37[6:0] ? phv_data_84 : _GEN_2254; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2256 = 7'h55 == total_offset_37[6:0] ? phv_data_85 : _GEN_2255; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2257 = 7'h56 == total_offset_37[6:0] ? phv_data_86 : _GEN_2256; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2258 = 7'h57 == total_offset_37[6:0] ? phv_data_87 : _GEN_2257; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2259 = 7'h58 == total_offset_37[6:0] ? phv_data_88 : _GEN_2258; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2260 = 7'h59 == total_offset_37[6:0] ? phv_data_89 : _GEN_2259; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2261 = 7'h5a == total_offset_37[6:0] ? phv_data_90 : _GEN_2260; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2262 = 7'h5b == total_offset_37[6:0] ? phv_data_91 : _GEN_2261; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2263 = 7'h5c == total_offset_37[6:0] ? phv_data_92 : _GEN_2262; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2264 = 7'h5d == total_offset_37[6:0] ? phv_data_93 : _GEN_2263; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2265 = 7'h5e == total_offset_37[6:0] ? phv_data_94 : _GEN_2264; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2266 = 7'h5f == total_offset_37[6:0] ? phv_data_95 : _GEN_2265; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes_4_5 = 8'h5 < length_2 ? _GEN_2266 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_38 = offset_2 + 8'h6; // @[executor.scala 158:57]
  wire [7:0] _GEN_2269 = 7'h1 == total_offset_38[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2270 = 7'h2 == total_offset_38[6:0] ? phv_data_2 : _GEN_2269; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2271 = 7'h3 == total_offset_38[6:0] ? phv_data_3 : _GEN_2270; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2272 = 7'h4 == total_offset_38[6:0] ? phv_data_4 : _GEN_2271; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2273 = 7'h5 == total_offset_38[6:0] ? phv_data_5 : _GEN_2272; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2274 = 7'h6 == total_offset_38[6:0] ? phv_data_6 : _GEN_2273; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2275 = 7'h7 == total_offset_38[6:0] ? phv_data_7 : _GEN_2274; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2276 = 7'h8 == total_offset_38[6:0] ? phv_data_8 : _GEN_2275; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2277 = 7'h9 == total_offset_38[6:0] ? phv_data_9 : _GEN_2276; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2278 = 7'ha == total_offset_38[6:0] ? phv_data_10 : _GEN_2277; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2279 = 7'hb == total_offset_38[6:0] ? phv_data_11 : _GEN_2278; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2280 = 7'hc == total_offset_38[6:0] ? phv_data_12 : _GEN_2279; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2281 = 7'hd == total_offset_38[6:0] ? phv_data_13 : _GEN_2280; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2282 = 7'he == total_offset_38[6:0] ? phv_data_14 : _GEN_2281; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2283 = 7'hf == total_offset_38[6:0] ? phv_data_15 : _GEN_2282; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2284 = 7'h10 == total_offset_38[6:0] ? phv_data_16 : _GEN_2283; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2285 = 7'h11 == total_offset_38[6:0] ? phv_data_17 : _GEN_2284; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2286 = 7'h12 == total_offset_38[6:0] ? phv_data_18 : _GEN_2285; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2287 = 7'h13 == total_offset_38[6:0] ? phv_data_19 : _GEN_2286; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2288 = 7'h14 == total_offset_38[6:0] ? phv_data_20 : _GEN_2287; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2289 = 7'h15 == total_offset_38[6:0] ? phv_data_21 : _GEN_2288; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2290 = 7'h16 == total_offset_38[6:0] ? phv_data_22 : _GEN_2289; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2291 = 7'h17 == total_offset_38[6:0] ? phv_data_23 : _GEN_2290; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2292 = 7'h18 == total_offset_38[6:0] ? phv_data_24 : _GEN_2291; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2293 = 7'h19 == total_offset_38[6:0] ? phv_data_25 : _GEN_2292; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2294 = 7'h1a == total_offset_38[6:0] ? phv_data_26 : _GEN_2293; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2295 = 7'h1b == total_offset_38[6:0] ? phv_data_27 : _GEN_2294; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2296 = 7'h1c == total_offset_38[6:0] ? phv_data_28 : _GEN_2295; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2297 = 7'h1d == total_offset_38[6:0] ? phv_data_29 : _GEN_2296; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2298 = 7'h1e == total_offset_38[6:0] ? phv_data_30 : _GEN_2297; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2299 = 7'h1f == total_offset_38[6:0] ? phv_data_31 : _GEN_2298; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2300 = 7'h20 == total_offset_38[6:0] ? phv_data_32 : _GEN_2299; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2301 = 7'h21 == total_offset_38[6:0] ? phv_data_33 : _GEN_2300; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2302 = 7'h22 == total_offset_38[6:0] ? phv_data_34 : _GEN_2301; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2303 = 7'h23 == total_offset_38[6:0] ? phv_data_35 : _GEN_2302; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2304 = 7'h24 == total_offset_38[6:0] ? phv_data_36 : _GEN_2303; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2305 = 7'h25 == total_offset_38[6:0] ? phv_data_37 : _GEN_2304; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2306 = 7'h26 == total_offset_38[6:0] ? phv_data_38 : _GEN_2305; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2307 = 7'h27 == total_offset_38[6:0] ? phv_data_39 : _GEN_2306; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2308 = 7'h28 == total_offset_38[6:0] ? phv_data_40 : _GEN_2307; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2309 = 7'h29 == total_offset_38[6:0] ? phv_data_41 : _GEN_2308; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2310 = 7'h2a == total_offset_38[6:0] ? phv_data_42 : _GEN_2309; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2311 = 7'h2b == total_offset_38[6:0] ? phv_data_43 : _GEN_2310; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2312 = 7'h2c == total_offset_38[6:0] ? phv_data_44 : _GEN_2311; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2313 = 7'h2d == total_offset_38[6:0] ? phv_data_45 : _GEN_2312; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2314 = 7'h2e == total_offset_38[6:0] ? phv_data_46 : _GEN_2313; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2315 = 7'h2f == total_offset_38[6:0] ? phv_data_47 : _GEN_2314; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2316 = 7'h30 == total_offset_38[6:0] ? phv_data_48 : _GEN_2315; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2317 = 7'h31 == total_offset_38[6:0] ? phv_data_49 : _GEN_2316; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2318 = 7'h32 == total_offset_38[6:0] ? phv_data_50 : _GEN_2317; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2319 = 7'h33 == total_offset_38[6:0] ? phv_data_51 : _GEN_2318; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2320 = 7'h34 == total_offset_38[6:0] ? phv_data_52 : _GEN_2319; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2321 = 7'h35 == total_offset_38[6:0] ? phv_data_53 : _GEN_2320; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2322 = 7'h36 == total_offset_38[6:0] ? phv_data_54 : _GEN_2321; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2323 = 7'h37 == total_offset_38[6:0] ? phv_data_55 : _GEN_2322; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2324 = 7'h38 == total_offset_38[6:0] ? phv_data_56 : _GEN_2323; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2325 = 7'h39 == total_offset_38[6:0] ? phv_data_57 : _GEN_2324; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2326 = 7'h3a == total_offset_38[6:0] ? phv_data_58 : _GEN_2325; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2327 = 7'h3b == total_offset_38[6:0] ? phv_data_59 : _GEN_2326; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2328 = 7'h3c == total_offset_38[6:0] ? phv_data_60 : _GEN_2327; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2329 = 7'h3d == total_offset_38[6:0] ? phv_data_61 : _GEN_2328; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2330 = 7'h3e == total_offset_38[6:0] ? phv_data_62 : _GEN_2329; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2331 = 7'h3f == total_offset_38[6:0] ? phv_data_63 : _GEN_2330; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2332 = 7'h40 == total_offset_38[6:0] ? phv_data_64 : _GEN_2331; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2333 = 7'h41 == total_offset_38[6:0] ? phv_data_65 : _GEN_2332; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2334 = 7'h42 == total_offset_38[6:0] ? phv_data_66 : _GEN_2333; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2335 = 7'h43 == total_offset_38[6:0] ? phv_data_67 : _GEN_2334; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2336 = 7'h44 == total_offset_38[6:0] ? phv_data_68 : _GEN_2335; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2337 = 7'h45 == total_offset_38[6:0] ? phv_data_69 : _GEN_2336; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2338 = 7'h46 == total_offset_38[6:0] ? phv_data_70 : _GEN_2337; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2339 = 7'h47 == total_offset_38[6:0] ? phv_data_71 : _GEN_2338; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2340 = 7'h48 == total_offset_38[6:0] ? phv_data_72 : _GEN_2339; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2341 = 7'h49 == total_offset_38[6:0] ? phv_data_73 : _GEN_2340; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2342 = 7'h4a == total_offset_38[6:0] ? phv_data_74 : _GEN_2341; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2343 = 7'h4b == total_offset_38[6:0] ? phv_data_75 : _GEN_2342; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2344 = 7'h4c == total_offset_38[6:0] ? phv_data_76 : _GEN_2343; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2345 = 7'h4d == total_offset_38[6:0] ? phv_data_77 : _GEN_2344; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2346 = 7'h4e == total_offset_38[6:0] ? phv_data_78 : _GEN_2345; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2347 = 7'h4f == total_offset_38[6:0] ? phv_data_79 : _GEN_2346; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2348 = 7'h50 == total_offset_38[6:0] ? phv_data_80 : _GEN_2347; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2349 = 7'h51 == total_offset_38[6:0] ? phv_data_81 : _GEN_2348; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2350 = 7'h52 == total_offset_38[6:0] ? phv_data_82 : _GEN_2349; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2351 = 7'h53 == total_offset_38[6:0] ? phv_data_83 : _GEN_2350; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2352 = 7'h54 == total_offset_38[6:0] ? phv_data_84 : _GEN_2351; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2353 = 7'h55 == total_offset_38[6:0] ? phv_data_85 : _GEN_2352; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2354 = 7'h56 == total_offset_38[6:0] ? phv_data_86 : _GEN_2353; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2355 = 7'h57 == total_offset_38[6:0] ? phv_data_87 : _GEN_2354; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2356 = 7'h58 == total_offset_38[6:0] ? phv_data_88 : _GEN_2355; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2357 = 7'h59 == total_offset_38[6:0] ? phv_data_89 : _GEN_2356; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2358 = 7'h5a == total_offset_38[6:0] ? phv_data_90 : _GEN_2357; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2359 = 7'h5b == total_offset_38[6:0] ? phv_data_91 : _GEN_2358; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2360 = 7'h5c == total_offset_38[6:0] ? phv_data_92 : _GEN_2359; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2361 = 7'h5d == total_offset_38[6:0] ? phv_data_93 : _GEN_2360; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2362 = 7'h5e == total_offset_38[6:0] ? phv_data_94 : _GEN_2361; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2363 = 7'h5f == total_offset_38[6:0] ? phv_data_95 : _GEN_2362; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes_4_6 = 8'h6 < length_2 ? _GEN_2363 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_39 = offset_2 + 8'h7; // @[executor.scala 158:57]
  wire [7:0] _GEN_2366 = 7'h1 == total_offset_39[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2367 = 7'h2 == total_offset_39[6:0] ? phv_data_2 : _GEN_2366; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2368 = 7'h3 == total_offset_39[6:0] ? phv_data_3 : _GEN_2367; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2369 = 7'h4 == total_offset_39[6:0] ? phv_data_4 : _GEN_2368; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2370 = 7'h5 == total_offset_39[6:0] ? phv_data_5 : _GEN_2369; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2371 = 7'h6 == total_offset_39[6:0] ? phv_data_6 : _GEN_2370; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2372 = 7'h7 == total_offset_39[6:0] ? phv_data_7 : _GEN_2371; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2373 = 7'h8 == total_offset_39[6:0] ? phv_data_8 : _GEN_2372; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2374 = 7'h9 == total_offset_39[6:0] ? phv_data_9 : _GEN_2373; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2375 = 7'ha == total_offset_39[6:0] ? phv_data_10 : _GEN_2374; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2376 = 7'hb == total_offset_39[6:0] ? phv_data_11 : _GEN_2375; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2377 = 7'hc == total_offset_39[6:0] ? phv_data_12 : _GEN_2376; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2378 = 7'hd == total_offset_39[6:0] ? phv_data_13 : _GEN_2377; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2379 = 7'he == total_offset_39[6:0] ? phv_data_14 : _GEN_2378; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2380 = 7'hf == total_offset_39[6:0] ? phv_data_15 : _GEN_2379; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2381 = 7'h10 == total_offset_39[6:0] ? phv_data_16 : _GEN_2380; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2382 = 7'h11 == total_offset_39[6:0] ? phv_data_17 : _GEN_2381; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2383 = 7'h12 == total_offset_39[6:0] ? phv_data_18 : _GEN_2382; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2384 = 7'h13 == total_offset_39[6:0] ? phv_data_19 : _GEN_2383; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2385 = 7'h14 == total_offset_39[6:0] ? phv_data_20 : _GEN_2384; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2386 = 7'h15 == total_offset_39[6:0] ? phv_data_21 : _GEN_2385; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2387 = 7'h16 == total_offset_39[6:0] ? phv_data_22 : _GEN_2386; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2388 = 7'h17 == total_offset_39[6:0] ? phv_data_23 : _GEN_2387; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2389 = 7'h18 == total_offset_39[6:0] ? phv_data_24 : _GEN_2388; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2390 = 7'h19 == total_offset_39[6:0] ? phv_data_25 : _GEN_2389; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2391 = 7'h1a == total_offset_39[6:0] ? phv_data_26 : _GEN_2390; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2392 = 7'h1b == total_offset_39[6:0] ? phv_data_27 : _GEN_2391; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2393 = 7'h1c == total_offset_39[6:0] ? phv_data_28 : _GEN_2392; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2394 = 7'h1d == total_offset_39[6:0] ? phv_data_29 : _GEN_2393; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2395 = 7'h1e == total_offset_39[6:0] ? phv_data_30 : _GEN_2394; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2396 = 7'h1f == total_offset_39[6:0] ? phv_data_31 : _GEN_2395; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2397 = 7'h20 == total_offset_39[6:0] ? phv_data_32 : _GEN_2396; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2398 = 7'h21 == total_offset_39[6:0] ? phv_data_33 : _GEN_2397; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2399 = 7'h22 == total_offset_39[6:0] ? phv_data_34 : _GEN_2398; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2400 = 7'h23 == total_offset_39[6:0] ? phv_data_35 : _GEN_2399; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2401 = 7'h24 == total_offset_39[6:0] ? phv_data_36 : _GEN_2400; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2402 = 7'h25 == total_offset_39[6:0] ? phv_data_37 : _GEN_2401; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2403 = 7'h26 == total_offset_39[6:0] ? phv_data_38 : _GEN_2402; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2404 = 7'h27 == total_offset_39[6:0] ? phv_data_39 : _GEN_2403; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2405 = 7'h28 == total_offset_39[6:0] ? phv_data_40 : _GEN_2404; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2406 = 7'h29 == total_offset_39[6:0] ? phv_data_41 : _GEN_2405; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2407 = 7'h2a == total_offset_39[6:0] ? phv_data_42 : _GEN_2406; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2408 = 7'h2b == total_offset_39[6:0] ? phv_data_43 : _GEN_2407; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2409 = 7'h2c == total_offset_39[6:0] ? phv_data_44 : _GEN_2408; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2410 = 7'h2d == total_offset_39[6:0] ? phv_data_45 : _GEN_2409; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2411 = 7'h2e == total_offset_39[6:0] ? phv_data_46 : _GEN_2410; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2412 = 7'h2f == total_offset_39[6:0] ? phv_data_47 : _GEN_2411; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2413 = 7'h30 == total_offset_39[6:0] ? phv_data_48 : _GEN_2412; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2414 = 7'h31 == total_offset_39[6:0] ? phv_data_49 : _GEN_2413; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2415 = 7'h32 == total_offset_39[6:0] ? phv_data_50 : _GEN_2414; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2416 = 7'h33 == total_offset_39[6:0] ? phv_data_51 : _GEN_2415; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2417 = 7'h34 == total_offset_39[6:0] ? phv_data_52 : _GEN_2416; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2418 = 7'h35 == total_offset_39[6:0] ? phv_data_53 : _GEN_2417; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2419 = 7'h36 == total_offset_39[6:0] ? phv_data_54 : _GEN_2418; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2420 = 7'h37 == total_offset_39[6:0] ? phv_data_55 : _GEN_2419; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2421 = 7'h38 == total_offset_39[6:0] ? phv_data_56 : _GEN_2420; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2422 = 7'h39 == total_offset_39[6:0] ? phv_data_57 : _GEN_2421; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2423 = 7'h3a == total_offset_39[6:0] ? phv_data_58 : _GEN_2422; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2424 = 7'h3b == total_offset_39[6:0] ? phv_data_59 : _GEN_2423; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2425 = 7'h3c == total_offset_39[6:0] ? phv_data_60 : _GEN_2424; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2426 = 7'h3d == total_offset_39[6:0] ? phv_data_61 : _GEN_2425; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2427 = 7'h3e == total_offset_39[6:0] ? phv_data_62 : _GEN_2426; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2428 = 7'h3f == total_offset_39[6:0] ? phv_data_63 : _GEN_2427; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2429 = 7'h40 == total_offset_39[6:0] ? phv_data_64 : _GEN_2428; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2430 = 7'h41 == total_offset_39[6:0] ? phv_data_65 : _GEN_2429; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2431 = 7'h42 == total_offset_39[6:0] ? phv_data_66 : _GEN_2430; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2432 = 7'h43 == total_offset_39[6:0] ? phv_data_67 : _GEN_2431; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2433 = 7'h44 == total_offset_39[6:0] ? phv_data_68 : _GEN_2432; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2434 = 7'h45 == total_offset_39[6:0] ? phv_data_69 : _GEN_2433; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2435 = 7'h46 == total_offset_39[6:0] ? phv_data_70 : _GEN_2434; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2436 = 7'h47 == total_offset_39[6:0] ? phv_data_71 : _GEN_2435; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2437 = 7'h48 == total_offset_39[6:0] ? phv_data_72 : _GEN_2436; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2438 = 7'h49 == total_offset_39[6:0] ? phv_data_73 : _GEN_2437; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2439 = 7'h4a == total_offset_39[6:0] ? phv_data_74 : _GEN_2438; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2440 = 7'h4b == total_offset_39[6:0] ? phv_data_75 : _GEN_2439; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2441 = 7'h4c == total_offset_39[6:0] ? phv_data_76 : _GEN_2440; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2442 = 7'h4d == total_offset_39[6:0] ? phv_data_77 : _GEN_2441; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2443 = 7'h4e == total_offset_39[6:0] ? phv_data_78 : _GEN_2442; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2444 = 7'h4f == total_offset_39[6:0] ? phv_data_79 : _GEN_2443; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2445 = 7'h50 == total_offset_39[6:0] ? phv_data_80 : _GEN_2444; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2446 = 7'h51 == total_offset_39[6:0] ? phv_data_81 : _GEN_2445; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2447 = 7'h52 == total_offset_39[6:0] ? phv_data_82 : _GEN_2446; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2448 = 7'h53 == total_offset_39[6:0] ? phv_data_83 : _GEN_2447; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2449 = 7'h54 == total_offset_39[6:0] ? phv_data_84 : _GEN_2448; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2450 = 7'h55 == total_offset_39[6:0] ? phv_data_85 : _GEN_2449; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2451 = 7'h56 == total_offset_39[6:0] ? phv_data_86 : _GEN_2450; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2452 = 7'h57 == total_offset_39[6:0] ? phv_data_87 : _GEN_2451; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2453 = 7'h58 == total_offset_39[6:0] ? phv_data_88 : _GEN_2452; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2454 = 7'h59 == total_offset_39[6:0] ? phv_data_89 : _GEN_2453; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2455 = 7'h5a == total_offset_39[6:0] ? phv_data_90 : _GEN_2454; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2456 = 7'h5b == total_offset_39[6:0] ? phv_data_91 : _GEN_2455; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2457 = 7'h5c == total_offset_39[6:0] ? phv_data_92 : _GEN_2456; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2458 = 7'h5d == total_offset_39[6:0] ? phv_data_93 : _GEN_2457; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2459 = 7'h5e == total_offset_39[6:0] ? phv_data_94 : _GEN_2458; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2460 = 7'h5f == total_offset_39[6:0] ? phv_data_95 : _GEN_2459; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes_4_7 = 8'h7 < length_2 ? _GEN_2460 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [63:0] _io_field_out_2_T = {bytes_4_0,bytes_4_1,bytes_4_2,bytes_4_3,bytes_4_4,bytes_4_5,bytes_4_6,bytes_4_7}; // @[Cat.scala 30:58]
  wire [2:0] args_offset_2 = io_field_out_2_lo[13:11]; // @[primitive.scala 34:52]
  wire [2:0] args_length_2 = io_field_out_2_lo[10:8]; // @[primitive.scala 35:52]
  wire [8:0] _total_offset_T_40 = {{6'd0}, args_offset_2}; // @[executor.scala 173:60]
  wire [7:0] total_offset_40 = _total_offset_T_40[7:0]; // @[executor.scala 173:60]
  wire [7:0] _GEN_3400 = {{5'd0}, args_length_2}; // @[executor.scala 174:48]
  wire [7:0] _GEN_2463 = 3'h1 == total_offset_40[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2464 = 3'h2 == total_offset_40[2:0] ? args_2 : _GEN_2463; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2465 = 3'h3 == total_offset_40[2:0] ? args_3 : _GEN_2464; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2466 = 3'h4 == total_offset_40[2:0] ? args_4 : _GEN_2465; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2467 = 3'h5 == total_offset_40[2:0] ? args_5 : _GEN_2466; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2468 = 3'h6 == total_offset_40[2:0] ? args_6 : _GEN_2467; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_5_0 = 8'h0 < _GEN_3400 ? _GEN_2468 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [7:0] _GEN_3401 = {{5'd0}, args_offset_2}; // @[executor.scala 173:60]
  wire [7:0] total_offset_41 = _GEN_3401 + 8'h1; // @[executor.scala 173:60]
  wire [7:0] _GEN_2471 = 3'h1 == total_offset_41[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2472 = 3'h2 == total_offset_41[2:0] ? args_2 : _GEN_2471; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2473 = 3'h3 == total_offset_41[2:0] ? args_3 : _GEN_2472; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2474 = 3'h4 == total_offset_41[2:0] ? args_4 : _GEN_2473; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2475 = 3'h5 == total_offset_41[2:0] ? args_5 : _GEN_2474; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2476 = 3'h6 == total_offset_41[2:0] ? args_6 : _GEN_2475; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_5_1 = 8'h1 < _GEN_3400 ? _GEN_2476 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [7:0] total_offset_42 = _GEN_3401 + 8'h2; // @[executor.scala 173:60]
  wire [7:0] _GEN_2479 = 3'h1 == total_offset_42[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2480 = 3'h2 == total_offset_42[2:0] ? args_2 : _GEN_2479; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2481 = 3'h3 == total_offset_42[2:0] ? args_3 : _GEN_2480; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2482 = 3'h4 == total_offset_42[2:0] ? args_4 : _GEN_2481; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2483 = 3'h5 == total_offset_42[2:0] ? args_5 : _GEN_2482; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2484 = 3'h6 == total_offset_42[2:0] ? args_6 : _GEN_2483; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_5_2 = 8'h2 < _GEN_3400 ? _GEN_2484 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [7:0] total_offset_43 = _GEN_3401 + 8'h3; // @[executor.scala 173:60]
  wire [7:0] _GEN_2487 = 3'h1 == total_offset_43[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2488 = 3'h2 == total_offset_43[2:0] ? args_2 : _GEN_2487; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2489 = 3'h3 == total_offset_43[2:0] ? args_3 : _GEN_2488; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2490 = 3'h4 == total_offset_43[2:0] ? args_4 : _GEN_2489; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2491 = 3'h5 == total_offset_43[2:0] ? args_5 : _GEN_2490; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2492 = 3'h6 == total_offset_43[2:0] ? args_6 : _GEN_2491; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_5_3 = 8'h3 < _GEN_3400 ? _GEN_2492 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [7:0] total_offset_44 = _GEN_3401 + 8'h4; // @[executor.scala 173:60]
  wire [7:0] _GEN_2495 = 3'h1 == total_offset_44[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2496 = 3'h2 == total_offset_44[2:0] ? args_2 : _GEN_2495; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2497 = 3'h3 == total_offset_44[2:0] ? args_3 : _GEN_2496; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2498 = 3'h4 == total_offset_44[2:0] ? args_4 : _GEN_2497; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2499 = 3'h5 == total_offset_44[2:0] ? args_5 : _GEN_2498; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2500 = 3'h6 == total_offset_44[2:0] ? args_6 : _GEN_2499; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_5_4 = 8'h4 < _GEN_3400 ? _GEN_2500 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [7:0] total_offset_45 = _GEN_3401 + 8'h5; // @[executor.scala 173:60]
  wire [7:0] _GEN_2503 = 3'h1 == total_offset_45[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2504 = 3'h2 == total_offset_45[2:0] ? args_2 : _GEN_2503; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2505 = 3'h3 == total_offset_45[2:0] ? args_3 : _GEN_2504; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2506 = 3'h4 == total_offset_45[2:0] ? args_4 : _GEN_2505; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2507 = 3'h5 == total_offset_45[2:0] ? args_5 : _GEN_2506; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2508 = 3'h6 == total_offset_45[2:0] ? args_6 : _GEN_2507; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_5_5 = 8'h5 < _GEN_3400 ? _GEN_2508 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [7:0] total_offset_46 = _GEN_3401 + 8'h6; // @[executor.scala 173:60]
  wire [7:0] _GEN_2511 = 3'h1 == total_offset_46[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2512 = 3'h2 == total_offset_46[2:0] ? args_2 : _GEN_2511; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2513 = 3'h3 == total_offset_46[2:0] ? args_3 : _GEN_2512; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2514 = 3'h4 == total_offset_46[2:0] ? args_4 : _GEN_2513; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2515 = 3'h5 == total_offset_46[2:0] ? args_5 : _GEN_2514; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_2516 = 3'h6 == total_offset_46[2:0] ? args_6 : _GEN_2515; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_5_6 = 8'h6 < _GEN_3400 ? _GEN_2516 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [63:0] _io_field_out_2_T_1 = {bytes_5_0,bytes_5_1,bytes_5_2,bytes_5_3,bytes_5_4,bytes_5_5,bytes_5_6,8'h0}; // @[Cat.scala 30:58]
  wire [49:0] io_field_out_2_hi_12 = io_field_out_2_lo[13] ? 50'h3ffffffffffff : 50'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _io_field_out_2_T_4 = {io_field_out_2_hi_12,io_field_out_2_lo}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_2526 = 4'ha == opcode_2 ? _io_field_out_2_T_1 : _io_field_out_2_T_4; // @[executor.scala 167:55 executor.scala 180:41 executor.scala 183:41]
  wire [63:0] _GEN_2527 = from_header_2 ? _io_field_out_2_T : _GEN_2526; // @[executor.scala 152:36 executor.scala 165:37]
  wire [3:0] opcode_3 = vliw_3[31:28]; // @[primitive.scala 9:44]
  wire [13:0] io_field_out_3_lo = vliw_3[13:0]; // @[primitive.scala 11:44]
  wire  from_header_3 = length_3 != 8'h0; // @[executor.scala 151:45]
  wire [8:0] _total_offset_T_48 = {{1'd0}, offset_3}; // @[executor.scala 158:57]
  wire [7:0] total_offset_48 = _total_offset_T_48[7:0]; // @[executor.scala 158:57]
  wire [7:0] _GEN_2530 = 7'h1 == total_offset_48[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2531 = 7'h2 == total_offset_48[6:0] ? phv_data_2 : _GEN_2530; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2532 = 7'h3 == total_offset_48[6:0] ? phv_data_3 : _GEN_2531; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2533 = 7'h4 == total_offset_48[6:0] ? phv_data_4 : _GEN_2532; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2534 = 7'h5 == total_offset_48[6:0] ? phv_data_5 : _GEN_2533; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2535 = 7'h6 == total_offset_48[6:0] ? phv_data_6 : _GEN_2534; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2536 = 7'h7 == total_offset_48[6:0] ? phv_data_7 : _GEN_2535; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2537 = 7'h8 == total_offset_48[6:0] ? phv_data_8 : _GEN_2536; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2538 = 7'h9 == total_offset_48[6:0] ? phv_data_9 : _GEN_2537; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2539 = 7'ha == total_offset_48[6:0] ? phv_data_10 : _GEN_2538; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2540 = 7'hb == total_offset_48[6:0] ? phv_data_11 : _GEN_2539; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2541 = 7'hc == total_offset_48[6:0] ? phv_data_12 : _GEN_2540; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2542 = 7'hd == total_offset_48[6:0] ? phv_data_13 : _GEN_2541; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2543 = 7'he == total_offset_48[6:0] ? phv_data_14 : _GEN_2542; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2544 = 7'hf == total_offset_48[6:0] ? phv_data_15 : _GEN_2543; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2545 = 7'h10 == total_offset_48[6:0] ? phv_data_16 : _GEN_2544; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2546 = 7'h11 == total_offset_48[6:0] ? phv_data_17 : _GEN_2545; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2547 = 7'h12 == total_offset_48[6:0] ? phv_data_18 : _GEN_2546; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2548 = 7'h13 == total_offset_48[6:0] ? phv_data_19 : _GEN_2547; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2549 = 7'h14 == total_offset_48[6:0] ? phv_data_20 : _GEN_2548; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2550 = 7'h15 == total_offset_48[6:0] ? phv_data_21 : _GEN_2549; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2551 = 7'h16 == total_offset_48[6:0] ? phv_data_22 : _GEN_2550; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2552 = 7'h17 == total_offset_48[6:0] ? phv_data_23 : _GEN_2551; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2553 = 7'h18 == total_offset_48[6:0] ? phv_data_24 : _GEN_2552; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2554 = 7'h19 == total_offset_48[6:0] ? phv_data_25 : _GEN_2553; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2555 = 7'h1a == total_offset_48[6:0] ? phv_data_26 : _GEN_2554; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2556 = 7'h1b == total_offset_48[6:0] ? phv_data_27 : _GEN_2555; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2557 = 7'h1c == total_offset_48[6:0] ? phv_data_28 : _GEN_2556; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2558 = 7'h1d == total_offset_48[6:0] ? phv_data_29 : _GEN_2557; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2559 = 7'h1e == total_offset_48[6:0] ? phv_data_30 : _GEN_2558; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2560 = 7'h1f == total_offset_48[6:0] ? phv_data_31 : _GEN_2559; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2561 = 7'h20 == total_offset_48[6:0] ? phv_data_32 : _GEN_2560; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2562 = 7'h21 == total_offset_48[6:0] ? phv_data_33 : _GEN_2561; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2563 = 7'h22 == total_offset_48[6:0] ? phv_data_34 : _GEN_2562; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2564 = 7'h23 == total_offset_48[6:0] ? phv_data_35 : _GEN_2563; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2565 = 7'h24 == total_offset_48[6:0] ? phv_data_36 : _GEN_2564; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2566 = 7'h25 == total_offset_48[6:0] ? phv_data_37 : _GEN_2565; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2567 = 7'h26 == total_offset_48[6:0] ? phv_data_38 : _GEN_2566; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2568 = 7'h27 == total_offset_48[6:0] ? phv_data_39 : _GEN_2567; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2569 = 7'h28 == total_offset_48[6:0] ? phv_data_40 : _GEN_2568; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2570 = 7'h29 == total_offset_48[6:0] ? phv_data_41 : _GEN_2569; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2571 = 7'h2a == total_offset_48[6:0] ? phv_data_42 : _GEN_2570; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2572 = 7'h2b == total_offset_48[6:0] ? phv_data_43 : _GEN_2571; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2573 = 7'h2c == total_offset_48[6:0] ? phv_data_44 : _GEN_2572; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2574 = 7'h2d == total_offset_48[6:0] ? phv_data_45 : _GEN_2573; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2575 = 7'h2e == total_offset_48[6:0] ? phv_data_46 : _GEN_2574; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2576 = 7'h2f == total_offset_48[6:0] ? phv_data_47 : _GEN_2575; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2577 = 7'h30 == total_offset_48[6:0] ? phv_data_48 : _GEN_2576; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2578 = 7'h31 == total_offset_48[6:0] ? phv_data_49 : _GEN_2577; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2579 = 7'h32 == total_offset_48[6:0] ? phv_data_50 : _GEN_2578; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2580 = 7'h33 == total_offset_48[6:0] ? phv_data_51 : _GEN_2579; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2581 = 7'h34 == total_offset_48[6:0] ? phv_data_52 : _GEN_2580; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2582 = 7'h35 == total_offset_48[6:0] ? phv_data_53 : _GEN_2581; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2583 = 7'h36 == total_offset_48[6:0] ? phv_data_54 : _GEN_2582; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2584 = 7'h37 == total_offset_48[6:0] ? phv_data_55 : _GEN_2583; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2585 = 7'h38 == total_offset_48[6:0] ? phv_data_56 : _GEN_2584; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2586 = 7'h39 == total_offset_48[6:0] ? phv_data_57 : _GEN_2585; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2587 = 7'h3a == total_offset_48[6:0] ? phv_data_58 : _GEN_2586; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2588 = 7'h3b == total_offset_48[6:0] ? phv_data_59 : _GEN_2587; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2589 = 7'h3c == total_offset_48[6:0] ? phv_data_60 : _GEN_2588; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2590 = 7'h3d == total_offset_48[6:0] ? phv_data_61 : _GEN_2589; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2591 = 7'h3e == total_offset_48[6:0] ? phv_data_62 : _GEN_2590; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2592 = 7'h3f == total_offset_48[6:0] ? phv_data_63 : _GEN_2591; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2593 = 7'h40 == total_offset_48[6:0] ? phv_data_64 : _GEN_2592; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2594 = 7'h41 == total_offset_48[6:0] ? phv_data_65 : _GEN_2593; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2595 = 7'h42 == total_offset_48[6:0] ? phv_data_66 : _GEN_2594; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2596 = 7'h43 == total_offset_48[6:0] ? phv_data_67 : _GEN_2595; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2597 = 7'h44 == total_offset_48[6:0] ? phv_data_68 : _GEN_2596; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2598 = 7'h45 == total_offset_48[6:0] ? phv_data_69 : _GEN_2597; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2599 = 7'h46 == total_offset_48[6:0] ? phv_data_70 : _GEN_2598; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2600 = 7'h47 == total_offset_48[6:0] ? phv_data_71 : _GEN_2599; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2601 = 7'h48 == total_offset_48[6:0] ? phv_data_72 : _GEN_2600; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2602 = 7'h49 == total_offset_48[6:0] ? phv_data_73 : _GEN_2601; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2603 = 7'h4a == total_offset_48[6:0] ? phv_data_74 : _GEN_2602; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2604 = 7'h4b == total_offset_48[6:0] ? phv_data_75 : _GEN_2603; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2605 = 7'h4c == total_offset_48[6:0] ? phv_data_76 : _GEN_2604; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2606 = 7'h4d == total_offset_48[6:0] ? phv_data_77 : _GEN_2605; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2607 = 7'h4e == total_offset_48[6:0] ? phv_data_78 : _GEN_2606; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2608 = 7'h4f == total_offset_48[6:0] ? phv_data_79 : _GEN_2607; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2609 = 7'h50 == total_offset_48[6:0] ? phv_data_80 : _GEN_2608; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2610 = 7'h51 == total_offset_48[6:0] ? phv_data_81 : _GEN_2609; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2611 = 7'h52 == total_offset_48[6:0] ? phv_data_82 : _GEN_2610; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2612 = 7'h53 == total_offset_48[6:0] ? phv_data_83 : _GEN_2611; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2613 = 7'h54 == total_offset_48[6:0] ? phv_data_84 : _GEN_2612; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2614 = 7'h55 == total_offset_48[6:0] ? phv_data_85 : _GEN_2613; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2615 = 7'h56 == total_offset_48[6:0] ? phv_data_86 : _GEN_2614; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2616 = 7'h57 == total_offset_48[6:0] ? phv_data_87 : _GEN_2615; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2617 = 7'h58 == total_offset_48[6:0] ? phv_data_88 : _GEN_2616; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2618 = 7'h59 == total_offset_48[6:0] ? phv_data_89 : _GEN_2617; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2619 = 7'h5a == total_offset_48[6:0] ? phv_data_90 : _GEN_2618; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2620 = 7'h5b == total_offset_48[6:0] ? phv_data_91 : _GEN_2619; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2621 = 7'h5c == total_offset_48[6:0] ? phv_data_92 : _GEN_2620; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2622 = 7'h5d == total_offset_48[6:0] ? phv_data_93 : _GEN_2621; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2623 = 7'h5e == total_offset_48[6:0] ? phv_data_94 : _GEN_2622; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2624 = 7'h5f == total_offset_48[6:0] ? phv_data_95 : _GEN_2623; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes_6_0 = 8'h0 < length_3 ? _GEN_2624 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_49 = offset_3 + 8'h1; // @[executor.scala 158:57]
  wire [7:0] _GEN_2627 = 7'h1 == total_offset_49[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2628 = 7'h2 == total_offset_49[6:0] ? phv_data_2 : _GEN_2627; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2629 = 7'h3 == total_offset_49[6:0] ? phv_data_3 : _GEN_2628; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2630 = 7'h4 == total_offset_49[6:0] ? phv_data_4 : _GEN_2629; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2631 = 7'h5 == total_offset_49[6:0] ? phv_data_5 : _GEN_2630; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2632 = 7'h6 == total_offset_49[6:0] ? phv_data_6 : _GEN_2631; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2633 = 7'h7 == total_offset_49[6:0] ? phv_data_7 : _GEN_2632; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2634 = 7'h8 == total_offset_49[6:0] ? phv_data_8 : _GEN_2633; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2635 = 7'h9 == total_offset_49[6:0] ? phv_data_9 : _GEN_2634; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2636 = 7'ha == total_offset_49[6:0] ? phv_data_10 : _GEN_2635; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2637 = 7'hb == total_offset_49[6:0] ? phv_data_11 : _GEN_2636; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2638 = 7'hc == total_offset_49[6:0] ? phv_data_12 : _GEN_2637; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2639 = 7'hd == total_offset_49[6:0] ? phv_data_13 : _GEN_2638; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2640 = 7'he == total_offset_49[6:0] ? phv_data_14 : _GEN_2639; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2641 = 7'hf == total_offset_49[6:0] ? phv_data_15 : _GEN_2640; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2642 = 7'h10 == total_offset_49[6:0] ? phv_data_16 : _GEN_2641; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2643 = 7'h11 == total_offset_49[6:0] ? phv_data_17 : _GEN_2642; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2644 = 7'h12 == total_offset_49[6:0] ? phv_data_18 : _GEN_2643; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2645 = 7'h13 == total_offset_49[6:0] ? phv_data_19 : _GEN_2644; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2646 = 7'h14 == total_offset_49[6:0] ? phv_data_20 : _GEN_2645; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2647 = 7'h15 == total_offset_49[6:0] ? phv_data_21 : _GEN_2646; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2648 = 7'h16 == total_offset_49[6:0] ? phv_data_22 : _GEN_2647; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2649 = 7'h17 == total_offset_49[6:0] ? phv_data_23 : _GEN_2648; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2650 = 7'h18 == total_offset_49[6:0] ? phv_data_24 : _GEN_2649; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2651 = 7'h19 == total_offset_49[6:0] ? phv_data_25 : _GEN_2650; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2652 = 7'h1a == total_offset_49[6:0] ? phv_data_26 : _GEN_2651; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2653 = 7'h1b == total_offset_49[6:0] ? phv_data_27 : _GEN_2652; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2654 = 7'h1c == total_offset_49[6:0] ? phv_data_28 : _GEN_2653; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2655 = 7'h1d == total_offset_49[6:0] ? phv_data_29 : _GEN_2654; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2656 = 7'h1e == total_offset_49[6:0] ? phv_data_30 : _GEN_2655; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2657 = 7'h1f == total_offset_49[6:0] ? phv_data_31 : _GEN_2656; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2658 = 7'h20 == total_offset_49[6:0] ? phv_data_32 : _GEN_2657; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2659 = 7'h21 == total_offset_49[6:0] ? phv_data_33 : _GEN_2658; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2660 = 7'h22 == total_offset_49[6:0] ? phv_data_34 : _GEN_2659; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2661 = 7'h23 == total_offset_49[6:0] ? phv_data_35 : _GEN_2660; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2662 = 7'h24 == total_offset_49[6:0] ? phv_data_36 : _GEN_2661; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2663 = 7'h25 == total_offset_49[6:0] ? phv_data_37 : _GEN_2662; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2664 = 7'h26 == total_offset_49[6:0] ? phv_data_38 : _GEN_2663; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2665 = 7'h27 == total_offset_49[6:0] ? phv_data_39 : _GEN_2664; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2666 = 7'h28 == total_offset_49[6:0] ? phv_data_40 : _GEN_2665; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2667 = 7'h29 == total_offset_49[6:0] ? phv_data_41 : _GEN_2666; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2668 = 7'h2a == total_offset_49[6:0] ? phv_data_42 : _GEN_2667; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2669 = 7'h2b == total_offset_49[6:0] ? phv_data_43 : _GEN_2668; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2670 = 7'h2c == total_offset_49[6:0] ? phv_data_44 : _GEN_2669; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2671 = 7'h2d == total_offset_49[6:0] ? phv_data_45 : _GEN_2670; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2672 = 7'h2e == total_offset_49[6:0] ? phv_data_46 : _GEN_2671; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2673 = 7'h2f == total_offset_49[6:0] ? phv_data_47 : _GEN_2672; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2674 = 7'h30 == total_offset_49[6:0] ? phv_data_48 : _GEN_2673; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2675 = 7'h31 == total_offset_49[6:0] ? phv_data_49 : _GEN_2674; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2676 = 7'h32 == total_offset_49[6:0] ? phv_data_50 : _GEN_2675; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2677 = 7'h33 == total_offset_49[6:0] ? phv_data_51 : _GEN_2676; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2678 = 7'h34 == total_offset_49[6:0] ? phv_data_52 : _GEN_2677; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2679 = 7'h35 == total_offset_49[6:0] ? phv_data_53 : _GEN_2678; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2680 = 7'h36 == total_offset_49[6:0] ? phv_data_54 : _GEN_2679; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2681 = 7'h37 == total_offset_49[6:0] ? phv_data_55 : _GEN_2680; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2682 = 7'h38 == total_offset_49[6:0] ? phv_data_56 : _GEN_2681; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2683 = 7'h39 == total_offset_49[6:0] ? phv_data_57 : _GEN_2682; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2684 = 7'h3a == total_offset_49[6:0] ? phv_data_58 : _GEN_2683; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2685 = 7'h3b == total_offset_49[6:0] ? phv_data_59 : _GEN_2684; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2686 = 7'h3c == total_offset_49[6:0] ? phv_data_60 : _GEN_2685; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2687 = 7'h3d == total_offset_49[6:0] ? phv_data_61 : _GEN_2686; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2688 = 7'h3e == total_offset_49[6:0] ? phv_data_62 : _GEN_2687; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2689 = 7'h3f == total_offset_49[6:0] ? phv_data_63 : _GEN_2688; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2690 = 7'h40 == total_offset_49[6:0] ? phv_data_64 : _GEN_2689; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2691 = 7'h41 == total_offset_49[6:0] ? phv_data_65 : _GEN_2690; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2692 = 7'h42 == total_offset_49[6:0] ? phv_data_66 : _GEN_2691; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2693 = 7'h43 == total_offset_49[6:0] ? phv_data_67 : _GEN_2692; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2694 = 7'h44 == total_offset_49[6:0] ? phv_data_68 : _GEN_2693; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2695 = 7'h45 == total_offset_49[6:0] ? phv_data_69 : _GEN_2694; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2696 = 7'h46 == total_offset_49[6:0] ? phv_data_70 : _GEN_2695; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2697 = 7'h47 == total_offset_49[6:0] ? phv_data_71 : _GEN_2696; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2698 = 7'h48 == total_offset_49[6:0] ? phv_data_72 : _GEN_2697; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2699 = 7'h49 == total_offset_49[6:0] ? phv_data_73 : _GEN_2698; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2700 = 7'h4a == total_offset_49[6:0] ? phv_data_74 : _GEN_2699; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2701 = 7'h4b == total_offset_49[6:0] ? phv_data_75 : _GEN_2700; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2702 = 7'h4c == total_offset_49[6:0] ? phv_data_76 : _GEN_2701; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2703 = 7'h4d == total_offset_49[6:0] ? phv_data_77 : _GEN_2702; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2704 = 7'h4e == total_offset_49[6:0] ? phv_data_78 : _GEN_2703; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2705 = 7'h4f == total_offset_49[6:0] ? phv_data_79 : _GEN_2704; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2706 = 7'h50 == total_offset_49[6:0] ? phv_data_80 : _GEN_2705; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2707 = 7'h51 == total_offset_49[6:0] ? phv_data_81 : _GEN_2706; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2708 = 7'h52 == total_offset_49[6:0] ? phv_data_82 : _GEN_2707; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2709 = 7'h53 == total_offset_49[6:0] ? phv_data_83 : _GEN_2708; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2710 = 7'h54 == total_offset_49[6:0] ? phv_data_84 : _GEN_2709; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2711 = 7'h55 == total_offset_49[6:0] ? phv_data_85 : _GEN_2710; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2712 = 7'h56 == total_offset_49[6:0] ? phv_data_86 : _GEN_2711; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2713 = 7'h57 == total_offset_49[6:0] ? phv_data_87 : _GEN_2712; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2714 = 7'h58 == total_offset_49[6:0] ? phv_data_88 : _GEN_2713; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2715 = 7'h59 == total_offset_49[6:0] ? phv_data_89 : _GEN_2714; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2716 = 7'h5a == total_offset_49[6:0] ? phv_data_90 : _GEN_2715; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2717 = 7'h5b == total_offset_49[6:0] ? phv_data_91 : _GEN_2716; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2718 = 7'h5c == total_offset_49[6:0] ? phv_data_92 : _GEN_2717; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2719 = 7'h5d == total_offset_49[6:0] ? phv_data_93 : _GEN_2718; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2720 = 7'h5e == total_offset_49[6:0] ? phv_data_94 : _GEN_2719; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2721 = 7'h5f == total_offset_49[6:0] ? phv_data_95 : _GEN_2720; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes_6_1 = 8'h1 < length_3 ? _GEN_2721 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_50 = offset_3 + 8'h2; // @[executor.scala 158:57]
  wire [7:0] _GEN_2724 = 7'h1 == total_offset_50[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2725 = 7'h2 == total_offset_50[6:0] ? phv_data_2 : _GEN_2724; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2726 = 7'h3 == total_offset_50[6:0] ? phv_data_3 : _GEN_2725; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2727 = 7'h4 == total_offset_50[6:0] ? phv_data_4 : _GEN_2726; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2728 = 7'h5 == total_offset_50[6:0] ? phv_data_5 : _GEN_2727; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2729 = 7'h6 == total_offset_50[6:0] ? phv_data_6 : _GEN_2728; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2730 = 7'h7 == total_offset_50[6:0] ? phv_data_7 : _GEN_2729; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2731 = 7'h8 == total_offset_50[6:0] ? phv_data_8 : _GEN_2730; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2732 = 7'h9 == total_offset_50[6:0] ? phv_data_9 : _GEN_2731; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2733 = 7'ha == total_offset_50[6:0] ? phv_data_10 : _GEN_2732; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2734 = 7'hb == total_offset_50[6:0] ? phv_data_11 : _GEN_2733; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2735 = 7'hc == total_offset_50[6:0] ? phv_data_12 : _GEN_2734; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2736 = 7'hd == total_offset_50[6:0] ? phv_data_13 : _GEN_2735; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2737 = 7'he == total_offset_50[6:0] ? phv_data_14 : _GEN_2736; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2738 = 7'hf == total_offset_50[6:0] ? phv_data_15 : _GEN_2737; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2739 = 7'h10 == total_offset_50[6:0] ? phv_data_16 : _GEN_2738; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2740 = 7'h11 == total_offset_50[6:0] ? phv_data_17 : _GEN_2739; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2741 = 7'h12 == total_offset_50[6:0] ? phv_data_18 : _GEN_2740; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2742 = 7'h13 == total_offset_50[6:0] ? phv_data_19 : _GEN_2741; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2743 = 7'h14 == total_offset_50[6:0] ? phv_data_20 : _GEN_2742; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2744 = 7'h15 == total_offset_50[6:0] ? phv_data_21 : _GEN_2743; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2745 = 7'h16 == total_offset_50[6:0] ? phv_data_22 : _GEN_2744; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2746 = 7'h17 == total_offset_50[6:0] ? phv_data_23 : _GEN_2745; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2747 = 7'h18 == total_offset_50[6:0] ? phv_data_24 : _GEN_2746; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2748 = 7'h19 == total_offset_50[6:0] ? phv_data_25 : _GEN_2747; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2749 = 7'h1a == total_offset_50[6:0] ? phv_data_26 : _GEN_2748; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2750 = 7'h1b == total_offset_50[6:0] ? phv_data_27 : _GEN_2749; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2751 = 7'h1c == total_offset_50[6:0] ? phv_data_28 : _GEN_2750; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2752 = 7'h1d == total_offset_50[6:0] ? phv_data_29 : _GEN_2751; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2753 = 7'h1e == total_offset_50[6:0] ? phv_data_30 : _GEN_2752; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2754 = 7'h1f == total_offset_50[6:0] ? phv_data_31 : _GEN_2753; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2755 = 7'h20 == total_offset_50[6:0] ? phv_data_32 : _GEN_2754; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2756 = 7'h21 == total_offset_50[6:0] ? phv_data_33 : _GEN_2755; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2757 = 7'h22 == total_offset_50[6:0] ? phv_data_34 : _GEN_2756; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2758 = 7'h23 == total_offset_50[6:0] ? phv_data_35 : _GEN_2757; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2759 = 7'h24 == total_offset_50[6:0] ? phv_data_36 : _GEN_2758; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2760 = 7'h25 == total_offset_50[6:0] ? phv_data_37 : _GEN_2759; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2761 = 7'h26 == total_offset_50[6:0] ? phv_data_38 : _GEN_2760; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2762 = 7'h27 == total_offset_50[6:0] ? phv_data_39 : _GEN_2761; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2763 = 7'h28 == total_offset_50[6:0] ? phv_data_40 : _GEN_2762; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2764 = 7'h29 == total_offset_50[6:0] ? phv_data_41 : _GEN_2763; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2765 = 7'h2a == total_offset_50[6:0] ? phv_data_42 : _GEN_2764; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2766 = 7'h2b == total_offset_50[6:0] ? phv_data_43 : _GEN_2765; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2767 = 7'h2c == total_offset_50[6:0] ? phv_data_44 : _GEN_2766; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2768 = 7'h2d == total_offset_50[6:0] ? phv_data_45 : _GEN_2767; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2769 = 7'h2e == total_offset_50[6:0] ? phv_data_46 : _GEN_2768; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2770 = 7'h2f == total_offset_50[6:0] ? phv_data_47 : _GEN_2769; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2771 = 7'h30 == total_offset_50[6:0] ? phv_data_48 : _GEN_2770; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2772 = 7'h31 == total_offset_50[6:0] ? phv_data_49 : _GEN_2771; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2773 = 7'h32 == total_offset_50[6:0] ? phv_data_50 : _GEN_2772; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2774 = 7'h33 == total_offset_50[6:0] ? phv_data_51 : _GEN_2773; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2775 = 7'h34 == total_offset_50[6:0] ? phv_data_52 : _GEN_2774; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2776 = 7'h35 == total_offset_50[6:0] ? phv_data_53 : _GEN_2775; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2777 = 7'h36 == total_offset_50[6:0] ? phv_data_54 : _GEN_2776; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2778 = 7'h37 == total_offset_50[6:0] ? phv_data_55 : _GEN_2777; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2779 = 7'h38 == total_offset_50[6:0] ? phv_data_56 : _GEN_2778; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2780 = 7'h39 == total_offset_50[6:0] ? phv_data_57 : _GEN_2779; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2781 = 7'h3a == total_offset_50[6:0] ? phv_data_58 : _GEN_2780; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2782 = 7'h3b == total_offset_50[6:0] ? phv_data_59 : _GEN_2781; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2783 = 7'h3c == total_offset_50[6:0] ? phv_data_60 : _GEN_2782; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2784 = 7'h3d == total_offset_50[6:0] ? phv_data_61 : _GEN_2783; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2785 = 7'h3e == total_offset_50[6:0] ? phv_data_62 : _GEN_2784; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2786 = 7'h3f == total_offset_50[6:0] ? phv_data_63 : _GEN_2785; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2787 = 7'h40 == total_offset_50[6:0] ? phv_data_64 : _GEN_2786; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2788 = 7'h41 == total_offset_50[6:0] ? phv_data_65 : _GEN_2787; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2789 = 7'h42 == total_offset_50[6:0] ? phv_data_66 : _GEN_2788; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2790 = 7'h43 == total_offset_50[6:0] ? phv_data_67 : _GEN_2789; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2791 = 7'h44 == total_offset_50[6:0] ? phv_data_68 : _GEN_2790; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2792 = 7'h45 == total_offset_50[6:0] ? phv_data_69 : _GEN_2791; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2793 = 7'h46 == total_offset_50[6:0] ? phv_data_70 : _GEN_2792; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2794 = 7'h47 == total_offset_50[6:0] ? phv_data_71 : _GEN_2793; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2795 = 7'h48 == total_offset_50[6:0] ? phv_data_72 : _GEN_2794; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2796 = 7'h49 == total_offset_50[6:0] ? phv_data_73 : _GEN_2795; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2797 = 7'h4a == total_offset_50[6:0] ? phv_data_74 : _GEN_2796; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2798 = 7'h4b == total_offset_50[6:0] ? phv_data_75 : _GEN_2797; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2799 = 7'h4c == total_offset_50[6:0] ? phv_data_76 : _GEN_2798; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2800 = 7'h4d == total_offset_50[6:0] ? phv_data_77 : _GEN_2799; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2801 = 7'h4e == total_offset_50[6:0] ? phv_data_78 : _GEN_2800; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2802 = 7'h4f == total_offset_50[6:0] ? phv_data_79 : _GEN_2801; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2803 = 7'h50 == total_offset_50[6:0] ? phv_data_80 : _GEN_2802; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2804 = 7'h51 == total_offset_50[6:0] ? phv_data_81 : _GEN_2803; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2805 = 7'h52 == total_offset_50[6:0] ? phv_data_82 : _GEN_2804; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2806 = 7'h53 == total_offset_50[6:0] ? phv_data_83 : _GEN_2805; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2807 = 7'h54 == total_offset_50[6:0] ? phv_data_84 : _GEN_2806; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2808 = 7'h55 == total_offset_50[6:0] ? phv_data_85 : _GEN_2807; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2809 = 7'h56 == total_offset_50[6:0] ? phv_data_86 : _GEN_2808; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2810 = 7'h57 == total_offset_50[6:0] ? phv_data_87 : _GEN_2809; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2811 = 7'h58 == total_offset_50[6:0] ? phv_data_88 : _GEN_2810; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2812 = 7'h59 == total_offset_50[6:0] ? phv_data_89 : _GEN_2811; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2813 = 7'h5a == total_offset_50[6:0] ? phv_data_90 : _GEN_2812; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2814 = 7'h5b == total_offset_50[6:0] ? phv_data_91 : _GEN_2813; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2815 = 7'h5c == total_offset_50[6:0] ? phv_data_92 : _GEN_2814; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2816 = 7'h5d == total_offset_50[6:0] ? phv_data_93 : _GEN_2815; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2817 = 7'h5e == total_offset_50[6:0] ? phv_data_94 : _GEN_2816; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2818 = 7'h5f == total_offset_50[6:0] ? phv_data_95 : _GEN_2817; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes_6_2 = 8'h2 < length_3 ? _GEN_2818 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_51 = offset_3 + 8'h3; // @[executor.scala 158:57]
  wire [7:0] _GEN_2821 = 7'h1 == total_offset_51[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2822 = 7'h2 == total_offset_51[6:0] ? phv_data_2 : _GEN_2821; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2823 = 7'h3 == total_offset_51[6:0] ? phv_data_3 : _GEN_2822; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2824 = 7'h4 == total_offset_51[6:0] ? phv_data_4 : _GEN_2823; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2825 = 7'h5 == total_offset_51[6:0] ? phv_data_5 : _GEN_2824; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2826 = 7'h6 == total_offset_51[6:0] ? phv_data_6 : _GEN_2825; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2827 = 7'h7 == total_offset_51[6:0] ? phv_data_7 : _GEN_2826; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2828 = 7'h8 == total_offset_51[6:0] ? phv_data_8 : _GEN_2827; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2829 = 7'h9 == total_offset_51[6:0] ? phv_data_9 : _GEN_2828; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2830 = 7'ha == total_offset_51[6:0] ? phv_data_10 : _GEN_2829; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2831 = 7'hb == total_offset_51[6:0] ? phv_data_11 : _GEN_2830; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2832 = 7'hc == total_offset_51[6:0] ? phv_data_12 : _GEN_2831; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2833 = 7'hd == total_offset_51[6:0] ? phv_data_13 : _GEN_2832; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2834 = 7'he == total_offset_51[6:0] ? phv_data_14 : _GEN_2833; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2835 = 7'hf == total_offset_51[6:0] ? phv_data_15 : _GEN_2834; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2836 = 7'h10 == total_offset_51[6:0] ? phv_data_16 : _GEN_2835; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2837 = 7'h11 == total_offset_51[6:0] ? phv_data_17 : _GEN_2836; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2838 = 7'h12 == total_offset_51[6:0] ? phv_data_18 : _GEN_2837; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2839 = 7'h13 == total_offset_51[6:0] ? phv_data_19 : _GEN_2838; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2840 = 7'h14 == total_offset_51[6:0] ? phv_data_20 : _GEN_2839; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2841 = 7'h15 == total_offset_51[6:0] ? phv_data_21 : _GEN_2840; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2842 = 7'h16 == total_offset_51[6:0] ? phv_data_22 : _GEN_2841; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2843 = 7'h17 == total_offset_51[6:0] ? phv_data_23 : _GEN_2842; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2844 = 7'h18 == total_offset_51[6:0] ? phv_data_24 : _GEN_2843; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2845 = 7'h19 == total_offset_51[6:0] ? phv_data_25 : _GEN_2844; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2846 = 7'h1a == total_offset_51[6:0] ? phv_data_26 : _GEN_2845; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2847 = 7'h1b == total_offset_51[6:0] ? phv_data_27 : _GEN_2846; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2848 = 7'h1c == total_offset_51[6:0] ? phv_data_28 : _GEN_2847; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2849 = 7'h1d == total_offset_51[6:0] ? phv_data_29 : _GEN_2848; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2850 = 7'h1e == total_offset_51[6:0] ? phv_data_30 : _GEN_2849; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2851 = 7'h1f == total_offset_51[6:0] ? phv_data_31 : _GEN_2850; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2852 = 7'h20 == total_offset_51[6:0] ? phv_data_32 : _GEN_2851; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2853 = 7'h21 == total_offset_51[6:0] ? phv_data_33 : _GEN_2852; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2854 = 7'h22 == total_offset_51[6:0] ? phv_data_34 : _GEN_2853; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2855 = 7'h23 == total_offset_51[6:0] ? phv_data_35 : _GEN_2854; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2856 = 7'h24 == total_offset_51[6:0] ? phv_data_36 : _GEN_2855; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2857 = 7'h25 == total_offset_51[6:0] ? phv_data_37 : _GEN_2856; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2858 = 7'h26 == total_offset_51[6:0] ? phv_data_38 : _GEN_2857; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2859 = 7'h27 == total_offset_51[6:0] ? phv_data_39 : _GEN_2858; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2860 = 7'h28 == total_offset_51[6:0] ? phv_data_40 : _GEN_2859; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2861 = 7'h29 == total_offset_51[6:0] ? phv_data_41 : _GEN_2860; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2862 = 7'h2a == total_offset_51[6:0] ? phv_data_42 : _GEN_2861; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2863 = 7'h2b == total_offset_51[6:0] ? phv_data_43 : _GEN_2862; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2864 = 7'h2c == total_offset_51[6:0] ? phv_data_44 : _GEN_2863; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2865 = 7'h2d == total_offset_51[6:0] ? phv_data_45 : _GEN_2864; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2866 = 7'h2e == total_offset_51[6:0] ? phv_data_46 : _GEN_2865; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2867 = 7'h2f == total_offset_51[6:0] ? phv_data_47 : _GEN_2866; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2868 = 7'h30 == total_offset_51[6:0] ? phv_data_48 : _GEN_2867; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2869 = 7'h31 == total_offset_51[6:0] ? phv_data_49 : _GEN_2868; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2870 = 7'h32 == total_offset_51[6:0] ? phv_data_50 : _GEN_2869; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2871 = 7'h33 == total_offset_51[6:0] ? phv_data_51 : _GEN_2870; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2872 = 7'h34 == total_offset_51[6:0] ? phv_data_52 : _GEN_2871; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2873 = 7'h35 == total_offset_51[6:0] ? phv_data_53 : _GEN_2872; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2874 = 7'h36 == total_offset_51[6:0] ? phv_data_54 : _GEN_2873; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2875 = 7'h37 == total_offset_51[6:0] ? phv_data_55 : _GEN_2874; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2876 = 7'h38 == total_offset_51[6:0] ? phv_data_56 : _GEN_2875; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2877 = 7'h39 == total_offset_51[6:0] ? phv_data_57 : _GEN_2876; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2878 = 7'h3a == total_offset_51[6:0] ? phv_data_58 : _GEN_2877; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2879 = 7'h3b == total_offset_51[6:0] ? phv_data_59 : _GEN_2878; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2880 = 7'h3c == total_offset_51[6:0] ? phv_data_60 : _GEN_2879; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2881 = 7'h3d == total_offset_51[6:0] ? phv_data_61 : _GEN_2880; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2882 = 7'h3e == total_offset_51[6:0] ? phv_data_62 : _GEN_2881; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2883 = 7'h3f == total_offset_51[6:0] ? phv_data_63 : _GEN_2882; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2884 = 7'h40 == total_offset_51[6:0] ? phv_data_64 : _GEN_2883; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2885 = 7'h41 == total_offset_51[6:0] ? phv_data_65 : _GEN_2884; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2886 = 7'h42 == total_offset_51[6:0] ? phv_data_66 : _GEN_2885; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2887 = 7'h43 == total_offset_51[6:0] ? phv_data_67 : _GEN_2886; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2888 = 7'h44 == total_offset_51[6:0] ? phv_data_68 : _GEN_2887; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2889 = 7'h45 == total_offset_51[6:0] ? phv_data_69 : _GEN_2888; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2890 = 7'h46 == total_offset_51[6:0] ? phv_data_70 : _GEN_2889; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2891 = 7'h47 == total_offset_51[6:0] ? phv_data_71 : _GEN_2890; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2892 = 7'h48 == total_offset_51[6:0] ? phv_data_72 : _GEN_2891; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2893 = 7'h49 == total_offset_51[6:0] ? phv_data_73 : _GEN_2892; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2894 = 7'h4a == total_offset_51[6:0] ? phv_data_74 : _GEN_2893; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2895 = 7'h4b == total_offset_51[6:0] ? phv_data_75 : _GEN_2894; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2896 = 7'h4c == total_offset_51[6:0] ? phv_data_76 : _GEN_2895; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2897 = 7'h4d == total_offset_51[6:0] ? phv_data_77 : _GEN_2896; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2898 = 7'h4e == total_offset_51[6:0] ? phv_data_78 : _GEN_2897; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2899 = 7'h4f == total_offset_51[6:0] ? phv_data_79 : _GEN_2898; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2900 = 7'h50 == total_offset_51[6:0] ? phv_data_80 : _GEN_2899; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2901 = 7'h51 == total_offset_51[6:0] ? phv_data_81 : _GEN_2900; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2902 = 7'h52 == total_offset_51[6:0] ? phv_data_82 : _GEN_2901; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2903 = 7'h53 == total_offset_51[6:0] ? phv_data_83 : _GEN_2902; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2904 = 7'h54 == total_offset_51[6:0] ? phv_data_84 : _GEN_2903; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2905 = 7'h55 == total_offset_51[6:0] ? phv_data_85 : _GEN_2904; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2906 = 7'h56 == total_offset_51[6:0] ? phv_data_86 : _GEN_2905; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2907 = 7'h57 == total_offset_51[6:0] ? phv_data_87 : _GEN_2906; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2908 = 7'h58 == total_offset_51[6:0] ? phv_data_88 : _GEN_2907; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2909 = 7'h59 == total_offset_51[6:0] ? phv_data_89 : _GEN_2908; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2910 = 7'h5a == total_offset_51[6:0] ? phv_data_90 : _GEN_2909; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2911 = 7'h5b == total_offset_51[6:0] ? phv_data_91 : _GEN_2910; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2912 = 7'h5c == total_offset_51[6:0] ? phv_data_92 : _GEN_2911; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2913 = 7'h5d == total_offset_51[6:0] ? phv_data_93 : _GEN_2912; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2914 = 7'h5e == total_offset_51[6:0] ? phv_data_94 : _GEN_2913; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2915 = 7'h5f == total_offset_51[6:0] ? phv_data_95 : _GEN_2914; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes_6_3 = 8'h3 < length_3 ? _GEN_2915 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_52 = offset_3 + 8'h4; // @[executor.scala 158:57]
  wire [7:0] _GEN_2918 = 7'h1 == total_offset_52[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2919 = 7'h2 == total_offset_52[6:0] ? phv_data_2 : _GEN_2918; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2920 = 7'h3 == total_offset_52[6:0] ? phv_data_3 : _GEN_2919; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2921 = 7'h4 == total_offset_52[6:0] ? phv_data_4 : _GEN_2920; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2922 = 7'h5 == total_offset_52[6:0] ? phv_data_5 : _GEN_2921; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2923 = 7'h6 == total_offset_52[6:0] ? phv_data_6 : _GEN_2922; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2924 = 7'h7 == total_offset_52[6:0] ? phv_data_7 : _GEN_2923; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2925 = 7'h8 == total_offset_52[6:0] ? phv_data_8 : _GEN_2924; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2926 = 7'h9 == total_offset_52[6:0] ? phv_data_9 : _GEN_2925; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2927 = 7'ha == total_offset_52[6:0] ? phv_data_10 : _GEN_2926; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2928 = 7'hb == total_offset_52[6:0] ? phv_data_11 : _GEN_2927; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2929 = 7'hc == total_offset_52[6:0] ? phv_data_12 : _GEN_2928; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2930 = 7'hd == total_offset_52[6:0] ? phv_data_13 : _GEN_2929; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2931 = 7'he == total_offset_52[6:0] ? phv_data_14 : _GEN_2930; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2932 = 7'hf == total_offset_52[6:0] ? phv_data_15 : _GEN_2931; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2933 = 7'h10 == total_offset_52[6:0] ? phv_data_16 : _GEN_2932; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2934 = 7'h11 == total_offset_52[6:0] ? phv_data_17 : _GEN_2933; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2935 = 7'h12 == total_offset_52[6:0] ? phv_data_18 : _GEN_2934; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2936 = 7'h13 == total_offset_52[6:0] ? phv_data_19 : _GEN_2935; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2937 = 7'h14 == total_offset_52[6:0] ? phv_data_20 : _GEN_2936; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2938 = 7'h15 == total_offset_52[6:0] ? phv_data_21 : _GEN_2937; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2939 = 7'h16 == total_offset_52[6:0] ? phv_data_22 : _GEN_2938; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2940 = 7'h17 == total_offset_52[6:0] ? phv_data_23 : _GEN_2939; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2941 = 7'h18 == total_offset_52[6:0] ? phv_data_24 : _GEN_2940; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2942 = 7'h19 == total_offset_52[6:0] ? phv_data_25 : _GEN_2941; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2943 = 7'h1a == total_offset_52[6:0] ? phv_data_26 : _GEN_2942; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2944 = 7'h1b == total_offset_52[6:0] ? phv_data_27 : _GEN_2943; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2945 = 7'h1c == total_offset_52[6:0] ? phv_data_28 : _GEN_2944; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2946 = 7'h1d == total_offset_52[6:0] ? phv_data_29 : _GEN_2945; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2947 = 7'h1e == total_offset_52[6:0] ? phv_data_30 : _GEN_2946; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2948 = 7'h1f == total_offset_52[6:0] ? phv_data_31 : _GEN_2947; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2949 = 7'h20 == total_offset_52[6:0] ? phv_data_32 : _GEN_2948; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2950 = 7'h21 == total_offset_52[6:0] ? phv_data_33 : _GEN_2949; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2951 = 7'h22 == total_offset_52[6:0] ? phv_data_34 : _GEN_2950; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2952 = 7'h23 == total_offset_52[6:0] ? phv_data_35 : _GEN_2951; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2953 = 7'h24 == total_offset_52[6:0] ? phv_data_36 : _GEN_2952; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2954 = 7'h25 == total_offset_52[6:0] ? phv_data_37 : _GEN_2953; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2955 = 7'h26 == total_offset_52[6:0] ? phv_data_38 : _GEN_2954; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2956 = 7'h27 == total_offset_52[6:0] ? phv_data_39 : _GEN_2955; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2957 = 7'h28 == total_offset_52[6:0] ? phv_data_40 : _GEN_2956; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2958 = 7'h29 == total_offset_52[6:0] ? phv_data_41 : _GEN_2957; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2959 = 7'h2a == total_offset_52[6:0] ? phv_data_42 : _GEN_2958; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2960 = 7'h2b == total_offset_52[6:0] ? phv_data_43 : _GEN_2959; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2961 = 7'h2c == total_offset_52[6:0] ? phv_data_44 : _GEN_2960; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2962 = 7'h2d == total_offset_52[6:0] ? phv_data_45 : _GEN_2961; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2963 = 7'h2e == total_offset_52[6:0] ? phv_data_46 : _GEN_2962; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2964 = 7'h2f == total_offset_52[6:0] ? phv_data_47 : _GEN_2963; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2965 = 7'h30 == total_offset_52[6:0] ? phv_data_48 : _GEN_2964; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2966 = 7'h31 == total_offset_52[6:0] ? phv_data_49 : _GEN_2965; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2967 = 7'h32 == total_offset_52[6:0] ? phv_data_50 : _GEN_2966; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2968 = 7'h33 == total_offset_52[6:0] ? phv_data_51 : _GEN_2967; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2969 = 7'h34 == total_offset_52[6:0] ? phv_data_52 : _GEN_2968; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2970 = 7'h35 == total_offset_52[6:0] ? phv_data_53 : _GEN_2969; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2971 = 7'h36 == total_offset_52[6:0] ? phv_data_54 : _GEN_2970; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2972 = 7'h37 == total_offset_52[6:0] ? phv_data_55 : _GEN_2971; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2973 = 7'h38 == total_offset_52[6:0] ? phv_data_56 : _GEN_2972; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2974 = 7'h39 == total_offset_52[6:0] ? phv_data_57 : _GEN_2973; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2975 = 7'h3a == total_offset_52[6:0] ? phv_data_58 : _GEN_2974; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2976 = 7'h3b == total_offset_52[6:0] ? phv_data_59 : _GEN_2975; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2977 = 7'h3c == total_offset_52[6:0] ? phv_data_60 : _GEN_2976; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2978 = 7'h3d == total_offset_52[6:0] ? phv_data_61 : _GEN_2977; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2979 = 7'h3e == total_offset_52[6:0] ? phv_data_62 : _GEN_2978; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2980 = 7'h3f == total_offset_52[6:0] ? phv_data_63 : _GEN_2979; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2981 = 7'h40 == total_offset_52[6:0] ? phv_data_64 : _GEN_2980; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2982 = 7'h41 == total_offset_52[6:0] ? phv_data_65 : _GEN_2981; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2983 = 7'h42 == total_offset_52[6:0] ? phv_data_66 : _GEN_2982; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2984 = 7'h43 == total_offset_52[6:0] ? phv_data_67 : _GEN_2983; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2985 = 7'h44 == total_offset_52[6:0] ? phv_data_68 : _GEN_2984; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2986 = 7'h45 == total_offset_52[6:0] ? phv_data_69 : _GEN_2985; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2987 = 7'h46 == total_offset_52[6:0] ? phv_data_70 : _GEN_2986; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2988 = 7'h47 == total_offset_52[6:0] ? phv_data_71 : _GEN_2987; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2989 = 7'h48 == total_offset_52[6:0] ? phv_data_72 : _GEN_2988; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2990 = 7'h49 == total_offset_52[6:0] ? phv_data_73 : _GEN_2989; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2991 = 7'h4a == total_offset_52[6:0] ? phv_data_74 : _GEN_2990; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2992 = 7'h4b == total_offset_52[6:0] ? phv_data_75 : _GEN_2991; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2993 = 7'h4c == total_offset_52[6:0] ? phv_data_76 : _GEN_2992; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2994 = 7'h4d == total_offset_52[6:0] ? phv_data_77 : _GEN_2993; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2995 = 7'h4e == total_offset_52[6:0] ? phv_data_78 : _GEN_2994; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2996 = 7'h4f == total_offset_52[6:0] ? phv_data_79 : _GEN_2995; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2997 = 7'h50 == total_offset_52[6:0] ? phv_data_80 : _GEN_2996; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2998 = 7'h51 == total_offset_52[6:0] ? phv_data_81 : _GEN_2997; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_2999 = 7'h52 == total_offset_52[6:0] ? phv_data_82 : _GEN_2998; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3000 = 7'h53 == total_offset_52[6:0] ? phv_data_83 : _GEN_2999; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3001 = 7'h54 == total_offset_52[6:0] ? phv_data_84 : _GEN_3000; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3002 = 7'h55 == total_offset_52[6:0] ? phv_data_85 : _GEN_3001; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3003 = 7'h56 == total_offset_52[6:0] ? phv_data_86 : _GEN_3002; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3004 = 7'h57 == total_offset_52[6:0] ? phv_data_87 : _GEN_3003; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3005 = 7'h58 == total_offset_52[6:0] ? phv_data_88 : _GEN_3004; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3006 = 7'h59 == total_offset_52[6:0] ? phv_data_89 : _GEN_3005; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3007 = 7'h5a == total_offset_52[6:0] ? phv_data_90 : _GEN_3006; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3008 = 7'h5b == total_offset_52[6:0] ? phv_data_91 : _GEN_3007; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3009 = 7'h5c == total_offset_52[6:0] ? phv_data_92 : _GEN_3008; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3010 = 7'h5d == total_offset_52[6:0] ? phv_data_93 : _GEN_3009; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3011 = 7'h5e == total_offset_52[6:0] ? phv_data_94 : _GEN_3010; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3012 = 7'h5f == total_offset_52[6:0] ? phv_data_95 : _GEN_3011; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes_6_4 = 8'h4 < length_3 ? _GEN_3012 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_53 = offset_3 + 8'h5; // @[executor.scala 158:57]
  wire [7:0] _GEN_3015 = 7'h1 == total_offset_53[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3016 = 7'h2 == total_offset_53[6:0] ? phv_data_2 : _GEN_3015; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3017 = 7'h3 == total_offset_53[6:0] ? phv_data_3 : _GEN_3016; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3018 = 7'h4 == total_offset_53[6:0] ? phv_data_4 : _GEN_3017; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3019 = 7'h5 == total_offset_53[6:0] ? phv_data_5 : _GEN_3018; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3020 = 7'h6 == total_offset_53[6:0] ? phv_data_6 : _GEN_3019; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3021 = 7'h7 == total_offset_53[6:0] ? phv_data_7 : _GEN_3020; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3022 = 7'h8 == total_offset_53[6:0] ? phv_data_8 : _GEN_3021; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3023 = 7'h9 == total_offset_53[6:0] ? phv_data_9 : _GEN_3022; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3024 = 7'ha == total_offset_53[6:0] ? phv_data_10 : _GEN_3023; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3025 = 7'hb == total_offset_53[6:0] ? phv_data_11 : _GEN_3024; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3026 = 7'hc == total_offset_53[6:0] ? phv_data_12 : _GEN_3025; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3027 = 7'hd == total_offset_53[6:0] ? phv_data_13 : _GEN_3026; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3028 = 7'he == total_offset_53[6:0] ? phv_data_14 : _GEN_3027; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3029 = 7'hf == total_offset_53[6:0] ? phv_data_15 : _GEN_3028; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3030 = 7'h10 == total_offset_53[6:0] ? phv_data_16 : _GEN_3029; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3031 = 7'h11 == total_offset_53[6:0] ? phv_data_17 : _GEN_3030; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3032 = 7'h12 == total_offset_53[6:0] ? phv_data_18 : _GEN_3031; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3033 = 7'h13 == total_offset_53[6:0] ? phv_data_19 : _GEN_3032; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3034 = 7'h14 == total_offset_53[6:0] ? phv_data_20 : _GEN_3033; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3035 = 7'h15 == total_offset_53[6:0] ? phv_data_21 : _GEN_3034; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3036 = 7'h16 == total_offset_53[6:0] ? phv_data_22 : _GEN_3035; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3037 = 7'h17 == total_offset_53[6:0] ? phv_data_23 : _GEN_3036; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3038 = 7'h18 == total_offset_53[6:0] ? phv_data_24 : _GEN_3037; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3039 = 7'h19 == total_offset_53[6:0] ? phv_data_25 : _GEN_3038; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3040 = 7'h1a == total_offset_53[6:0] ? phv_data_26 : _GEN_3039; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3041 = 7'h1b == total_offset_53[6:0] ? phv_data_27 : _GEN_3040; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3042 = 7'h1c == total_offset_53[6:0] ? phv_data_28 : _GEN_3041; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3043 = 7'h1d == total_offset_53[6:0] ? phv_data_29 : _GEN_3042; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3044 = 7'h1e == total_offset_53[6:0] ? phv_data_30 : _GEN_3043; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3045 = 7'h1f == total_offset_53[6:0] ? phv_data_31 : _GEN_3044; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3046 = 7'h20 == total_offset_53[6:0] ? phv_data_32 : _GEN_3045; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3047 = 7'h21 == total_offset_53[6:0] ? phv_data_33 : _GEN_3046; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3048 = 7'h22 == total_offset_53[6:0] ? phv_data_34 : _GEN_3047; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3049 = 7'h23 == total_offset_53[6:0] ? phv_data_35 : _GEN_3048; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3050 = 7'h24 == total_offset_53[6:0] ? phv_data_36 : _GEN_3049; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3051 = 7'h25 == total_offset_53[6:0] ? phv_data_37 : _GEN_3050; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3052 = 7'h26 == total_offset_53[6:0] ? phv_data_38 : _GEN_3051; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3053 = 7'h27 == total_offset_53[6:0] ? phv_data_39 : _GEN_3052; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3054 = 7'h28 == total_offset_53[6:0] ? phv_data_40 : _GEN_3053; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3055 = 7'h29 == total_offset_53[6:0] ? phv_data_41 : _GEN_3054; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3056 = 7'h2a == total_offset_53[6:0] ? phv_data_42 : _GEN_3055; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3057 = 7'h2b == total_offset_53[6:0] ? phv_data_43 : _GEN_3056; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3058 = 7'h2c == total_offset_53[6:0] ? phv_data_44 : _GEN_3057; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3059 = 7'h2d == total_offset_53[6:0] ? phv_data_45 : _GEN_3058; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3060 = 7'h2e == total_offset_53[6:0] ? phv_data_46 : _GEN_3059; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3061 = 7'h2f == total_offset_53[6:0] ? phv_data_47 : _GEN_3060; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3062 = 7'h30 == total_offset_53[6:0] ? phv_data_48 : _GEN_3061; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3063 = 7'h31 == total_offset_53[6:0] ? phv_data_49 : _GEN_3062; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3064 = 7'h32 == total_offset_53[6:0] ? phv_data_50 : _GEN_3063; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3065 = 7'h33 == total_offset_53[6:0] ? phv_data_51 : _GEN_3064; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3066 = 7'h34 == total_offset_53[6:0] ? phv_data_52 : _GEN_3065; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3067 = 7'h35 == total_offset_53[6:0] ? phv_data_53 : _GEN_3066; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3068 = 7'h36 == total_offset_53[6:0] ? phv_data_54 : _GEN_3067; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3069 = 7'h37 == total_offset_53[6:0] ? phv_data_55 : _GEN_3068; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3070 = 7'h38 == total_offset_53[6:0] ? phv_data_56 : _GEN_3069; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3071 = 7'h39 == total_offset_53[6:0] ? phv_data_57 : _GEN_3070; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3072 = 7'h3a == total_offset_53[6:0] ? phv_data_58 : _GEN_3071; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3073 = 7'h3b == total_offset_53[6:0] ? phv_data_59 : _GEN_3072; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3074 = 7'h3c == total_offset_53[6:0] ? phv_data_60 : _GEN_3073; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3075 = 7'h3d == total_offset_53[6:0] ? phv_data_61 : _GEN_3074; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3076 = 7'h3e == total_offset_53[6:0] ? phv_data_62 : _GEN_3075; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3077 = 7'h3f == total_offset_53[6:0] ? phv_data_63 : _GEN_3076; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3078 = 7'h40 == total_offset_53[6:0] ? phv_data_64 : _GEN_3077; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3079 = 7'h41 == total_offset_53[6:0] ? phv_data_65 : _GEN_3078; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3080 = 7'h42 == total_offset_53[6:0] ? phv_data_66 : _GEN_3079; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3081 = 7'h43 == total_offset_53[6:0] ? phv_data_67 : _GEN_3080; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3082 = 7'h44 == total_offset_53[6:0] ? phv_data_68 : _GEN_3081; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3083 = 7'h45 == total_offset_53[6:0] ? phv_data_69 : _GEN_3082; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3084 = 7'h46 == total_offset_53[6:0] ? phv_data_70 : _GEN_3083; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3085 = 7'h47 == total_offset_53[6:0] ? phv_data_71 : _GEN_3084; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3086 = 7'h48 == total_offset_53[6:0] ? phv_data_72 : _GEN_3085; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3087 = 7'h49 == total_offset_53[6:0] ? phv_data_73 : _GEN_3086; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3088 = 7'h4a == total_offset_53[6:0] ? phv_data_74 : _GEN_3087; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3089 = 7'h4b == total_offset_53[6:0] ? phv_data_75 : _GEN_3088; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3090 = 7'h4c == total_offset_53[6:0] ? phv_data_76 : _GEN_3089; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3091 = 7'h4d == total_offset_53[6:0] ? phv_data_77 : _GEN_3090; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3092 = 7'h4e == total_offset_53[6:0] ? phv_data_78 : _GEN_3091; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3093 = 7'h4f == total_offset_53[6:0] ? phv_data_79 : _GEN_3092; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3094 = 7'h50 == total_offset_53[6:0] ? phv_data_80 : _GEN_3093; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3095 = 7'h51 == total_offset_53[6:0] ? phv_data_81 : _GEN_3094; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3096 = 7'h52 == total_offset_53[6:0] ? phv_data_82 : _GEN_3095; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3097 = 7'h53 == total_offset_53[6:0] ? phv_data_83 : _GEN_3096; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3098 = 7'h54 == total_offset_53[6:0] ? phv_data_84 : _GEN_3097; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3099 = 7'h55 == total_offset_53[6:0] ? phv_data_85 : _GEN_3098; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3100 = 7'h56 == total_offset_53[6:0] ? phv_data_86 : _GEN_3099; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3101 = 7'h57 == total_offset_53[6:0] ? phv_data_87 : _GEN_3100; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3102 = 7'h58 == total_offset_53[6:0] ? phv_data_88 : _GEN_3101; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3103 = 7'h59 == total_offset_53[6:0] ? phv_data_89 : _GEN_3102; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3104 = 7'h5a == total_offset_53[6:0] ? phv_data_90 : _GEN_3103; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3105 = 7'h5b == total_offset_53[6:0] ? phv_data_91 : _GEN_3104; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3106 = 7'h5c == total_offset_53[6:0] ? phv_data_92 : _GEN_3105; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3107 = 7'h5d == total_offset_53[6:0] ? phv_data_93 : _GEN_3106; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3108 = 7'h5e == total_offset_53[6:0] ? phv_data_94 : _GEN_3107; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3109 = 7'h5f == total_offset_53[6:0] ? phv_data_95 : _GEN_3108; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes_6_5 = 8'h5 < length_3 ? _GEN_3109 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_54 = offset_3 + 8'h6; // @[executor.scala 158:57]
  wire [7:0] _GEN_3112 = 7'h1 == total_offset_54[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3113 = 7'h2 == total_offset_54[6:0] ? phv_data_2 : _GEN_3112; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3114 = 7'h3 == total_offset_54[6:0] ? phv_data_3 : _GEN_3113; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3115 = 7'h4 == total_offset_54[6:0] ? phv_data_4 : _GEN_3114; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3116 = 7'h5 == total_offset_54[6:0] ? phv_data_5 : _GEN_3115; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3117 = 7'h6 == total_offset_54[6:0] ? phv_data_6 : _GEN_3116; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3118 = 7'h7 == total_offset_54[6:0] ? phv_data_7 : _GEN_3117; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3119 = 7'h8 == total_offset_54[6:0] ? phv_data_8 : _GEN_3118; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3120 = 7'h9 == total_offset_54[6:0] ? phv_data_9 : _GEN_3119; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3121 = 7'ha == total_offset_54[6:0] ? phv_data_10 : _GEN_3120; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3122 = 7'hb == total_offset_54[6:0] ? phv_data_11 : _GEN_3121; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3123 = 7'hc == total_offset_54[6:0] ? phv_data_12 : _GEN_3122; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3124 = 7'hd == total_offset_54[6:0] ? phv_data_13 : _GEN_3123; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3125 = 7'he == total_offset_54[6:0] ? phv_data_14 : _GEN_3124; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3126 = 7'hf == total_offset_54[6:0] ? phv_data_15 : _GEN_3125; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3127 = 7'h10 == total_offset_54[6:0] ? phv_data_16 : _GEN_3126; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3128 = 7'h11 == total_offset_54[6:0] ? phv_data_17 : _GEN_3127; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3129 = 7'h12 == total_offset_54[6:0] ? phv_data_18 : _GEN_3128; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3130 = 7'h13 == total_offset_54[6:0] ? phv_data_19 : _GEN_3129; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3131 = 7'h14 == total_offset_54[6:0] ? phv_data_20 : _GEN_3130; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3132 = 7'h15 == total_offset_54[6:0] ? phv_data_21 : _GEN_3131; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3133 = 7'h16 == total_offset_54[6:0] ? phv_data_22 : _GEN_3132; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3134 = 7'h17 == total_offset_54[6:0] ? phv_data_23 : _GEN_3133; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3135 = 7'h18 == total_offset_54[6:0] ? phv_data_24 : _GEN_3134; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3136 = 7'h19 == total_offset_54[6:0] ? phv_data_25 : _GEN_3135; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3137 = 7'h1a == total_offset_54[6:0] ? phv_data_26 : _GEN_3136; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3138 = 7'h1b == total_offset_54[6:0] ? phv_data_27 : _GEN_3137; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3139 = 7'h1c == total_offset_54[6:0] ? phv_data_28 : _GEN_3138; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3140 = 7'h1d == total_offset_54[6:0] ? phv_data_29 : _GEN_3139; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3141 = 7'h1e == total_offset_54[6:0] ? phv_data_30 : _GEN_3140; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3142 = 7'h1f == total_offset_54[6:0] ? phv_data_31 : _GEN_3141; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3143 = 7'h20 == total_offset_54[6:0] ? phv_data_32 : _GEN_3142; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3144 = 7'h21 == total_offset_54[6:0] ? phv_data_33 : _GEN_3143; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3145 = 7'h22 == total_offset_54[6:0] ? phv_data_34 : _GEN_3144; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3146 = 7'h23 == total_offset_54[6:0] ? phv_data_35 : _GEN_3145; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3147 = 7'h24 == total_offset_54[6:0] ? phv_data_36 : _GEN_3146; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3148 = 7'h25 == total_offset_54[6:0] ? phv_data_37 : _GEN_3147; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3149 = 7'h26 == total_offset_54[6:0] ? phv_data_38 : _GEN_3148; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3150 = 7'h27 == total_offset_54[6:0] ? phv_data_39 : _GEN_3149; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3151 = 7'h28 == total_offset_54[6:0] ? phv_data_40 : _GEN_3150; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3152 = 7'h29 == total_offset_54[6:0] ? phv_data_41 : _GEN_3151; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3153 = 7'h2a == total_offset_54[6:0] ? phv_data_42 : _GEN_3152; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3154 = 7'h2b == total_offset_54[6:0] ? phv_data_43 : _GEN_3153; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3155 = 7'h2c == total_offset_54[6:0] ? phv_data_44 : _GEN_3154; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3156 = 7'h2d == total_offset_54[6:0] ? phv_data_45 : _GEN_3155; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3157 = 7'h2e == total_offset_54[6:0] ? phv_data_46 : _GEN_3156; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3158 = 7'h2f == total_offset_54[6:0] ? phv_data_47 : _GEN_3157; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3159 = 7'h30 == total_offset_54[6:0] ? phv_data_48 : _GEN_3158; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3160 = 7'h31 == total_offset_54[6:0] ? phv_data_49 : _GEN_3159; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3161 = 7'h32 == total_offset_54[6:0] ? phv_data_50 : _GEN_3160; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3162 = 7'h33 == total_offset_54[6:0] ? phv_data_51 : _GEN_3161; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3163 = 7'h34 == total_offset_54[6:0] ? phv_data_52 : _GEN_3162; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3164 = 7'h35 == total_offset_54[6:0] ? phv_data_53 : _GEN_3163; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3165 = 7'h36 == total_offset_54[6:0] ? phv_data_54 : _GEN_3164; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3166 = 7'h37 == total_offset_54[6:0] ? phv_data_55 : _GEN_3165; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3167 = 7'h38 == total_offset_54[6:0] ? phv_data_56 : _GEN_3166; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3168 = 7'h39 == total_offset_54[6:0] ? phv_data_57 : _GEN_3167; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3169 = 7'h3a == total_offset_54[6:0] ? phv_data_58 : _GEN_3168; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3170 = 7'h3b == total_offset_54[6:0] ? phv_data_59 : _GEN_3169; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3171 = 7'h3c == total_offset_54[6:0] ? phv_data_60 : _GEN_3170; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3172 = 7'h3d == total_offset_54[6:0] ? phv_data_61 : _GEN_3171; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3173 = 7'h3e == total_offset_54[6:0] ? phv_data_62 : _GEN_3172; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3174 = 7'h3f == total_offset_54[6:0] ? phv_data_63 : _GEN_3173; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3175 = 7'h40 == total_offset_54[6:0] ? phv_data_64 : _GEN_3174; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3176 = 7'h41 == total_offset_54[6:0] ? phv_data_65 : _GEN_3175; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3177 = 7'h42 == total_offset_54[6:0] ? phv_data_66 : _GEN_3176; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3178 = 7'h43 == total_offset_54[6:0] ? phv_data_67 : _GEN_3177; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3179 = 7'h44 == total_offset_54[6:0] ? phv_data_68 : _GEN_3178; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3180 = 7'h45 == total_offset_54[6:0] ? phv_data_69 : _GEN_3179; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3181 = 7'h46 == total_offset_54[6:0] ? phv_data_70 : _GEN_3180; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3182 = 7'h47 == total_offset_54[6:0] ? phv_data_71 : _GEN_3181; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3183 = 7'h48 == total_offset_54[6:0] ? phv_data_72 : _GEN_3182; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3184 = 7'h49 == total_offset_54[6:0] ? phv_data_73 : _GEN_3183; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3185 = 7'h4a == total_offset_54[6:0] ? phv_data_74 : _GEN_3184; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3186 = 7'h4b == total_offset_54[6:0] ? phv_data_75 : _GEN_3185; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3187 = 7'h4c == total_offset_54[6:0] ? phv_data_76 : _GEN_3186; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3188 = 7'h4d == total_offset_54[6:0] ? phv_data_77 : _GEN_3187; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3189 = 7'h4e == total_offset_54[6:0] ? phv_data_78 : _GEN_3188; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3190 = 7'h4f == total_offset_54[6:0] ? phv_data_79 : _GEN_3189; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3191 = 7'h50 == total_offset_54[6:0] ? phv_data_80 : _GEN_3190; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3192 = 7'h51 == total_offset_54[6:0] ? phv_data_81 : _GEN_3191; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3193 = 7'h52 == total_offset_54[6:0] ? phv_data_82 : _GEN_3192; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3194 = 7'h53 == total_offset_54[6:0] ? phv_data_83 : _GEN_3193; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3195 = 7'h54 == total_offset_54[6:0] ? phv_data_84 : _GEN_3194; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3196 = 7'h55 == total_offset_54[6:0] ? phv_data_85 : _GEN_3195; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3197 = 7'h56 == total_offset_54[6:0] ? phv_data_86 : _GEN_3196; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3198 = 7'h57 == total_offset_54[6:0] ? phv_data_87 : _GEN_3197; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3199 = 7'h58 == total_offset_54[6:0] ? phv_data_88 : _GEN_3198; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3200 = 7'h59 == total_offset_54[6:0] ? phv_data_89 : _GEN_3199; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3201 = 7'h5a == total_offset_54[6:0] ? phv_data_90 : _GEN_3200; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3202 = 7'h5b == total_offset_54[6:0] ? phv_data_91 : _GEN_3201; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3203 = 7'h5c == total_offset_54[6:0] ? phv_data_92 : _GEN_3202; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3204 = 7'h5d == total_offset_54[6:0] ? phv_data_93 : _GEN_3203; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3205 = 7'h5e == total_offset_54[6:0] ? phv_data_94 : _GEN_3204; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3206 = 7'h5f == total_offset_54[6:0] ? phv_data_95 : _GEN_3205; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes_6_6 = 8'h6 < length_3 ? _GEN_3206 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [7:0] total_offset_55 = offset_3 + 8'h7; // @[executor.scala 158:57]
  wire [7:0] _GEN_3209 = 7'h1 == total_offset_55[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3210 = 7'h2 == total_offset_55[6:0] ? phv_data_2 : _GEN_3209; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3211 = 7'h3 == total_offset_55[6:0] ? phv_data_3 : _GEN_3210; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3212 = 7'h4 == total_offset_55[6:0] ? phv_data_4 : _GEN_3211; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3213 = 7'h5 == total_offset_55[6:0] ? phv_data_5 : _GEN_3212; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3214 = 7'h6 == total_offset_55[6:0] ? phv_data_6 : _GEN_3213; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3215 = 7'h7 == total_offset_55[6:0] ? phv_data_7 : _GEN_3214; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3216 = 7'h8 == total_offset_55[6:0] ? phv_data_8 : _GEN_3215; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3217 = 7'h9 == total_offset_55[6:0] ? phv_data_9 : _GEN_3216; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3218 = 7'ha == total_offset_55[6:0] ? phv_data_10 : _GEN_3217; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3219 = 7'hb == total_offset_55[6:0] ? phv_data_11 : _GEN_3218; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3220 = 7'hc == total_offset_55[6:0] ? phv_data_12 : _GEN_3219; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3221 = 7'hd == total_offset_55[6:0] ? phv_data_13 : _GEN_3220; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3222 = 7'he == total_offset_55[6:0] ? phv_data_14 : _GEN_3221; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3223 = 7'hf == total_offset_55[6:0] ? phv_data_15 : _GEN_3222; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3224 = 7'h10 == total_offset_55[6:0] ? phv_data_16 : _GEN_3223; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3225 = 7'h11 == total_offset_55[6:0] ? phv_data_17 : _GEN_3224; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3226 = 7'h12 == total_offset_55[6:0] ? phv_data_18 : _GEN_3225; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3227 = 7'h13 == total_offset_55[6:0] ? phv_data_19 : _GEN_3226; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3228 = 7'h14 == total_offset_55[6:0] ? phv_data_20 : _GEN_3227; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3229 = 7'h15 == total_offset_55[6:0] ? phv_data_21 : _GEN_3228; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3230 = 7'h16 == total_offset_55[6:0] ? phv_data_22 : _GEN_3229; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3231 = 7'h17 == total_offset_55[6:0] ? phv_data_23 : _GEN_3230; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3232 = 7'h18 == total_offset_55[6:0] ? phv_data_24 : _GEN_3231; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3233 = 7'h19 == total_offset_55[6:0] ? phv_data_25 : _GEN_3232; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3234 = 7'h1a == total_offset_55[6:0] ? phv_data_26 : _GEN_3233; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3235 = 7'h1b == total_offset_55[6:0] ? phv_data_27 : _GEN_3234; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3236 = 7'h1c == total_offset_55[6:0] ? phv_data_28 : _GEN_3235; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3237 = 7'h1d == total_offset_55[6:0] ? phv_data_29 : _GEN_3236; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3238 = 7'h1e == total_offset_55[6:0] ? phv_data_30 : _GEN_3237; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3239 = 7'h1f == total_offset_55[6:0] ? phv_data_31 : _GEN_3238; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3240 = 7'h20 == total_offset_55[6:0] ? phv_data_32 : _GEN_3239; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3241 = 7'h21 == total_offset_55[6:0] ? phv_data_33 : _GEN_3240; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3242 = 7'h22 == total_offset_55[6:0] ? phv_data_34 : _GEN_3241; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3243 = 7'h23 == total_offset_55[6:0] ? phv_data_35 : _GEN_3242; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3244 = 7'h24 == total_offset_55[6:0] ? phv_data_36 : _GEN_3243; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3245 = 7'h25 == total_offset_55[6:0] ? phv_data_37 : _GEN_3244; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3246 = 7'h26 == total_offset_55[6:0] ? phv_data_38 : _GEN_3245; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3247 = 7'h27 == total_offset_55[6:0] ? phv_data_39 : _GEN_3246; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3248 = 7'h28 == total_offset_55[6:0] ? phv_data_40 : _GEN_3247; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3249 = 7'h29 == total_offset_55[6:0] ? phv_data_41 : _GEN_3248; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3250 = 7'h2a == total_offset_55[6:0] ? phv_data_42 : _GEN_3249; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3251 = 7'h2b == total_offset_55[6:0] ? phv_data_43 : _GEN_3250; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3252 = 7'h2c == total_offset_55[6:0] ? phv_data_44 : _GEN_3251; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3253 = 7'h2d == total_offset_55[6:0] ? phv_data_45 : _GEN_3252; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3254 = 7'h2e == total_offset_55[6:0] ? phv_data_46 : _GEN_3253; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3255 = 7'h2f == total_offset_55[6:0] ? phv_data_47 : _GEN_3254; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3256 = 7'h30 == total_offset_55[6:0] ? phv_data_48 : _GEN_3255; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3257 = 7'h31 == total_offset_55[6:0] ? phv_data_49 : _GEN_3256; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3258 = 7'h32 == total_offset_55[6:0] ? phv_data_50 : _GEN_3257; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3259 = 7'h33 == total_offset_55[6:0] ? phv_data_51 : _GEN_3258; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3260 = 7'h34 == total_offset_55[6:0] ? phv_data_52 : _GEN_3259; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3261 = 7'h35 == total_offset_55[6:0] ? phv_data_53 : _GEN_3260; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3262 = 7'h36 == total_offset_55[6:0] ? phv_data_54 : _GEN_3261; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3263 = 7'h37 == total_offset_55[6:0] ? phv_data_55 : _GEN_3262; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3264 = 7'h38 == total_offset_55[6:0] ? phv_data_56 : _GEN_3263; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3265 = 7'h39 == total_offset_55[6:0] ? phv_data_57 : _GEN_3264; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3266 = 7'h3a == total_offset_55[6:0] ? phv_data_58 : _GEN_3265; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3267 = 7'h3b == total_offset_55[6:0] ? phv_data_59 : _GEN_3266; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3268 = 7'h3c == total_offset_55[6:0] ? phv_data_60 : _GEN_3267; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3269 = 7'h3d == total_offset_55[6:0] ? phv_data_61 : _GEN_3268; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3270 = 7'h3e == total_offset_55[6:0] ? phv_data_62 : _GEN_3269; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3271 = 7'h3f == total_offset_55[6:0] ? phv_data_63 : _GEN_3270; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3272 = 7'h40 == total_offset_55[6:0] ? phv_data_64 : _GEN_3271; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3273 = 7'h41 == total_offset_55[6:0] ? phv_data_65 : _GEN_3272; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3274 = 7'h42 == total_offset_55[6:0] ? phv_data_66 : _GEN_3273; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3275 = 7'h43 == total_offset_55[6:0] ? phv_data_67 : _GEN_3274; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3276 = 7'h44 == total_offset_55[6:0] ? phv_data_68 : _GEN_3275; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3277 = 7'h45 == total_offset_55[6:0] ? phv_data_69 : _GEN_3276; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3278 = 7'h46 == total_offset_55[6:0] ? phv_data_70 : _GEN_3277; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3279 = 7'h47 == total_offset_55[6:0] ? phv_data_71 : _GEN_3278; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3280 = 7'h48 == total_offset_55[6:0] ? phv_data_72 : _GEN_3279; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3281 = 7'h49 == total_offset_55[6:0] ? phv_data_73 : _GEN_3280; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3282 = 7'h4a == total_offset_55[6:0] ? phv_data_74 : _GEN_3281; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3283 = 7'h4b == total_offset_55[6:0] ? phv_data_75 : _GEN_3282; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3284 = 7'h4c == total_offset_55[6:0] ? phv_data_76 : _GEN_3283; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3285 = 7'h4d == total_offset_55[6:0] ? phv_data_77 : _GEN_3284; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3286 = 7'h4e == total_offset_55[6:0] ? phv_data_78 : _GEN_3285; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3287 = 7'h4f == total_offset_55[6:0] ? phv_data_79 : _GEN_3286; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3288 = 7'h50 == total_offset_55[6:0] ? phv_data_80 : _GEN_3287; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3289 = 7'h51 == total_offset_55[6:0] ? phv_data_81 : _GEN_3288; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3290 = 7'h52 == total_offset_55[6:0] ? phv_data_82 : _GEN_3289; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3291 = 7'h53 == total_offset_55[6:0] ? phv_data_83 : _GEN_3290; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3292 = 7'h54 == total_offset_55[6:0] ? phv_data_84 : _GEN_3291; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3293 = 7'h55 == total_offset_55[6:0] ? phv_data_85 : _GEN_3292; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3294 = 7'h56 == total_offset_55[6:0] ? phv_data_86 : _GEN_3293; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3295 = 7'h57 == total_offset_55[6:0] ? phv_data_87 : _GEN_3294; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3296 = 7'h58 == total_offset_55[6:0] ? phv_data_88 : _GEN_3295; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3297 = 7'h59 == total_offset_55[6:0] ? phv_data_89 : _GEN_3296; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3298 = 7'h5a == total_offset_55[6:0] ? phv_data_90 : _GEN_3297; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3299 = 7'h5b == total_offset_55[6:0] ? phv_data_91 : _GEN_3298; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3300 = 7'h5c == total_offset_55[6:0] ? phv_data_92 : _GEN_3299; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3301 = 7'h5d == total_offset_55[6:0] ? phv_data_93 : _GEN_3300; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3302 = 7'h5e == total_offset_55[6:0] ? phv_data_94 : _GEN_3301; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] _GEN_3303 = 7'h5f == total_offset_55[6:0] ? phv_data_95 : _GEN_3302; // @[executor.scala 160:38 executor.scala 160:38]
  wire [7:0] bytes_6_7 = 8'h7 < length_3 ? _GEN_3303 : 8'h0; // @[executor.scala 159:60 executor.scala 160:38 executor.scala 162:38]
  wire [63:0] _io_field_out_3_T = {bytes_6_0,bytes_6_1,bytes_6_2,bytes_6_3,bytes_6_4,bytes_6_5,bytes_6_6,bytes_6_7}; // @[Cat.scala 30:58]
  wire [2:0] args_offset_3 = io_field_out_3_lo[13:11]; // @[primitive.scala 34:52]
  wire [2:0] args_length_3 = io_field_out_3_lo[10:8]; // @[primitive.scala 35:52]
  wire [8:0] _total_offset_T_56 = {{6'd0}, args_offset_3}; // @[executor.scala 173:60]
  wire [7:0] total_offset_56 = _total_offset_T_56[7:0]; // @[executor.scala 173:60]
  wire [7:0] _GEN_3414 = {{5'd0}, args_length_3}; // @[executor.scala 174:48]
  wire [7:0] _GEN_3306 = 3'h1 == total_offset_56[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3307 = 3'h2 == total_offset_56[2:0] ? args_2 : _GEN_3306; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3308 = 3'h3 == total_offset_56[2:0] ? args_3 : _GEN_3307; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3309 = 3'h4 == total_offset_56[2:0] ? args_4 : _GEN_3308; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3310 = 3'h5 == total_offset_56[2:0] ? args_5 : _GEN_3309; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3311 = 3'h6 == total_offset_56[2:0] ? args_6 : _GEN_3310; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_7_0 = 8'h0 < _GEN_3414 ? _GEN_3311 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [7:0] _GEN_3415 = {{5'd0}, args_offset_3}; // @[executor.scala 173:60]
  wire [7:0] total_offset_57 = _GEN_3415 + 8'h1; // @[executor.scala 173:60]
  wire [7:0] _GEN_3314 = 3'h1 == total_offset_57[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3315 = 3'h2 == total_offset_57[2:0] ? args_2 : _GEN_3314; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3316 = 3'h3 == total_offset_57[2:0] ? args_3 : _GEN_3315; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3317 = 3'h4 == total_offset_57[2:0] ? args_4 : _GEN_3316; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3318 = 3'h5 == total_offset_57[2:0] ? args_5 : _GEN_3317; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3319 = 3'h6 == total_offset_57[2:0] ? args_6 : _GEN_3318; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_7_1 = 8'h1 < _GEN_3414 ? _GEN_3319 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [7:0] total_offset_58 = _GEN_3415 + 8'h2; // @[executor.scala 173:60]
  wire [7:0] _GEN_3322 = 3'h1 == total_offset_58[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3323 = 3'h2 == total_offset_58[2:0] ? args_2 : _GEN_3322; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3324 = 3'h3 == total_offset_58[2:0] ? args_3 : _GEN_3323; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3325 = 3'h4 == total_offset_58[2:0] ? args_4 : _GEN_3324; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3326 = 3'h5 == total_offset_58[2:0] ? args_5 : _GEN_3325; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3327 = 3'h6 == total_offset_58[2:0] ? args_6 : _GEN_3326; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_7_2 = 8'h2 < _GEN_3414 ? _GEN_3327 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [7:0] total_offset_59 = _GEN_3415 + 8'h3; // @[executor.scala 173:60]
  wire [7:0] _GEN_3330 = 3'h1 == total_offset_59[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3331 = 3'h2 == total_offset_59[2:0] ? args_2 : _GEN_3330; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3332 = 3'h3 == total_offset_59[2:0] ? args_3 : _GEN_3331; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3333 = 3'h4 == total_offset_59[2:0] ? args_4 : _GEN_3332; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3334 = 3'h5 == total_offset_59[2:0] ? args_5 : _GEN_3333; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3335 = 3'h6 == total_offset_59[2:0] ? args_6 : _GEN_3334; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_7_3 = 8'h3 < _GEN_3414 ? _GEN_3335 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [7:0] total_offset_60 = _GEN_3415 + 8'h4; // @[executor.scala 173:60]
  wire [7:0] _GEN_3338 = 3'h1 == total_offset_60[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3339 = 3'h2 == total_offset_60[2:0] ? args_2 : _GEN_3338; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3340 = 3'h3 == total_offset_60[2:0] ? args_3 : _GEN_3339; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3341 = 3'h4 == total_offset_60[2:0] ? args_4 : _GEN_3340; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3342 = 3'h5 == total_offset_60[2:0] ? args_5 : _GEN_3341; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3343 = 3'h6 == total_offset_60[2:0] ? args_6 : _GEN_3342; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_7_4 = 8'h4 < _GEN_3414 ? _GEN_3343 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [7:0] total_offset_61 = _GEN_3415 + 8'h5; // @[executor.scala 173:60]
  wire [7:0] _GEN_3346 = 3'h1 == total_offset_61[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3347 = 3'h2 == total_offset_61[2:0] ? args_2 : _GEN_3346; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3348 = 3'h3 == total_offset_61[2:0] ? args_3 : _GEN_3347; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3349 = 3'h4 == total_offset_61[2:0] ? args_4 : _GEN_3348; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3350 = 3'h5 == total_offset_61[2:0] ? args_5 : _GEN_3349; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3351 = 3'h6 == total_offset_61[2:0] ? args_6 : _GEN_3350; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_7_5 = 8'h5 < _GEN_3414 ? _GEN_3351 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [7:0] total_offset_62 = _GEN_3415 + 8'h6; // @[executor.scala 173:60]
  wire [7:0] _GEN_3354 = 3'h1 == total_offset_62[2:0] ? args_1 : args_0; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3355 = 3'h2 == total_offset_62[2:0] ? args_2 : _GEN_3354; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3356 = 3'h3 == total_offset_62[2:0] ? args_3 : _GEN_3355; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3357 = 3'h4 == total_offset_62[2:0] ? args_4 : _GEN_3356; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3358 = 3'h5 == total_offset_62[2:0] ? args_5 : _GEN_3357; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] _GEN_3359 = 3'h6 == total_offset_62[2:0] ? args_6 : _GEN_3358; // @[executor.scala 175:42 executor.scala 175:42]
  wire [7:0] bytes_7_6 = 8'h6 < _GEN_3414 ? _GEN_3359 : 8'h0; // @[executor.scala 174:63 executor.scala 175:42 executor.scala 177:42]
  wire [63:0] _io_field_out_3_T_1 = {bytes_7_0,bytes_7_1,bytes_7_2,bytes_7_3,bytes_7_4,bytes_7_5,bytes_7_6,8'h0}; // @[Cat.scala 30:58]
  wire [49:0] io_field_out_3_hi_12 = io_field_out_3_lo[13] ? 50'h3ffffffffffff : 50'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _io_field_out_3_T_4 = {io_field_out_3_hi_12,io_field_out_3_lo}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_3369 = 4'ha == opcode_3 ? _io_field_out_3_T_1 : _io_field_out_3_T_4; // @[executor.scala 167:55 executor.scala 180:41 executor.scala 183:41]
  wire [63:0] _GEN_3370 = from_header_3 ? _io_field_out_3_T : _GEN_3369; // @[executor.scala 152:36 executor.scala 165:37]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[executor.scala 130:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[executor.scala 130:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[executor.scala 130:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[executor.scala 130:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[executor.scala 130:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[executor.scala 130:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[executor.scala 130:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[executor.scala 130:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[executor.scala 130:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[executor.scala 130:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[executor.scala 130:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[executor.scala 130:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[executor.scala 130:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[executor.scala 130:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[executor.scala 130:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[executor.scala 130:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[executor.scala 130:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[executor.scala 130:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[executor.scala 130:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[executor.scala 130:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[executor.scala 130:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[executor.scala 130:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[executor.scala 130:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[executor.scala 130:25]
  assign io_vliw_out_0 = vliw_0; // @[executor.scala 137:21]
  assign io_vliw_out_1 = vliw_1; // @[executor.scala 137:21]
  assign io_vliw_out_2 = vliw_2; // @[executor.scala 137:21]
  assign io_vliw_out_3 = vliw_3; // @[executor.scala 137:21]
  assign io_field_out_0 = phv_is_valid_processor ? _GEN_841 : 64'h0; // @[executor.scala 150:43 executor.scala 149:29]
  assign io_field_out_1 = phv_is_valid_processor ? _GEN_1684 : 64'h0; // @[executor.scala 150:43 executor.scala 149:29]
  assign io_field_out_2 = phv_is_valid_processor ? _GEN_2527 : 64'h0; // @[executor.scala 150:43 executor.scala 149:29]
  assign io_field_out_3 = phv_is_valid_processor ? _GEN_3370 : 64'h0; // @[executor.scala 150:43 executor.scala 149:29]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[executor.scala 129:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[executor.scala 129:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[executor.scala 129:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[executor.scala 129:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[executor.scala 129:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[executor.scala 129:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[executor.scala 129:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[executor.scala 129:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[executor.scala 129:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[executor.scala 129:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[executor.scala 129:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[executor.scala 129:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[executor.scala 129:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[executor.scala 129:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[executor.scala 129:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[executor.scala 129:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[executor.scala 129:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[executor.scala 129:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[executor.scala 129:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[executor.scala 129:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[executor.scala 129:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[executor.scala 129:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[executor.scala 129:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[executor.scala 129:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[executor.scala 129:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[executor.scala 129:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[executor.scala 129:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[executor.scala 129:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[executor.scala 129:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[executor.scala 129:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[executor.scala 129:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[executor.scala 129:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[executor.scala 129:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[executor.scala 129:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[executor.scala 129:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[executor.scala 129:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[executor.scala 129:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[executor.scala 129:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[executor.scala 129:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[executor.scala 129:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[executor.scala 129:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[executor.scala 129:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[executor.scala 129:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[executor.scala 129:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[executor.scala 129:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[executor.scala 129:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[executor.scala 129:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[executor.scala 129:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[executor.scala 129:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[executor.scala 129:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[executor.scala 129:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[executor.scala 129:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[executor.scala 129:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[executor.scala 129:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[executor.scala 129:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[executor.scala 129:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[executor.scala 129:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[executor.scala 129:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[executor.scala 129:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[executor.scala 129:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[executor.scala 129:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[executor.scala 129:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[executor.scala 129:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[executor.scala 129:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[executor.scala 129:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[executor.scala 129:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[executor.scala 129:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[executor.scala 129:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[executor.scala 129:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[executor.scala 129:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[executor.scala 129:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[executor.scala 129:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[executor.scala 129:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[executor.scala 129:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[executor.scala 129:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[executor.scala 129:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[executor.scala 129:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[executor.scala 129:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[executor.scala 129:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[executor.scala 129:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[executor.scala 129:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[executor.scala 129:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[executor.scala 129:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[executor.scala 129:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[executor.scala 129:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[executor.scala 129:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[executor.scala 129:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[executor.scala 129:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[executor.scala 129:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[executor.scala 129:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[executor.scala 129:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[executor.scala 129:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[executor.scala 129:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[executor.scala 129:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[executor.scala 129:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[executor.scala 129:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[executor.scala 129:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[executor.scala 129:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[executor.scala 129:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[executor.scala 129:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[executor.scala 129:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[executor.scala 129:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[executor.scala 129:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[executor.scala 129:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[executor.scala 129:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[executor.scala 129:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[executor.scala 129:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[executor.scala 129:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[executor.scala 129:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[executor.scala 129:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[executor.scala 129:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[executor.scala 129:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[executor.scala 129:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[executor.scala 129:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[executor.scala 129:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[executor.scala 129:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[executor.scala 129:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[executor.scala 129:13]
    args_0 <= io_args_in_0; // @[executor.scala 133:14]
    args_1 <= io_args_in_1; // @[executor.scala 133:14]
    args_2 <= io_args_in_2; // @[executor.scala 133:14]
    args_3 <= io_args_in_3; // @[executor.scala 133:14]
    args_4 <= io_args_in_4; // @[executor.scala 133:14]
    args_5 <= io_args_in_5; // @[executor.scala 133:14]
    args_6 <= io_args_in_6; // @[executor.scala 133:14]
    vliw_0 <= io_vliw_in_0; // @[executor.scala 136:14]
    vliw_1 <= io_vliw_in_1; // @[executor.scala 136:14]
    vliw_2 <= io_vliw_in_2; // @[executor.scala 136:14]
    vliw_3 <= io_vliw_in_3; // @[executor.scala 136:14]
    offset_0 <= io_offset_in_0; // @[executor.scala 141:16]
    offset_1 <= io_offset_in_1; // @[executor.scala 141:16]
    offset_2 <= io_offset_in_2; // @[executor.scala 141:16]
    offset_3 <= io_offset_in_3; // @[executor.scala 141:16]
    length_0 <= io_length_in_0; // @[executor.scala 142:16]
    length_1 <= io_length_in_1; // @[executor.scala 142:16]
    length_2 <= io_length_in_2; // @[executor.scala 142:16]
    length_3 <= io_length_in_3; // @[executor.scala 142:16]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_header_0 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  phv_header_1 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  phv_header_2 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  phv_header_3 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  phv_header_4 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  phv_header_5 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  phv_header_6 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  phv_header_7 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  phv_header_8 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  phv_header_9 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  phv_header_10 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  phv_header_11 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  phv_header_12 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  phv_header_13 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  phv_header_14 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  phv_header_15 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  phv_next_config_id = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  args_0 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  args_1 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  args_2 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  args_3 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  args_4 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  args_5 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  args_6 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  vliw_0 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  vliw_1 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  vliw_2 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  vliw_3 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  offset_0 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  offset_1 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  offset_2 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  offset_3 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  length_0 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  length_1 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  length_2 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  length_3 = _RAND_136[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
