module Processor(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [7:0]  io_pipe_phv_in_data_160,
  input  [7:0]  io_pipe_phv_in_data_161,
  input  [7:0]  io_pipe_phv_in_data_162,
  input  [7:0]  io_pipe_phv_in_data_163,
  input  [7:0]  io_pipe_phv_in_data_164,
  input  [7:0]  io_pipe_phv_in_data_165,
  input  [7:0]  io_pipe_phv_in_data_166,
  input  [7:0]  io_pipe_phv_in_data_167,
  input  [7:0]  io_pipe_phv_in_data_168,
  input  [7:0]  io_pipe_phv_in_data_169,
  input  [7:0]  io_pipe_phv_in_data_170,
  input  [7:0]  io_pipe_phv_in_data_171,
  input  [7:0]  io_pipe_phv_in_data_172,
  input  [7:0]  io_pipe_phv_in_data_173,
  input  [7:0]  io_pipe_phv_in_data_174,
  input  [7:0]  io_pipe_phv_in_data_175,
  input  [7:0]  io_pipe_phv_in_data_176,
  input  [7:0]  io_pipe_phv_in_data_177,
  input  [7:0]  io_pipe_phv_in_data_178,
  input  [7:0]  io_pipe_phv_in_data_179,
  input  [7:0]  io_pipe_phv_in_data_180,
  input  [7:0]  io_pipe_phv_in_data_181,
  input  [7:0]  io_pipe_phv_in_data_182,
  input  [7:0]  io_pipe_phv_in_data_183,
  input  [7:0]  io_pipe_phv_in_data_184,
  input  [7:0]  io_pipe_phv_in_data_185,
  input  [7:0]  io_pipe_phv_in_data_186,
  input  [7:0]  io_pipe_phv_in_data_187,
  input  [7:0]  io_pipe_phv_in_data_188,
  input  [7:0]  io_pipe_phv_in_data_189,
  input  [7:0]  io_pipe_phv_in_data_190,
  input  [7:0]  io_pipe_phv_in_data_191,
  input  [7:0]  io_pipe_phv_in_data_192,
  input  [7:0]  io_pipe_phv_in_data_193,
  input  [7:0]  io_pipe_phv_in_data_194,
  input  [7:0]  io_pipe_phv_in_data_195,
  input  [7:0]  io_pipe_phv_in_data_196,
  input  [7:0]  io_pipe_phv_in_data_197,
  input  [7:0]  io_pipe_phv_in_data_198,
  input  [7:0]  io_pipe_phv_in_data_199,
  input  [7:0]  io_pipe_phv_in_data_200,
  input  [7:0]  io_pipe_phv_in_data_201,
  input  [7:0]  io_pipe_phv_in_data_202,
  input  [7:0]  io_pipe_phv_in_data_203,
  input  [7:0]  io_pipe_phv_in_data_204,
  input  [7:0]  io_pipe_phv_in_data_205,
  input  [7:0]  io_pipe_phv_in_data_206,
  input  [7:0]  io_pipe_phv_in_data_207,
  input  [7:0]  io_pipe_phv_in_data_208,
  input  [7:0]  io_pipe_phv_in_data_209,
  input  [7:0]  io_pipe_phv_in_data_210,
  input  [7:0]  io_pipe_phv_in_data_211,
  input  [7:0]  io_pipe_phv_in_data_212,
  input  [7:0]  io_pipe_phv_in_data_213,
  input  [7:0]  io_pipe_phv_in_data_214,
  input  [7:0]  io_pipe_phv_in_data_215,
  input  [7:0]  io_pipe_phv_in_data_216,
  input  [7:0]  io_pipe_phv_in_data_217,
  input  [7:0]  io_pipe_phv_in_data_218,
  input  [7:0]  io_pipe_phv_in_data_219,
  input  [7:0]  io_pipe_phv_in_data_220,
  input  [7:0]  io_pipe_phv_in_data_221,
  input  [7:0]  io_pipe_phv_in_data_222,
  input  [7:0]  io_pipe_phv_in_data_223,
  input  [7:0]  io_pipe_phv_in_data_224,
  input  [7:0]  io_pipe_phv_in_data_225,
  input  [7:0]  io_pipe_phv_in_data_226,
  input  [7:0]  io_pipe_phv_in_data_227,
  input  [7:0]  io_pipe_phv_in_data_228,
  input  [7:0]  io_pipe_phv_in_data_229,
  input  [7:0]  io_pipe_phv_in_data_230,
  input  [7:0]  io_pipe_phv_in_data_231,
  input  [7:0]  io_pipe_phv_in_data_232,
  input  [7:0]  io_pipe_phv_in_data_233,
  input  [7:0]  io_pipe_phv_in_data_234,
  input  [7:0]  io_pipe_phv_in_data_235,
  input  [7:0]  io_pipe_phv_in_data_236,
  input  [7:0]  io_pipe_phv_in_data_237,
  input  [7:0]  io_pipe_phv_in_data_238,
  input  [7:0]  io_pipe_phv_in_data_239,
  input  [7:0]  io_pipe_phv_in_data_240,
  input  [7:0]  io_pipe_phv_in_data_241,
  input  [7:0]  io_pipe_phv_in_data_242,
  input  [7:0]  io_pipe_phv_in_data_243,
  input  [7:0]  io_pipe_phv_in_data_244,
  input  [7:0]  io_pipe_phv_in_data_245,
  input  [7:0]  io_pipe_phv_in_data_246,
  input  [7:0]  io_pipe_phv_in_data_247,
  input  [7:0]  io_pipe_phv_in_data_248,
  input  [7:0]  io_pipe_phv_in_data_249,
  input  [7:0]  io_pipe_phv_in_data_250,
  input  [7:0]  io_pipe_phv_in_data_251,
  input  [7:0]  io_pipe_phv_in_data_252,
  input  [7:0]  io_pipe_phv_in_data_253,
  input  [7:0]  io_pipe_phv_in_data_254,
  input  [7:0]  io_pipe_phv_in_data_255,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [2:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [7:0]  io_pipe_phv_out_data_160,
  output [7:0]  io_pipe_phv_out_data_161,
  output [7:0]  io_pipe_phv_out_data_162,
  output [7:0]  io_pipe_phv_out_data_163,
  output [7:0]  io_pipe_phv_out_data_164,
  output [7:0]  io_pipe_phv_out_data_165,
  output [7:0]  io_pipe_phv_out_data_166,
  output [7:0]  io_pipe_phv_out_data_167,
  output [7:0]  io_pipe_phv_out_data_168,
  output [7:0]  io_pipe_phv_out_data_169,
  output [7:0]  io_pipe_phv_out_data_170,
  output [7:0]  io_pipe_phv_out_data_171,
  output [7:0]  io_pipe_phv_out_data_172,
  output [7:0]  io_pipe_phv_out_data_173,
  output [7:0]  io_pipe_phv_out_data_174,
  output [7:0]  io_pipe_phv_out_data_175,
  output [7:0]  io_pipe_phv_out_data_176,
  output [7:0]  io_pipe_phv_out_data_177,
  output [7:0]  io_pipe_phv_out_data_178,
  output [7:0]  io_pipe_phv_out_data_179,
  output [7:0]  io_pipe_phv_out_data_180,
  output [7:0]  io_pipe_phv_out_data_181,
  output [7:0]  io_pipe_phv_out_data_182,
  output [7:0]  io_pipe_phv_out_data_183,
  output [7:0]  io_pipe_phv_out_data_184,
  output [7:0]  io_pipe_phv_out_data_185,
  output [7:0]  io_pipe_phv_out_data_186,
  output [7:0]  io_pipe_phv_out_data_187,
  output [7:0]  io_pipe_phv_out_data_188,
  output [7:0]  io_pipe_phv_out_data_189,
  output [7:0]  io_pipe_phv_out_data_190,
  output [7:0]  io_pipe_phv_out_data_191,
  output [7:0]  io_pipe_phv_out_data_192,
  output [7:0]  io_pipe_phv_out_data_193,
  output [7:0]  io_pipe_phv_out_data_194,
  output [7:0]  io_pipe_phv_out_data_195,
  output [7:0]  io_pipe_phv_out_data_196,
  output [7:0]  io_pipe_phv_out_data_197,
  output [7:0]  io_pipe_phv_out_data_198,
  output [7:0]  io_pipe_phv_out_data_199,
  output [7:0]  io_pipe_phv_out_data_200,
  output [7:0]  io_pipe_phv_out_data_201,
  output [7:0]  io_pipe_phv_out_data_202,
  output [7:0]  io_pipe_phv_out_data_203,
  output [7:0]  io_pipe_phv_out_data_204,
  output [7:0]  io_pipe_phv_out_data_205,
  output [7:0]  io_pipe_phv_out_data_206,
  output [7:0]  io_pipe_phv_out_data_207,
  output [7:0]  io_pipe_phv_out_data_208,
  output [7:0]  io_pipe_phv_out_data_209,
  output [7:0]  io_pipe_phv_out_data_210,
  output [7:0]  io_pipe_phv_out_data_211,
  output [7:0]  io_pipe_phv_out_data_212,
  output [7:0]  io_pipe_phv_out_data_213,
  output [7:0]  io_pipe_phv_out_data_214,
  output [7:0]  io_pipe_phv_out_data_215,
  output [7:0]  io_pipe_phv_out_data_216,
  output [7:0]  io_pipe_phv_out_data_217,
  output [7:0]  io_pipe_phv_out_data_218,
  output [7:0]  io_pipe_phv_out_data_219,
  output [7:0]  io_pipe_phv_out_data_220,
  output [7:0]  io_pipe_phv_out_data_221,
  output [7:0]  io_pipe_phv_out_data_222,
  output [7:0]  io_pipe_phv_out_data_223,
  output [7:0]  io_pipe_phv_out_data_224,
  output [7:0]  io_pipe_phv_out_data_225,
  output [7:0]  io_pipe_phv_out_data_226,
  output [7:0]  io_pipe_phv_out_data_227,
  output [7:0]  io_pipe_phv_out_data_228,
  output [7:0]  io_pipe_phv_out_data_229,
  output [7:0]  io_pipe_phv_out_data_230,
  output [7:0]  io_pipe_phv_out_data_231,
  output [7:0]  io_pipe_phv_out_data_232,
  output [7:0]  io_pipe_phv_out_data_233,
  output [7:0]  io_pipe_phv_out_data_234,
  output [7:0]  io_pipe_phv_out_data_235,
  output [7:0]  io_pipe_phv_out_data_236,
  output [7:0]  io_pipe_phv_out_data_237,
  output [7:0]  io_pipe_phv_out_data_238,
  output [7:0]  io_pipe_phv_out_data_239,
  output [7:0]  io_pipe_phv_out_data_240,
  output [7:0]  io_pipe_phv_out_data_241,
  output [7:0]  io_pipe_phv_out_data_242,
  output [7:0]  io_pipe_phv_out_data_243,
  output [7:0]  io_pipe_phv_out_data_244,
  output [7:0]  io_pipe_phv_out_data_245,
  output [7:0]  io_pipe_phv_out_data_246,
  output [7:0]  io_pipe_phv_out_data_247,
  output [7:0]  io_pipe_phv_out_data_248,
  output [7:0]  io_pipe_phv_out_data_249,
  output [7:0]  io_pipe_phv_out_data_250,
  output [7:0]  io_pipe_phv_out_data_251,
  output [7:0]  io_pipe_phv_out_data_252,
  output [7:0]  io_pipe_phv_out_data_253,
  output [7:0]  io_pipe_phv_out_data_254,
  output [7:0]  io_pipe_phv_out_data_255,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [2:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  input         io_mod_par_mod_en,
  input         io_mod_par_mod_last_mau_id_mod,
  input  [1:0]  io_mod_par_mod_last_mau_id,
  input  [1:0]  io_mod_par_mod_cs,
  input         io_mod_par_mod_module_mod_state_id_mod,
  input  [7:0]  io_mod_par_mod_module_mod_state_id,
  input         io_mod_par_mod_module_mod_sram_w_cs,
  input         io_mod_par_mod_module_mod_sram_w_en,
  input  [7:0]  io_mod_par_mod_module_mod_sram_w_addr,
  input  [63:0] io_mod_par_mod_module_mod_sram_w_data,
  input         io_mod_mat_mod_en,
  input         io_mod_mat_mod_config_id,
  input  [7:0]  io_mod_mat_mod_key_mod_header_id,
  input  [7:0]  io_mod_mat_mod_key_mod_internal_offset,
  input  [7:0]  io_mod_mat_mod_key_mod_key_length,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_0,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_1,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_2,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_3,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_4,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_5,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_6,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_7,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_8,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_9,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_10,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_11,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_12,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_13,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_14,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_15,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_16,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_17,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_18,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_19,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_20,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_21,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_22,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_23,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_24,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_25,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_26,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_27,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_28,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_29,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_30,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_31,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_32,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_33,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_34,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_35,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_36,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_37,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_38,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_39,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_40,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_41,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_42,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_43,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_44,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_45,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_46,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_47,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_48,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_49,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_50,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_51,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_52,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_53,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_54,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_55,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_56,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_57,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_58,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_59,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_60,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_61,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_62,
  input  [5:0]  io_mod_mat_mod_table_mod_sram_id_table_63,
  input  [6:0]  io_mod_mat_mod_table_mod_table_width,
  input  [6:0]  io_mod_mat_mod_table_mod_table_depth,
  input         io_mod_act_mod_en_0,
  input         io_mod_act_mod_en_1,
  input  [7:0]  io_mod_act_mod_addr,
  input  [63:0] io_mod_act_mod_data_0,
  input  [63:0] io_mod_act_mod_data_1,
  output        io_mem_cluster_0_en,
  output [7:0]  io_mem_cluster_0_addr,
  input  [63:0] io_mem_cluster_0_data,
  output        io_mem_cluster_1_en,
  output [7:0]  io_mem_cluster_1_addr,
  input  [63:0] io_mem_cluster_1_data,
  output        io_mem_cluster_2_en,
  output [7:0]  io_mem_cluster_2_addr,
  input  [63:0] io_mem_cluster_2_data,
  output        io_mem_cluster_3_en,
  output [7:0]  io_mem_cluster_3_addr,
  input  [63:0] io_mem_cluster_3_data,
  output        io_mem_cluster_4_en,
  output [7:0]  io_mem_cluster_4_addr,
  input  [63:0] io_mem_cluster_4_data,
  output        io_mem_cluster_5_en,
  output [7:0]  io_mem_cluster_5_addr,
  input  [63:0] io_mem_cluster_5_data,
  output        io_mem_cluster_6_en,
  output [7:0]  io_mem_cluster_6_addr,
  input  [63:0] io_mem_cluster_6_data,
  output        io_mem_cluster_7_en,
  output [7:0]  io_mem_cluster_7_addr,
  input  [63:0] io_mem_cluster_7_data,
  output        io_mem_cluster_8_en,
  output [7:0]  io_mem_cluster_8_addr,
  input  [63:0] io_mem_cluster_8_data,
  output        io_mem_cluster_9_en,
  output [7:0]  io_mem_cluster_9_addr,
  input  [63:0] io_mem_cluster_9_data,
  output        io_mem_cluster_10_en,
  output [7:0]  io_mem_cluster_10_addr,
  input  [63:0] io_mem_cluster_10_data,
  output        io_mem_cluster_11_en,
  output [7:0]  io_mem_cluster_11_addr,
  input  [63:0] io_mem_cluster_11_data,
  output        io_mem_cluster_12_en,
  output [7:0]  io_mem_cluster_12_addr,
  input  [63:0] io_mem_cluster_12_data,
  output        io_mem_cluster_13_en,
  output [7:0]  io_mem_cluster_13_addr,
  input  [63:0] io_mem_cluster_13_data,
  output        io_mem_cluster_14_en,
  output [7:0]  io_mem_cluster_14_addr,
  input  [63:0] io_mem_cluster_14_data,
  output        io_mem_cluster_15_en,
  output [7:0]  io_mem_cluster_15_addr,
  input  [63:0] io_mem_cluster_15_data,
  output        io_mem_cluster_16_en,
  output [7:0]  io_mem_cluster_16_addr,
  input  [63:0] io_mem_cluster_16_data,
  output        io_mem_cluster_17_en,
  output [7:0]  io_mem_cluster_17_addr,
  input  [63:0] io_mem_cluster_17_data,
  output        io_mem_cluster_18_en,
  output [7:0]  io_mem_cluster_18_addr,
  input  [63:0] io_mem_cluster_18_data,
  output        io_mem_cluster_19_en,
  output [7:0]  io_mem_cluster_19_addr,
  input  [63:0] io_mem_cluster_19_data,
  output        io_mem_cluster_20_en,
  output [7:0]  io_mem_cluster_20_addr,
  input  [63:0] io_mem_cluster_20_data,
  output        io_mem_cluster_21_en,
  output [7:0]  io_mem_cluster_21_addr,
  input  [63:0] io_mem_cluster_21_data,
  output        io_mem_cluster_22_en,
  output [7:0]  io_mem_cluster_22_addr,
  input  [63:0] io_mem_cluster_22_data,
  output        io_mem_cluster_23_en,
  output [7:0]  io_mem_cluster_23_addr,
  input  [63:0] io_mem_cluster_23_data,
  output        io_mem_cluster_24_en,
  output [7:0]  io_mem_cluster_24_addr,
  input  [63:0] io_mem_cluster_24_data,
  output        io_mem_cluster_25_en,
  output [7:0]  io_mem_cluster_25_addr,
  input  [63:0] io_mem_cluster_25_data,
  output        io_mem_cluster_26_en,
  output [7:0]  io_mem_cluster_26_addr,
  input  [63:0] io_mem_cluster_26_data,
  output        io_mem_cluster_27_en,
  output [7:0]  io_mem_cluster_27_addr,
  input  [63:0] io_mem_cluster_27_data,
  output        io_mem_cluster_28_en,
  output [7:0]  io_mem_cluster_28_addr,
  input  [63:0] io_mem_cluster_28_data,
  output        io_mem_cluster_29_en,
  output [7:0]  io_mem_cluster_29_addr,
  input  [63:0] io_mem_cluster_29_data,
  output        io_mem_cluster_30_en,
  output [7:0]  io_mem_cluster_30_addr,
  input  [63:0] io_mem_cluster_30_data,
  output        io_mem_cluster_31_en,
  output [7:0]  io_mem_cluster_31_addr,
  input  [63:0] io_mem_cluster_31_data,
  output        io_mem_cluster_32_en,
  output [7:0]  io_mem_cluster_32_addr,
  input  [63:0] io_mem_cluster_32_data,
  output        io_mem_cluster_33_en,
  output [7:0]  io_mem_cluster_33_addr,
  input  [63:0] io_mem_cluster_33_data,
  output        io_mem_cluster_34_en,
  output [7:0]  io_mem_cluster_34_addr,
  input  [63:0] io_mem_cluster_34_data,
  output        io_mem_cluster_35_en,
  output [7:0]  io_mem_cluster_35_addr,
  input  [63:0] io_mem_cluster_35_data,
  output        io_mem_cluster_36_en,
  output [7:0]  io_mem_cluster_36_addr,
  input  [63:0] io_mem_cluster_36_data,
  output        io_mem_cluster_37_en,
  output [7:0]  io_mem_cluster_37_addr,
  input  [63:0] io_mem_cluster_37_data,
  output        io_mem_cluster_38_en,
  output [7:0]  io_mem_cluster_38_addr,
  input  [63:0] io_mem_cluster_38_data,
  output        io_mem_cluster_39_en,
  output [7:0]  io_mem_cluster_39_addr,
  input  [63:0] io_mem_cluster_39_data,
  output        io_mem_cluster_40_en,
  output [7:0]  io_mem_cluster_40_addr,
  input  [63:0] io_mem_cluster_40_data,
  output        io_mem_cluster_41_en,
  output [7:0]  io_mem_cluster_41_addr,
  input  [63:0] io_mem_cluster_41_data,
  output        io_mem_cluster_42_en,
  output [7:0]  io_mem_cluster_42_addr,
  input  [63:0] io_mem_cluster_42_data,
  output        io_mem_cluster_43_en,
  output [7:0]  io_mem_cluster_43_addr,
  input  [63:0] io_mem_cluster_43_data,
  output        io_mem_cluster_44_en,
  output [7:0]  io_mem_cluster_44_addr,
  input  [63:0] io_mem_cluster_44_data,
  output        io_mem_cluster_45_en,
  output [7:0]  io_mem_cluster_45_addr,
  input  [63:0] io_mem_cluster_45_data,
  output        io_mem_cluster_46_en,
  output [7:0]  io_mem_cluster_46_addr,
  input  [63:0] io_mem_cluster_46_data,
  output        io_mem_cluster_47_en,
  output [7:0]  io_mem_cluster_47_addr,
  input  [63:0] io_mem_cluster_47_data,
  output        io_mem_cluster_48_en,
  output [7:0]  io_mem_cluster_48_addr,
  input  [63:0] io_mem_cluster_48_data,
  output        io_mem_cluster_49_en,
  output [7:0]  io_mem_cluster_49_addr,
  input  [63:0] io_mem_cluster_49_data,
  output        io_mem_cluster_50_en,
  output [7:0]  io_mem_cluster_50_addr,
  input  [63:0] io_mem_cluster_50_data,
  output        io_mem_cluster_51_en,
  output [7:0]  io_mem_cluster_51_addr,
  input  [63:0] io_mem_cluster_51_data,
  output        io_mem_cluster_52_en,
  output [7:0]  io_mem_cluster_52_addr,
  input  [63:0] io_mem_cluster_52_data,
  output        io_mem_cluster_53_en,
  output [7:0]  io_mem_cluster_53_addr,
  input  [63:0] io_mem_cluster_53_data,
  output        io_mem_cluster_54_en,
  output [7:0]  io_mem_cluster_54_addr,
  input  [63:0] io_mem_cluster_54_data,
  output        io_mem_cluster_55_en,
  output [7:0]  io_mem_cluster_55_addr,
  input  [63:0] io_mem_cluster_55_data,
  output        io_mem_cluster_56_en,
  output [7:0]  io_mem_cluster_56_addr,
  input  [63:0] io_mem_cluster_56_data,
  output        io_mem_cluster_57_en,
  output [7:0]  io_mem_cluster_57_addr,
  input  [63:0] io_mem_cluster_57_data,
  output        io_mem_cluster_58_en,
  output [7:0]  io_mem_cluster_58_addr,
  input  [63:0] io_mem_cluster_58_data,
  output        io_mem_cluster_59_en,
  output [7:0]  io_mem_cluster_59_addr,
  input  [63:0] io_mem_cluster_59_data,
  output        io_mem_cluster_60_en,
  output [7:0]  io_mem_cluster_60_addr,
  input  [63:0] io_mem_cluster_60_data,
  output        io_mem_cluster_61_en,
  output [7:0]  io_mem_cluster_61_addr,
  input  [63:0] io_mem_cluster_61_data,
  output        io_mem_cluster_62_en,
  output [7:0]  io_mem_cluster_62_addr,
  input  [63:0] io_mem_cluster_62_data,
  output        io_mem_cluster_63_en,
  output [7:0]  io_mem_cluster_63_addr,
  input  [63:0] io_mem_cluster_63_data
);
  wire  PAR_clock; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_0; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_1; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_2; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_3; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_4; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_5; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_6; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_7; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_8; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_9; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_10; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_11; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_12; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_13; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_14; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_15; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_16; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_17; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_18; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_19; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_20; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_21; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_22; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_23; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_24; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_25; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_26; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_27; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_28; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_29; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_30; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_31; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_32; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_33; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_34; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_35; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_36; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_37; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_38; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_39; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_40; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_41; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_42; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_43; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_44; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_45; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_46; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_47; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_48; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_49; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_50; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_51; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_52; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_53; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_54; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_55; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_56; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_57; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_58; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_59; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_60; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_61; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_62; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_63; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_64; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_65; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_66; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_67; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_68; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_69; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_70; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_71; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_72; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_73; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_74; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_75; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_76; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_77; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_78; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_79; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_80; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_81; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_82; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_83; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_84; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_85; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_86; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_87; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_88; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_89; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_90; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_91; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_92; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_93; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_94; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_95; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_96; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_97; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_98; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_99; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_100; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_101; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_102; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_103; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_104; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_105; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_106; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_107; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_108; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_109; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_110; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_111; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_112; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_113; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_114; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_115; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_116; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_117; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_118; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_119; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_120; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_121; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_122; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_123; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_124; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_125; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_126; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_127; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_128; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_129; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_130; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_131; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_132; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_133; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_134; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_135; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_136; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_137; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_138; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_139; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_140; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_141; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_142; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_143; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_144; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_145; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_146; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_147; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_148; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_149; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_150; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_151; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_152; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_153; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_154; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_155; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_156; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_157; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_158; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_159; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_160; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_161; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_162; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_163; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_164; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_165; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_166; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_167; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_168; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_169; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_170; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_171; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_172; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_173; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_174; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_175; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_176; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_177; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_178; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_179; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_180; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_181; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_182; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_183; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_184; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_185; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_186; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_187; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_188; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_189; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_190; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_191; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_192; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_193; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_194; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_195; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_196; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_197; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_198; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_199; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_200; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_201; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_202; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_203; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_204; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_205; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_206; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_207; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_208; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_209; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_210; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_211; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_212; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_213; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_214; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_215; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_216; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_217; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_218; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_219; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_220; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_221; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_222; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_223; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_224; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_225; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_226; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_227; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_228; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_229; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_230; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_231; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_232; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_233; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_234; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_235; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_236; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_237; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_238; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_239; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_240; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_241; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_242; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_243; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_244; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_245; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_246; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_247; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_248; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_249; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_250; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_251; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_252; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_253; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_254; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_255; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_0; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_1; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_2; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_3; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_4; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_5; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_6; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_7; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_8; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_9; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_10; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_11; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_12; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_13; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_14; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_15; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_parse_current_state; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_parse_current_offset; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_parse_transition_field; // @[processor.scala 13:21]
  wire [2:0] PAR_io_pipe_phv_in_next_processor_id; // @[processor.scala 13:21]
  wire  PAR_io_pipe_phv_in_next_config_id; // @[processor.scala 13:21]
  wire  PAR_io_pipe_phv_in_is_valid_processor; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_0; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_1; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_2; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_3; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_4; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_5; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_6; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_7; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_8; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_9; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_10; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_11; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_12; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_13; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_14; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_15; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_16; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_17; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_18; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_19; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_20; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_21; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_22; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_23; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_24; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_25; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_26; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_27; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_28; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_29; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_30; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_31; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_32; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_33; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_34; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_35; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_36; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_37; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_38; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_39; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_40; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_41; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_42; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_43; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_44; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_45; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_46; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_47; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_48; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_49; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_50; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_51; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_52; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_53; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_54; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_55; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_56; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_57; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_58; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_59; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_60; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_61; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_62; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_63; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_64; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_65; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_66; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_67; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_68; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_69; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_70; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_71; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_72; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_73; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_74; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_75; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_76; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_77; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_78; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_79; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_80; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_81; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_82; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_83; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_84; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_85; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_86; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_87; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_88; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_89; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_90; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_91; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_92; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_93; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_94; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_95; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_96; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_97; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_98; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_99; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_100; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_101; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_102; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_103; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_104; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_105; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_106; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_107; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_108; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_109; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_110; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_111; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_112; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_113; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_114; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_115; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_116; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_117; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_118; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_119; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_120; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_121; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_122; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_123; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_124; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_125; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_126; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_127; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_128; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_129; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_130; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_131; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_132; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_133; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_134; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_135; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_136; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_137; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_138; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_139; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_140; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_141; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_142; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_143; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_144; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_145; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_146; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_147; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_148; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_149; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_150; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_151; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_152; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_153; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_154; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_155; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_156; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_157; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_158; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_159; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_160; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_161; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_162; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_163; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_164; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_165; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_166; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_167; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_168; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_169; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_170; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_171; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_172; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_173; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_174; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_175; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_176; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_177; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_178; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_179; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_180; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_181; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_182; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_183; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_184; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_185; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_186; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_187; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_188; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_189; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_190; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_191; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_192; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_193; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_194; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_195; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_196; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_197; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_198; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_199; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_200; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_201; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_202; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_203; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_204; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_205; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_206; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_207; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_208; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_209; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_210; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_211; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_212; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_213; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_214; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_215; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_216; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_217; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_218; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_219; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_220; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_221; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_222; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_223; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_224; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_225; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_226; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_227; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_228; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_229; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_230; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_231; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_232; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_233; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_234; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_235; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_236; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_237; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_238; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_239; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_240; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_241; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_242; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_243; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_244; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_245; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_246; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_247; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_248; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_249; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_250; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_251; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_252; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_253; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_254; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_255; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_0; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_1; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_2; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_3; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_4; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_5; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_6; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_7; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_8; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_9; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_10; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_11; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_12; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_13; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_14; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_15; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_parse_current_state; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_parse_current_offset; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_parse_transition_field; // @[processor.scala 13:21]
  wire [2:0] PAR_io_pipe_phv_out_next_processor_id; // @[processor.scala 13:21]
  wire  PAR_io_pipe_phv_out_next_config_id; // @[processor.scala 13:21]
  wire  PAR_io_pipe_phv_out_is_valid_processor; // @[processor.scala 13:21]
  wire  PAR_io_mod_en; // @[processor.scala 13:21]
  wire  PAR_io_mod_last_mau_id_mod; // @[processor.scala 13:21]
  wire [1:0] PAR_io_mod_last_mau_id; // @[processor.scala 13:21]
  wire [1:0] PAR_io_mod_cs; // @[processor.scala 13:21]
  wire  PAR_io_mod_module_mod_state_id_mod; // @[processor.scala 13:21]
  wire [7:0] PAR_io_mod_module_mod_state_id; // @[processor.scala 13:21]
  wire  PAR_io_mod_module_mod_sram_w_cs; // @[processor.scala 13:21]
  wire  PAR_io_mod_module_mod_sram_w_en; // @[processor.scala 13:21]
  wire [7:0] PAR_io_mod_module_mod_sram_w_addr; // @[processor.scala 13:21]
  wire [63:0] PAR_io_mod_module_mod_sram_w_data; // @[processor.scala 13:21]
  wire  MAT_clock; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_0; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_1; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_2; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_3; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_4; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_5; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_6; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_7; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_8; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_9; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_10; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_11; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_12; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_13; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_14; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_15; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_16; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_17; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_18; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_19; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_20; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_21; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_22; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_23; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_24; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_25; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_26; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_27; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_28; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_29; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_30; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_31; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_32; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_33; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_34; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_35; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_36; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_37; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_38; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_39; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_40; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_41; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_42; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_43; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_44; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_45; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_46; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_47; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_48; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_49; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_50; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_51; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_52; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_53; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_54; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_55; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_56; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_57; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_58; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_59; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_60; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_61; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_62; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_63; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_64; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_65; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_66; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_67; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_68; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_69; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_70; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_71; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_72; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_73; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_74; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_75; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_76; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_77; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_78; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_79; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_80; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_81; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_82; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_83; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_84; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_85; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_86; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_87; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_88; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_89; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_90; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_91; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_92; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_93; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_94; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_95; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_96; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_97; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_98; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_99; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_100; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_101; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_102; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_103; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_104; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_105; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_106; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_107; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_108; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_109; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_110; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_111; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_112; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_113; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_114; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_115; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_116; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_117; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_118; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_119; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_120; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_121; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_122; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_123; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_124; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_125; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_126; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_127; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_128; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_129; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_130; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_131; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_132; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_133; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_134; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_135; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_136; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_137; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_138; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_139; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_140; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_141; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_142; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_143; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_144; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_145; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_146; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_147; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_148; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_149; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_150; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_151; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_152; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_153; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_154; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_155; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_156; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_157; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_158; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_159; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_160; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_161; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_162; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_163; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_164; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_165; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_166; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_167; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_168; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_169; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_170; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_171; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_172; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_173; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_174; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_175; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_176; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_177; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_178; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_179; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_180; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_181; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_182; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_183; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_184; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_185; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_186; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_187; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_188; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_189; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_190; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_191; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_192; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_193; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_194; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_195; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_196; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_197; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_198; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_199; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_200; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_201; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_202; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_203; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_204; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_205; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_206; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_207; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_208; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_209; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_210; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_211; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_212; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_213; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_214; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_215; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_216; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_217; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_218; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_219; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_220; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_221; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_222; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_223; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_224; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_225; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_226; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_227; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_228; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_229; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_230; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_231; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_232; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_233; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_234; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_235; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_236; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_237; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_238; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_239; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_240; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_241; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_242; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_243; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_244; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_245; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_246; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_247; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_248; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_249; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_250; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_251; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_252; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_253; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_254; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_255; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_0; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_1; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_2; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_3; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_4; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_5; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_6; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_7; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_8; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_9; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_10; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_11; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_12; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_13; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_14; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_15; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_parse_current_state; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_parse_current_offset; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_parse_transition_field; // @[processor.scala 14:21]
  wire [2:0] MAT_io_pipe_phv_in_next_processor_id; // @[processor.scala 14:21]
  wire  MAT_io_pipe_phv_in_next_config_id; // @[processor.scala 14:21]
  wire  MAT_io_pipe_phv_in_is_valid_processor; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_0; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_1; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_2; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_3; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_4; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_5; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_6; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_7; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_8; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_9; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_10; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_11; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_12; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_13; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_14; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_15; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_16; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_17; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_18; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_19; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_20; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_21; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_22; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_23; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_24; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_25; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_26; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_27; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_28; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_29; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_30; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_31; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_32; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_33; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_34; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_35; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_36; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_37; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_38; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_39; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_40; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_41; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_42; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_43; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_44; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_45; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_46; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_47; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_48; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_49; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_50; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_51; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_52; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_53; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_54; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_55; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_56; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_57; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_58; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_59; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_60; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_61; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_62; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_63; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_64; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_65; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_66; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_67; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_68; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_69; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_70; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_71; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_72; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_73; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_74; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_75; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_76; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_77; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_78; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_79; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_80; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_81; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_82; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_83; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_84; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_85; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_86; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_87; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_88; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_89; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_90; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_91; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_92; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_93; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_94; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_95; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_96; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_97; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_98; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_99; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_100; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_101; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_102; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_103; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_104; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_105; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_106; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_107; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_108; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_109; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_110; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_111; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_112; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_113; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_114; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_115; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_116; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_117; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_118; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_119; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_120; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_121; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_122; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_123; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_124; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_125; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_126; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_127; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_128; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_129; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_130; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_131; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_132; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_133; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_134; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_135; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_136; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_137; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_138; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_139; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_140; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_141; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_142; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_143; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_144; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_145; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_146; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_147; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_148; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_149; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_150; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_151; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_152; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_153; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_154; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_155; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_156; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_157; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_158; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_159; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_160; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_161; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_162; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_163; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_164; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_165; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_166; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_167; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_168; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_169; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_170; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_171; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_172; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_173; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_174; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_175; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_176; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_177; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_178; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_179; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_180; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_181; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_182; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_183; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_184; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_185; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_186; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_187; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_188; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_189; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_190; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_191; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_192; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_193; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_194; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_195; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_196; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_197; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_198; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_199; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_200; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_201; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_202; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_203; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_204; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_205; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_206; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_207; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_208; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_209; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_210; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_211; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_212; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_213; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_214; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_215; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_216; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_217; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_218; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_219; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_220; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_221; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_222; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_223; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_224; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_225; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_226; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_227; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_228; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_229; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_230; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_231; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_232; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_233; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_234; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_235; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_236; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_237; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_238; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_239; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_240; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_241; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_242; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_243; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_244; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_245; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_246; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_247; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_248; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_249; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_250; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_251; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_252; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_253; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_254; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_255; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_0; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_1; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_2; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_3; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_4; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_5; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_6; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_7; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_8; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_9; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_10; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_11; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_12; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_13; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_14; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_15; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_parse_current_state; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_parse_current_offset; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_parse_transition_field; // @[processor.scala 14:21]
  wire [2:0] MAT_io_pipe_phv_out_next_processor_id; // @[processor.scala 14:21]
  wire  MAT_io_pipe_phv_out_next_config_id; // @[processor.scala 14:21]
  wire  MAT_io_pipe_phv_out_is_valid_processor; // @[processor.scala 14:21]
  wire  MAT_io_mod_en; // @[processor.scala 14:21]
  wire  MAT_io_mod_config_id; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mod_key_mod_header_id; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mod_key_mod_internal_offset; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mod_key_mod_key_length; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_0; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_1; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_2; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_3; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_4; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_5; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_6; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_7; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_8; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_9; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_10; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_11; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_12; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_13; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_14; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_15; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_16; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_17; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_18; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_19; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_20; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_21; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_22; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_23; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_24; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_25; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_26; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_27; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_28; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_29; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_30; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_31; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_32; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_33; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_34; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_35; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_36; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_37; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_38; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_39; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_40; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_41; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_42; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_43; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_44; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_45; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_46; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_47; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_48; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_49; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_50; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_51; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_52; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_53; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_54; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_55; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_56; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_57; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_58; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_59; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_60; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_61; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_62; // @[processor.scala 14:21]
  wire [5:0] MAT_io_mod_table_mod_sram_id_table_63; // @[processor.scala 14:21]
  wire [6:0] MAT_io_mod_table_mod_table_width; // @[processor.scala 14:21]
  wire [6:0] MAT_io_mod_table_mod_table_depth; // @[processor.scala 14:21]
  wire  MAT_io_hit; // @[processor.scala 14:21]
  wire [63:0] MAT_io_match_value; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_0_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_0_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_0_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_1_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_1_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_1_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_2_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_2_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_2_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_3_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_3_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_3_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_4_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_4_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_4_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_5_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_5_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_5_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_6_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_6_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_6_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_7_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_7_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_7_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_8_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_8_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_8_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_9_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_9_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_9_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_10_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_10_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_10_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_11_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_11_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_11_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_12_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_12_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_12_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_13_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_13_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_13_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_14_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_14_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_14_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_15_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_15_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_15_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_16_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_16_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_16_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_17_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_17_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_17_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_18_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_18_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_18_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_19_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_19_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_19_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_20_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_20_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_20_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_21_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_21_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_21_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_22_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_22_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_22_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_23_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_23_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_23_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_24_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_24_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_24_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_25_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_25_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_25_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_26_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_26_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_26_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_27_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_27_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_27_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_28_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_28_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_28_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_29_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_29_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_29_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_30_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_30_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_30_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_31_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_31_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_31_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_32_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_32_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_32_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_33_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_33_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_33_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_34_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_34_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_34_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_35_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_35_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_35_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_36_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_36_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_36_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_37_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_37_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_37_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_38_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_38_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_38_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_39_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_39_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_39_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_40_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_40_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_40_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_41_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_41_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_41_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_42_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_42_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_42_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_43_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_43_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_43_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_44_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_44_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_44_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_45_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_45_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_45_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_46_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_46_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_46_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_47_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_47_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_47_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_48_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_48_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_48_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_49_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_49_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_49_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_50_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_50_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_50_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_51_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_51_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_51_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_52_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_52_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_52_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_53_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_53_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_53_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_54_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_54_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_54_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_55_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_55_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_55_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_56_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_56_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_56_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_57_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_57_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_57_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_58_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_58_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_58_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_59_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_59_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_59_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_60_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_60_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_60_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_61_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_61_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_61_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_62_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_62_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_62_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_63_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_63_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_63_data; // @[processor.scala 14:21]
  wire  EXE_clock; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_0; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_1; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_2; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_3; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_4; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_5; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_6; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_7; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_8; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_9; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_10; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_11; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_12; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_13; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_14; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_15; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_16; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_17; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_18; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_19; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_20; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_21; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_22; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_23; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_24; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_25; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_26; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_27; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_28; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_29; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_30; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_31; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_32; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_33; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_34; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_35; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_36; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_37; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_38; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_39; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_40; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_41; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_42; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_43; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_44; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_45; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_46; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_47; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_48; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_49; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_50; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_51; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_52; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_53; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_54; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_55; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_56; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_57; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_58; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_59; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_60; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_61; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_62; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_63; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_64; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_65; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_66; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_67; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_68; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_69; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_70; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_71; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_72; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_73; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_74; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_75; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_76; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_77; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_78; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_79; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_80; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_81; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_82; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_83; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_84; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_85; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_86; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_87; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_88; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_89; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_90; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_91; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_92; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_93; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_94; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_95; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_96; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_97; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_98; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_99; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_100; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_101; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_102; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_103; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_104; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_105; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_106; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_107; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_108; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_109; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_110; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_111; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_112; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_113; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_114; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_115; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_116; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_117; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_118; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_119; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_120; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_121; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_122; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_123; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_124; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_125; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_126; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_127; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_128; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_129; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_130; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_131; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_132; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_133; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_134; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_135; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_136; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_137; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_138; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_139; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_140; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_141; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_142; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_143; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_144; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_145; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_146; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_147; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_148; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_149; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_150; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_151; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_152; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_153; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_154; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_155; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_156; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_157; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_158; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_159; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_160; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_161; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_162; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_163; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_164; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_165; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_166; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_167; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_168; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_169; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_170; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_171; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_172; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_173; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_174; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_175; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_176; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_177; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_178; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_179; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_180; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_181; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_182; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_183; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_184; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_185; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_186; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_187; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_188; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_189; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_190; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_191; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_192; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_193; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_194; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_195; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_196; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_197; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_198; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_199; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_200; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_201; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_202; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_203; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_204; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_205; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_206; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_207; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_208; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_209; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_210; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_211; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_212; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_213; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_214; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_215; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_216; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_217; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_218; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_219; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_220; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_221; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_222; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_223; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_224; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_225; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_226; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_227; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_228; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_229; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_230; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_231; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_232; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_233; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_234; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_235; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_236; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_237; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_238; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_239; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_240; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_241; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_242; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_243; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_244; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_245; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_246; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_247; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_248; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_249; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_250; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_251; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_252; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_253; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_254; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_255; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_0; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_1; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_2; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_3; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_4; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_5; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_6; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_7; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_8; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_9; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_10; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_11; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_12; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_13; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_14; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_15; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_parse_current_state; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_parse_current_offset; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_parse_transition_field; // @[processor.scala 15:21]
  wire [2:0] EXE_io_pipe_phv_in_next_processor_id; // @[processor.scala 15:21]
  wire  EXE_io_pipe_phv_in_next_config_id; // @[processor.scala 15:21]
  wire  EXE_io_pipe_phv_in_is_valid_processor; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_0; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_1; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_2; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_3; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_4; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_5; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_6; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_7; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_8; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_9; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_10; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_11; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_12; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_13; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_14; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_15; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_16; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_17; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_18; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_19; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_20; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_21; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_22; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_23; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_24; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_25; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_26; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_27; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_28; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_29; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_30; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_31; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_32; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_33; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_34; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_35; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_36; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_37; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_38; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_39; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_40; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_41; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_42; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_43; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_44; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_45; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_46; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_47; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_48; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_49; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_50; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_51; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_52; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_53; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_54; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_55; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_56; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_57; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_58; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_59; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_60; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_61; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_62; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_63; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_64; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_65; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_66; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_67; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_68; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_69; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_70; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_71; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_72; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_73; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_74; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_75; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_76; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_77; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_78; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_79; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_80; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_81; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_82; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_83; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_84; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_85; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_86; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_87; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_88; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_89; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_90; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_91; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_92; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_93; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_94; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_95; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_96; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_97; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_98; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_99; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_100; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_101; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_102; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_103; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_104; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_105; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_106; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_107; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_108; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_109; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_110; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_111; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_112; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_113; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_114; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_115; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_116; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_117; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_118; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_119; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_120; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_121; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_122; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_123; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_124; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_125; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_126; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_127; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_128; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_129; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_130; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_131; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_132; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_133; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_134; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_135; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_136; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_137; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_138; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_139; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_140; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_141; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_142; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_143; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_144; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_145; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_146; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_147; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_148; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_149; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_150; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_151; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_152; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_153; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_154; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_155; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_156; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_157; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_158; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_159; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_160; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_161; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_162; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_163; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_164; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_165; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_166; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_167; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_168; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_169; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_170; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_171; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_172; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_173; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_174; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_175; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_176; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_177; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_178; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_179; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_180; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_181; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_182; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_183; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_184; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_185; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_186; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_187; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_188; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_189; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_190; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_191; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_192; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_193; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_194; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_195; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_196; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_197; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_198; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_199; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_200; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_201; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_202; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_203; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_204; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_205; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_206; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_207; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_208; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_209; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_210; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_211; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_212; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_213; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_214; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_215; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_216; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_217; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_218; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_219; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_220; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_221; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_222; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_223; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_224; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_225; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_226; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_227; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_228; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_229; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_230; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_231; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_232; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_233; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_234; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_235; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_236; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_237; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_238; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_239; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_240; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_241; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_242; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_243; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_244; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_245; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_246; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_247; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_248; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_249; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_250; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_251; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_252; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_253; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_254; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_255; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_0; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_1; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_2; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_3; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_4; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_5; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_6; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_7; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_8; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_9; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_10; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_11; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_12; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_13; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_14; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_15; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_parse_current_state; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_parse_current_offset; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_parse_transition_field; // @[processor.scala 15:21]
  wire [2:0] EXE_io_pipe_phv_out_next_processor_id; // @[processor.scala 15:21]
  wire  EXE_io_pipe_phv_out_next_config_id; // @[processor.scala 15:21]
  wire  EXE_io_hit; // @[processor.scala 15:21]
  wire [63:0] EXE_io_match_value; // @[processor.scala 15:21]
  wire  EXE_io_action_mod_en_0; // @[processor.scala 15:21]
  wire  EXE_io_action_mod_en_1; // @[processor.scala 15:21]
  wire [7:0] EXE_io_action_mod_addr; // @[processor.scala 15:21]
  wire [63:0] EXE_io_action_mod_data_0; // @[processor.scala 15:21]
  wire [63:0] EXE_io_action_mod_data_1; // @[processor.scala 15:21]
  Parser PAR ( // @[processor.scala 13:21]
    .clock(PAR_clock),
    .io_pipe_phv_in_data_0(PAR_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(PAR_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(PAR_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(PAR_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(PAR_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(PAR_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(PAR_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(PAR_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(PAR_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(PAR_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(PAR_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(PAR_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(PAR_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(PAR_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(PAR_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(PAR_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(PAR_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(PAR_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(PAR_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(PAR_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(PAR_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(PAR_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(PAR_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(PAR_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(PAR_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(PAR_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(PAR_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(PAR_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(PAR_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(PAR_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(PAR_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(PAR_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(PAR_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(PAR_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(PAR_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(PAR_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(PAR_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(PAR_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(PAR_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(PAR_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(PAR_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(PAR_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(PAR_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(PAR_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(PAR_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(PAR_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(PAR_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(PAR_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(PAR_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(PAR_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(PAR_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(PAR_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(PAR_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(PAR_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(PAR_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(PAR_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(PAR_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(PAR_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(PAR_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(PAR_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(PAR_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(PAR_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(PAR_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(PAR_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(PAR_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(PAR_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(PAR_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(PAR_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(PAR_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(PAR_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(PAR_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(PAR_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(PAR_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(PAR_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(PAR_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(PAR_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(PAR_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(PAR_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(PAR_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(PAR_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(PAR_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(PAR_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(PAR_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(PAR_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(PAR_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(PAR_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(PAR_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(PAR_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(PAR_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(PAR_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(PAR_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(PAR_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(PAR_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(PAR_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(PAR_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(PAR_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(PAR_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(PAR_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(PAR_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(PAR_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(PAR_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(PAR_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(PAR_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(PAR_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(PAR_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(PAR_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(PAR_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(PAR_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(PAR_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(PAR_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(PAR_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(PAR_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(PAR_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(PAR_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(PAR_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(PAR_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(PAR_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(PAR_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(PAR_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(PAR_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(PAR_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(PAR_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(PAR_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(PAR_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(PAR_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(PAR_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(PAR_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(PAR_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(PAR_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(PAR_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(PAR_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(PAR_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(PAR_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(PAR_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(PAR_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(PAR_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(PAR_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(PAR_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(PAR_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(PAR_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(PAR_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(PAR_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(PAR_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(PAR_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(PAR_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(PAR_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(PAR_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(PAR_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(PAR_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(PAR_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(PAR_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(PAR_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(PAR_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(PAR_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(PAR_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(PAR_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(PAR_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(PAR_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(PAR_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(PAR_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(PAR_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(PAR_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(PAR_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(PAR_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(PAR_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(PAR_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(PAR_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(PAR_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(PAR_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(PAR_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(PAR_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(PAR_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(PAR_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(PAR_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(PAR_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(PAR_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(PAR_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(PAR_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(PAR_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(PAR_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(PAR_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(PAR_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(PAR_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(PAR_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(PAR_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(PAR_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(PAR_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(PAR_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(PAR_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(PAR_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(PAR_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(PAR_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(PAR_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(PAR_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(PAR_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(PAR_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(PAR_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(PAR_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(PAR_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(PAR_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(PAR_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(PAR_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(PAR_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(PAR_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(PAR_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(PAR_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(PAR_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(PAR_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(PAR_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(PAR_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(PAR_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(PAR_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(PAR_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(PAR_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(PAR_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(PAR_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(PAR_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(PAR_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(PAR_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(PAR_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(PAR_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(PAR_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(PAR_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(PAR_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(PAR_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(PAR_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(PAR_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(PAR_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(PAR_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(PAR_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(PAR_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(PAR_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(PAR_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(PAR_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(PAR_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(PAR_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(PAR_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(PAR_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(PAR_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(PAR_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(PAR_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(PAR_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(PAR_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(PAR_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(PAR_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(PAR_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(PAR_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(PAR_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(PAR_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(PAR_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(PAR_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(PAR_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(PAR_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(PAR_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(PAR_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(PAR_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(PAR_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(PAR_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(PAR_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(PAR_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(PAR_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(PAR_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(PAR_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(PAR_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(PAR_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(PAR_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(PAR_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(PAR_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(PAR_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(PAR_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(PAR_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(PAR_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(PAR_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(PAR_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(PAR_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(PAR_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(PAR_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(PAR_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(PAR_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(PAR_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(PAR_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(PAR_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(PAR_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(PAR_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(PAR_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(PAR_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(PAR_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(PAR_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(PAR_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(PAR_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(PAR_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(PAR_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(PAR_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(PAR_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(PAR_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(PAR_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(PAR_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(PAR_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(PAR_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(PAR_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(PAR_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(PAR_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(PAR_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(PAR_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(PAR_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(PAR_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(PAR_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(PAR_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(PAR_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(PAR_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(PAR_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(PAR_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(PAR_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(PAR_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(PAR_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(PAR_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(PAR_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(PAR_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(PAR_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(PAR_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(PAR_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(PAR_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(PAR_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(PAR_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(PAR_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(PAR_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(PAR_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(PAR_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(PAR_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(PAR_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(PAR_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(PAR_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(PAR_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(PAR_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(PAR_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(PAR_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(PAR_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(PAR_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(PAR_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(PAR_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(PAR_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(PAR_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(PAR_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(PAR_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(PAR_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(PAR_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(PAR_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(PAR_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(PAR_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(PAR_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(PAR_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(PAR_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(PAR_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(PAR_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(PAR_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(PAR_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(PAR_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(PAR_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(PAR_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(PAR_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(PAR_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(PAR_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(PAR_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(PAR_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(PAR_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(PAR_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(PAR_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(PAR_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(PAR_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(PAR_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(PAR_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(PAR_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(PAR_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(PAR_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(PAR_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(PAR_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(PAR_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(PAR_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(PAR_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(PAR_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(PAR_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(PAR_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(PAR_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(PAR_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(PAR_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(PAR_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(PAR_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(PAR_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(PAR_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(PAR_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(PAR_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(PAR_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(PAR_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(PAR_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(PAR_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(PAR_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(PAR_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(PAR_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(PAR_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(PAR_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(PAR_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(PAR_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(PAR_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(PAR_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(PAR_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(PAR_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(PAR_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(PAR_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(PAR_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(PAR_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(PAR_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(PAR_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(PAR_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(PAR_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(PAR_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(PAR_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(PAR_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(PAR_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(PAR_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(PAR_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(PAR_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(PAR_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(PAR_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(PAR_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(PAR_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(PAR_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(PAR_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(PAR_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(PAR_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(PAR_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(PAR_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(PAR_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(PAR_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(PAR_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(PAR_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(PAR_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(PAR_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(PAR_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(PAR_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(PAR_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(PAR_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(PAR_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(PAR_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(PAR_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(PAR_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(PAR_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(PAR_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(PAR_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(PAR_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(PAR_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(PAR_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(PAR_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(PAR_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(PAR_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(PAR_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(PAR_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(PAR_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(PAR_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(PAR_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(PAR_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(PAR_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(PAR_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(PAR_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(PAR_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(PAR_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(PAR_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(PAR_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(PAR_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(PAR_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(PAR_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(PAR_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(PAR_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(PAR_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(PAR_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(PAR_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(PAR_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(PAR_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(PAR_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(PAR_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(PAR_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(PAR_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(PAR_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(PAR_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(PAR_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(PAR_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(PAR_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(PAR_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(PAR_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(PAR_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(PAR_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(PAR_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(PAR_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(PAR_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(PAR_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(PAR_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(PAR_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(PAR_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(PAR_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(PAR_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(PAR_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(PAR_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(PAR_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(PAR_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(PAR_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(PAR_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(PAR_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(PAR_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(PAR_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(PAR_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(PAR_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(PAR_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(PAR_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(PAR_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(PAR_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(PAR_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(PAR_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(PAR_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(PAR_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(PAR_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(PAR_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(PAR_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(PAR_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(PAR_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(PAR_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(PAR_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(PAR_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(PAR_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(PAR_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(PAR_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(PAR_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(PAR_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(PAR_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(PAR_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(PAR_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(PAR_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(PAR_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(PAR_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(PAR_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(PAR_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(PAR_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(PAR_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(PAR_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(PAR_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(PAR_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(PAR_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(PAR_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(PAR_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(PAR_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(PAR_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(PAR_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(PAR_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(PAR_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(PAR_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(PAR_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(PAR_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(PAR_io_pipe_phv_out_is_valid_processor),
    .io_mod_en(PAR_io_mod_en),
    .io_mod_last_mau_id_mod(PAR_io_mod_last_mau_id_mod),
    .io_mod_last_mau_id(PAR_io_mod_last_mau_id),
    .io_mod_cs(PAR_io_mod_cs),
    .io_mod_module_mod_state_id_mod(PAR_io_mod_module_mod_state_id_mod),
    .io_mod_module_mod_state_id(PAR_io_mod_module_mod_state_id),
    .io_mod_module_mod_sram_w_cs(PAR_io_mod_module_mod_sram_w_cs),
    .io_mod_module_mod_sram_w_en(PAR_io_mod_module_mod_sram_w_en),
    .io_mod_module_mod_sram_w_addr(PAR_io_mod_module_mod_sram_w_addr),
    .io_mod_module_mod_sram_w_data(PAR_io_mod_module_mod_sram_w_data)
  );
  Matcher MAT ( // @[processor.scala 14:21]
    .clock(MAT_clock),
    .io_pipe_phv_in_data_0(MAT_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(MAT_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(MAT_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(MAT_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(MAT_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(MAT_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(MAT_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(MAT_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(MAT_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(MAT_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(MAT_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(MAT_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(MAT_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(MAT_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(MAT_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(MAT_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(MAT_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(MAT_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(MAT_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(MAT_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(MAT_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(MAT_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(MAT_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(MAT_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(MAT_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(MAT_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(MAT_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(MAT_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(MAT_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(MAT_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(MAT_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(MAT_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(MAT_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(MAT_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(MAT_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(MAT_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(MAT_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(MAT_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(MAT_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(MAT_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(MAT_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(MAT_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(MAT_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(MAT_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(MAT_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(MAT_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(MAT_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(MAT_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(MAT_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(MAT_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(MAT_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(MAT_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(MAT_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(MAT_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(MAT_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(MAT_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(MAT_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(MAT_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(MAT_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(MAT_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(MAT_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(MAT_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(MAT_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(MAT_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(MAT_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(MAT_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(MAT_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(MAT_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(MAT_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(MAT_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(MAT_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(MAT_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(MAT_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(MAT_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(MAT_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(MAT_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(MAT_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(MAT_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(MAT_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(MAT_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(MAT_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(MAT_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(MAT_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(MAT_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(MAT_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(MAT_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(MAT_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(MAT_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(MAT_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(MAT_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(MAT_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(MAT_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(MAT_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(MAT_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(MAT_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(MAT_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(MAT_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(MAT_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(MAT_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(MAT_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(MAT_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(MAT_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(MAT_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(MAT_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(MAT_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(MAT_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(MAT_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(MAT_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(MAT_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(MAT_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(MAT_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(MAT_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(MAT_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(MAT_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(MAT_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(MAT_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(MAT_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(MAT_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(MAT_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(MAT_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(MAT_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(MAT_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(MAT_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(MAT_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(MAT_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(MAT_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(MAT_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(MAT_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(MAT_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(MAT_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(MAT_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(MAT_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(MAT_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(MAT_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(MAT_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(MAT_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(MAT_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(MAT_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(MAT_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(MAT_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(MAT_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(MAT_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(MAT_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(MAT_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(MAT_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(MAT_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(MAT_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(MAT_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(MAT_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(MAT_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(MAT_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(MAT_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(MAT_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(MAT_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(MAT_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(MAT_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(MAT_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(MAT_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(MAT_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(MAT_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(MAT_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(MAT_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(MAT_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(MAT_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(MAT_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(MAT_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(MAT_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(MAT_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(MAT_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(MAT_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(MAT_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(MAT_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(MAT_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(MAT_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(MAT_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(MAT_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(MAT_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(MAT_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(MAT_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(MAT_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(MAT_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(MAT_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(MAT_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(MAT_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(MAT_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(MAT_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(MAT_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(MAT_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(MAT_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(MAT_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(MAT_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(MAT_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(MAT_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(MAT_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(MAT_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(MAT_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(MAT_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(MAT_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(MAT_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(MAT_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(MAT_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(MAT_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(MAT_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(MAT_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(MAT_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(MAT_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(MAT_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(MAT_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(MAT_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(MAT_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(MAT_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(MAT_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(MAT_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(MAT_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(MAT_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(MAT_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(MAT_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(MAT_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(MAT_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(MAT_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(MAT_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(MAT_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(MAT_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(MAT_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(MAT_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(MAT_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(MAT_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(MAT_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(MAT_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(MAT_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(MAT_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(MAT_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(MAT_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(MAT_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(MAT_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(MAT_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(MAT_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(MAT_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(MAT_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(MAT_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(MAT_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(MAT_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(MAT_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(MAT_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(MAT_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(MAT_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(MAT_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(MAT_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(MAT_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(MAT_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(MAT_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(MAT_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(MAT_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(MAT_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(MAT_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(MAT_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(MAT_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(MAT_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(MAT_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(MAT_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(MAT_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(MAT_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(MAT_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(MAT_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(MAT_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(MAT_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(MAT_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(MAT_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(MAT_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(MAT_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(MAT_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(MAT_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(MAT_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(MAT_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(MAT_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(MAT_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(MAT_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(MAT_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(MAT_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(MAT_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(MAT_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(MAT_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(MAT_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(MAT_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(MAT_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(MAT_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(MAT_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(MAT_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(MAT_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(MAT_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(MAT_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(MAT_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(MAT_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(MAT_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(MAT_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(MAT_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(MAT_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(MAT_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(MAT_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(MAT_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(MAT_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(MAT_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(MAT_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(MAT_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(MAT_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(MAT_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(MAT_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(MAT_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(MAT_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(MAT_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(MAT_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(MAT_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(MAT_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(MAT_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(MAT_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(MAT_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(MAT_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(MAT_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(MAT_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(MAT_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(MAT_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(MAT_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(MAT_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(MAT_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(MAT_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(MAT_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(MAT_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(MAT_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(MAT_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(MAT_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(MAT_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(MAT_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(MAT_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(MAT_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(MAT_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(MAT_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(MAT_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(MAT_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(MAT_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(MAT_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(MAT_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(MAT_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(MAT_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(MAT_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(MAT_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(MAT_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(MAT_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(MAT_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(MAT_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(MAT_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(MAT_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(MAT_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(MAT_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(MAT_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(MAT_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(MAT_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(MAT_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(MAT_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(MAT_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(MAT_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(MAT_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(MAT_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(MAT_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(MAT_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(MAT_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(MAT_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(MAT_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(MAT_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(MAT_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(MAT_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(MAT_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(MAT_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(MAT_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(MAT_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(MAT_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(MAT_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(MAT_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(MAT_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(MAT_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(MAT_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(MAT_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(MAT_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(MAT_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(MAT_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(MAT_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(MAT_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(MAT_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(MAT_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(MAT_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(MAT_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(MAT_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(MAT_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(MAT_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(MAT_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(MAT_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(MAT_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(MAT_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(MAT_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(MAT_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(MAT_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(MAT_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(MAT_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(MAT_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(MAT_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(MAT_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(MAT_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(MAT_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(MAT_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(MAT_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(MAT_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(MAT_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(MAT_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(MAT_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(MAT_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(MAT_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(MAT_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(MAT_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(MAT_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(MAT_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(MAT_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(MAT_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(MAT_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(MAT_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(MAT_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(MAT_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(MAT_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(MAT_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(MAT_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(MAT_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(MAT_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(MAT_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(MAT_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(MAT_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(MAT_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(MAT_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(MAT_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(MAT_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(MAT_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(MAT_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(MAT_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(MAT_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(MAT_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(MAT_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(MAT_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(MAT_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(MAT_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(MAT_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(MAT_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(MAT_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(MAT_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(MAT_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(MAT_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(MAT_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(MAT_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(MAT_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(MAT_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(MAT_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(MAT_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(MAT_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(MAT_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(MAT_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(MAT_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(MAT_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(MAT_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(MAT_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(MAT_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(MAT_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(MAT_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(MAT_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(MAT_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(MAT_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(MAT_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(MAT_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(MAT_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(MAT_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(MAT_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(MAT_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(MAT_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(MAT_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(MAT_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(MAT_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(MAT_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(MAT_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(MAT_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(MAT_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(MAT_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(MAT_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(MAT_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(MAT_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(MAT_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(MAT_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(MAT_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(MAT_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(MAT_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(MAT_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(MAT_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(MAT_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(MAT_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(MAT_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(MAT_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(MAT_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(MAT_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(MAT_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(MAT_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(MAT_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(MAT_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(MAT_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(MAT_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(MAT_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(MAT_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(MAT_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(MAT_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(MAT_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(MAT_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(MAT_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(MAT_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(MAT_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(MAT_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(MAT_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(MAT_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(MAT_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(MAT_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(MAT_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(MAT_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(MAT_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(MAT_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(MAT_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(MAT_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(MAT_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(MAT_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(MAT_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(MAT_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(MAT_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(MAT_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(MAT_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(MAT_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(MAT_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(MAT_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(MAT_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(MAT_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(MAT_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(MAT_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(MAT_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(MAT_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(MAT_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(MAT_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(MAT_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(MAT_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(MAT_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(MAT_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(MAT_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(MAT_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(MAT_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(MAT_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(MAT_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(MAT_io_pipe_phv_out_is_valid_processor),
    .io_mod_en(MAT_io_mod_en),
    .io_mod_config_id(MAT_io_mod_config_id),
    .io_mod_key_mod_header_id(MAT_io_mod_key_mod_header_id),
    .io_mod_key_mod_internal_offset(MAT_io_mod_key_mod_internal_offset),
    .io_mod_key_mod_key_length(MAT_io_mod_key_mod_key_length),
    .io_mod_table_mod_sram_id_table_0(MAT_io_mod_table_mod_sram_id_table_0),
    .io_mod_table_mod_sram_id_table_1(MAT_io_mod_table_mod_sram_id_table_1),
    .io_mod_table_mod_sram_id_table_2(MAT_io_mod_table_mod_sram_id_table_2),
    .io_mod_table_mod_sram_id_table_3(MAT_io_mod_table_mod_sram_id_table_3),
    .io_mod_table_mod_sram_id_table_4(MAT_io_mod_table_mod_sram_id_table_4),
    .io_mod_table_mod_sram_id_table_5(MAT_io_mod_table_mod_sram_id_table_5),
    .io_mod_table_mod_sram_id_table_6(MAT_io_mod_table_mod_sram_id_table_6),
    .io_mod_table_mod_sram_id_table_7(MAT_io_mod_table_mod_sram_id_table_7),
    .io_mod_table_mod_sram_id_table_8(MAT_io_mod_table_mod_sram_id_table_8),
    .io_mod_table_mod_sram_id_table_9(MAT_io_mod_table_mod_sram_id_table_9),
    .io_mod_table_mod_sram_id_table_10(MAT_io_mod_table_mod_sram_id_table_10),
    .io_mod_table_mod_sram_id_table_11(MAT_io_mod_table_mod_sram_id_table_11),
    .io_mod_table_mod_sram_id_table_12(MAT_io_mod_table_mod_sram_id_table_12),
    .io_mod_table_mod_sram_id_table_13(MAT_io_mod_table_mod_sram_id_table_13),
    .io_mod_table_mod_sram_id_table_14(MAT_io_mod_table_mod_sram_id_table_14),
    .io_mod_table_mod_sram_id_table_15(MAT_io_mod_table_mod_sram_id_table_15),
    .io_mod_table_mod_sram_id_table_16(MAT_io_mod_table_mod_sram_id_table_16),
    .io_mod_table_mod_sram_id_table_17(MAT_io_mod_table_mod_sram_id_table_17),
    .io_mod_table_mod_sram_id_table_18(MAT_io_mod_table_mod_sram_id_table_18),
    .io_mod_table_mod_sram_id_table_19(MAT_io_mod_table_mod_sram_id_table_19),
    .io_mod_table_mod_sram_id_table_20(MAT_io_mod_table_mod_sram_id_table_20),
    .io_mod_table_mod_sram_id_table_21(MAT_io_mod_table_mod_sram_id_table_21),
    .io_mod_table_mod_sram_id_table_22(MAT_io_mod_table_mod_sram_id_table_22),
    .io_mod_table_mod_sram_id_table_23(MAT_io_mod_table_mod_sram_id_table_23),
    .io_mod_table_mod_sram_id_table_24(MAT_io_mod_table_mod_sram_id_table_24),
    .io_mod_table_mod_sram_id_table_25(MAT_io_mod_table_mod_sram_id_table_25),
    .io_mod_table_mod_sram_id_table_26(MAT_io_mod_table_mod_sram_id_table_26),
    .io_mod_table_mod_sram_id_table_27(MAT_io_mod_table_mod_sram_id_table_27),
    .io_mod_table_mod_sram_id_table_28(MAT_io_mod_table_mod_sram_id_table_28),
    .io_mod_table_mod_sram_id_table_29(MAT_io_mod_table_mod_sram_id_table_29),
    .io_mod_table_mod_sram_id_table_30(MAT_io_mod_table_mod_sram_id_table_30),
    .io_mod_table_mod_sram_id_table_31(MAT_io_mod_table_mod_sram_id_table_31),
    .io_mod_table_mod_sram_id_table_32(MAT_io_mod_table_mod_sram_id_table_32),
    .io_mod_table_mod_sram_id_table_33(MAT_io_mod_table_mod_sram_id_table_33),
    .io_mod_table_mod_sram_id_table_34(MAT_io_mod_table_mod_sram_id_table_34),
    .io_mod_table_mod_sram_id_table_35(MAT_io_mod_table_mod_sram_id_table_35),
    .io_mod_table_mod_sram_id_table_36(MAT_io_mod_table_mod_sram_id_table_36),
    .io_mod_table_mod_sram_id_table_37(MAT_io_mod_table_mod_sram_id_table_37),
    .io_mod_table_mod_sram_id_table_38(MAT_io_mod_table_mod_sram_id_table_38),
    .io_mod_table_mod_sram_id_table_39(MAT_io_mod_table_mod_sram_id_table_39),
    .io_mod_table_mod_sram_id_table_40(MAT_io_mod_table_mod_sram_id_table_40),
    .io_mod_table_mod_sram_id_table_41(MAT_io_mod_table_mod_sram_id_table_41),
    .io_mod_table_mod_sram_id_table_42(MAT_io_mod_table_mod_sram_id_table_42),
    .io_mod_table_mod_sram_id_table_43(MAT_io_mod_table_mod_sram_id_table_43),
    .io_mod_table_mod_sram_id_table_44(MAT_io_mod_table_mod_sram_id_table_44),
    .io_mod_table_mod_sram_id_table_45(MAT_io_mod_table_mod_sram_id_table_45),
    .io_mod_table_mod_sram_id_table_46(MAT_io_mod_table_mod_sram_id_table_46),
    .io_mod_table_mod_sram_id_table_47(MAT_io_mod_table_mod_sram_id_table_47),
    .io_mod_table_mod_sram_id_table_48(MAT_io_mod_table_mod_sram_id_table_48),
    .io_mod_table_mod_sram_id_table_49(MAT_io_mod_table_mod_sram_id_table_49),
    .io_mod_table_mod_sram_id_table_50(MAT_io_mod_table_mod_sram_id_table_50),
    .io_mod_table_mod_sram_id_table_51(MAT_io_mod_table_mod_sram_id_table_51),
    .io_mod_table_mod_sram_id_table_52(MAT_io_mod_table_mod_sram_id_table_52),
    .io_mod_table_mod_sram_id_table_53(MAT_io_mod_table_mod_sram_id_table_53),
    .io_mod_table_mod_sram_id_table_54(MAT_io_mod_table_mod_sram_id_table_54),
    .io_mod_table_mod_sram_id_table_55(MAT_io_mod_table_mod_sram_id_table_55),
    .io_mod_table_mod_sram_id_table_56(MAT_io_mod_table_mod_sram_id_table_56),
    .io_mod_table_mod_sram_id_table_57(MAT_io_mod_table_mod_sram_id_table_57),
    .io_mod_table_mod_sram_id_table_58(MAT_io_mod_table_mod_sram_id_table_58),
    .io_mod_table_mod_sram_id_table_59(MAT_io_mod_table_mod_sram_id_table_59),
    .io_mod_table_mod_sram_id_table_60(MAT_io_mod_table_mod_sram_id_table_60),
    .io_mod_table_mod_sram_id_table_61(MAT_io_mod_table_mod_sram_id_table_61),
    .io_mod_table_mod_sram_id_table_62(MAT_io_mod_table_mod_sram_id_table_62),
    .io_mod_table_mod_sram_id_table_63(MAT_io_mod_table_mod_sram_id_table_63),
    .io_mod_table_mod_table_width(MAT_io_mod_table_mod_table_width),
    .io_mod_table_mod_table_depth(MAT_io_mod_table_mod_table_depth),
    .io_hit(MAT_io_hit),
    .io_match_value(MAT_io_match_value),
    .io_mem_cluster_0_en(MAT_io_mem_cluster_0_en),
    .io_mem_cluster_0_addr(MAT_io_mem_cluster_0_addr),
    .io_mem_cluster_0_data(MAT_io_mem_cluster_0_data),
    .io_mem_cluster_1_en(MAT_io_mem_cluster_1_en),
    .io_mem_cluster_1_addr(MAT_io_mem_cluster_1_addr),
    .io_mem_cluster_1_data(MAT_io_mem_cluster_1_data),
    .io_mem_cluster_2_en(MAT_io_mem_cluster_2_en),
    .io_mem_cluster_2_addr(MAT_io_mem_cluster_2_addr),
    .io_mem_cluster_2_data(MAT_io_mem_cluster_2_data),
    .io_mem_cluster_3_en(MAT_io_mem_cluster_3_en),
    .io_mem_cluster_3_addr(MAT_io_mem_cluster_3_addr),
    .io_mem_cluster_3_data(MAT_io_mem_cluster_3_data),
    .io_mem_cluster_4_en(MAT_io_mem_cluster_4_en),
    .io_mem_cluster_4_addr(MAT_io_mem_cluster_4_addr),
    .io_mem_cluster_4_data(MAT_io_mem_cluster_4_data),
    .io_mem_cluster_5_en(MAT_io_mem_cluster_5_en),
    .io_mem_cluster_5_addr(MAT_io_mem_cluster_5_addr),
    .io_mem_cluster_5_data(MAT_io_mem_cluster_5_data),
    .io_mem_cluster_6_en(MAT_io_mem_cluster_6_en),
    .io_mem_cluster_6_addr(MAT_io_mem_cluster_6_addr),
    .io_mem_cluster_6_data(MAT_io_mem_cluster_6_data),
    .io_mem_cluster_7_en(MAT_io_mem_cluster_7_en),
    .io_mem_cluster_7_addr(MAT_io_mem_cluster_7_addr),
    .io_mem_cluster_7_data(MAT_io_mem_cluster_7_data),
    .io_mem_cluster_8_en(MAT_io_mem_cluster_8_en),
    .io_mem_cluster_8_addr(MAT_io_mem_cluster_8_addr),
    .io_mem_cluster_8_data(MAT_io_mem_cluster_8_data),
    .io_mem_cluster_9_en(MAT_io_mem_cluster_9_en),
    .io_mem_cluster_9_addr(MAT_io_mem_cluster_9_addr),
    .io_mem_cluster_9_data(MAT_io_mem_cluster_9_data),
    .io_mem_cluster_10_en(MAT_io_mem_cluster_10_en),
    .io_mem_cluster_10_addr(MAT_io_mem_cluster_10_addr),
    .io_mem_cluster_10_data(MAT_io_mem_cluster_10_data),
    .io_mem_cluster_11_en(MAT_io_mem_cluster_11_en),
    .io_mem_cluster_11_addr(MAT_io_mem_cluster_11_addr),
    .io_mem_cluster_11_data(MAT_io_mem_cluster_11_data),
    .io_mem_cluster_12_en(MAT_io_mem_cluster_12_en),
    .io_mem_cluster_12_addr(MAT_io_mem_cluster_12_addr),
    .io_mem_cluster_12_data(MAT_io_mem_cluster_12_data),
    .io_mem_cluster_13_en(MAT_io_mem_cluster_13_en),
    .io_mem_cluster_13_addr(MAT_io_mem_cluster_13_addr),
    .io_mem_cluster_13_data(MAT_io_mem_cluster_13_data),
    .io_mem_cluster_14_en(MAT_io_mem_cluster_14_en),
    .io_mem_cluster_14_addr(MAT_io_mem_cluster_14_addr),
    .io_mem_cluster_14_data(MAT_io_mem_cluster_14_data),
    .io_mem_cluster_15_en(MAT_io_mem_cluster_15_en),
    .io_mem_cluster_15_addr(MAT_io_mem_cluster_15_addr),
    .io_mem_cluster_15_data(MAT_io_mem_cluster_15_data),
    .io_mem_cluster_16_en(MAT_io_mem_cluster_16_en),
    .io_mem_cluster_16_addr(MAT_io_mem_cluster_16_addr),
    .io_mem_cluster_16_data(MAT_io_mem_cluster_16_data),
    .io_mem_cluster_17_en(MAT_io_mem_cluster_17_en),
    .io_mem_cluster_17_addr(MAT_io_mem_cluster_17_addr),
    .io_mem_cluster_17_data(MAT_io_mem_cluster_17_data),
    .io_mem_cluster_18_en(MAT_io_mem_cluster_18_en),
    .io_mem_cluster_18_addr(MAT_io_mem_cluster_18_addr),
    .io_mem_cluster_18_data(MAT_io_mem_cluster_18_data),
    .io_mem_cluster_19_en(MAT_io_mem_cluster_19_en),
    .io_mem_cluster_19_addr(MAT_io_mem_cluster_19_addr),
    .io_mem_cluster_19_data(MAT_io_mem_cluster_19_data),
    .io_mem_cluster_20_en(MAT_io_mem_cluster_20_en),
    .io_mem_cluster_20_addr(MAT_io_mem_cluster_20_addr),
    .io_mem_cluster_20_data(MAT_io_mem_cluster_20_data),
    .io_mem_cluster_21_en(MAT_io_mem_cluster_21_en),
    .io_mem_cluster_21_addr(MAT_io_mem_cluster_21_addr),
    .io_mem_cluster_21_data(MAT_io_mem_cluster_21_data),
    .io_mem_cluster_22_en(MAT_io_mem_cluster_22_en),
    .io_mem_cluster_22_addr(MAT_io_mem_cluster_22_addr),
    .io_mem_cluster_22_data(MAT_io_mem_cluster_22_data),
    .io_mem_cluster_23_en(MAT_io_mem_cluster_23_en),
    .io_mem_cluster_23_addr(MAT_io_mem_cluster_23_addr),
    .io_mem_cluster_23_data(MAT_io_mem_cluster_23_data),
    .io_mem_cluster_24_en(MAT_io_mem_cluster_24_en),
    .io_mem_cluster_24_addr(MAT_io_mem_cluster_24_addr),
    .io_mem_cluster_24_data(MAT_io_mem_cluster_24_data),
    .io_mem_cluster_25_en(MAT_io_mem_cluster_25_en),
    .io_mem_cluster_25_addr(MAT_io_mem_cluster_25_addr),
    .io_mem_cluster_25_data(MAT_io_mem_cluster_25_data),
    .io_mem_cluster_26_en(MAT_io_mem_cluster_26_en),
    .io_mem_cluster_26_addr(MAT_io_mem_cluster_26_addr),
    .io_mem_cluster_26_data(MAT_io_mem_cluster_26_data),
    .io_mem_cluster_27_en(MAT_io_mem_cluster_27_en),
    .io_mem_cluster_27_addr(MAT_io_mem_cluster_27_addr),
    .io_mem_cluster_27_data(MAT_io_mem_cluster_27_data),
    .io_mem_cluster_28_en(MAT_io_mem_cluster_28_en),
    .io_mem_cluster_28_addr(MAT_io_mem_cluster_28_addr),
    .io_mem_cluster_28_data(MAT_io_mem_cluster_28_data),
    .io_mem_cluster_29_en(MAT_io_mem_cluster_29_en),
    .io_mem_cluster_29_addr(MAT_io_mem_cluster_29_addr),
    .io_mem_cluster_29_data(MAT_io_mem_cluster_29_data),
    .io_mem_cluster_30_en(MAT_io_mem_cluster_30_en),
    .io_mem_cluster_30_addr(MAT_io_mem_cluster_30_addr),
    .io_mem_cluster_30_data(MAT_io_mem_cluster_30_data),
    .io_mem_cluster_31_en(MAT_io_mem_cluster_31_en),
    .io_mem_cluster_31_addr(MAT_io_mem_cluster_31_addr),
    .io_mem_cluster_31_data(MAT_io_mem_cluster_31_data),
    .io_mem_cluster_32_en(MAT_io_mem_cluster_32_en),
    .io_mem_cluster_32_addr(MAT_io_mem_cluster_32_addr),
    .io_mem_cluster_32_data(MAT_io_mem_cluster_32_data),
    .io_mem_cluster_33_en(MAT_io_mem_cluster_33_en),
    .io_mem_cluster_33_addr(MAT_io_mem_cluster_33_addr),
    .io_mem_cluster_33_data(MAT_io_mem_cluster_33_data),
    .io_mem_cluster_34_en(MAT_io_mem_cluster_34_en),
    .io_mem_cluster_34_addr(MAT_io_mem_cluster_34_addr),
    .io_mem_cluster_34_data(MAT_io_mem_cluster_34_data),
    .io_mem_cluster_35_en(MAT_io_mem_cluster_35_en),
    .io_mem_cluster_35_addr(MAT_io_mem_cluster_35_addr),
    .io_mem_cluster_35_data(MAT_io_mem_cluster_35_data),
    .io_mem_cluster_36_en(MAT_io_mem_cluster_36_en),
    .io_mem_cluster_36_addr(MAT_io_mem_cluster_36_addr),
    .io_mem_cluster_36_data(MAT_io_mem_cluster_36_data),
    .io_mem_cluster_37_en(MAT_io_mem_cluster_37_en),
    .io_mem_cluster_37_addr(MAT_io_mem_cluster_37_addr),
    .io_mem_cluster_37_data(MAT_io_mem_cluster_37_data),
    .io_mem_cluster_38_en(MAT_io_mem_cluster_38_en),
    .io_mem_cluster_38_addr(MAT_io_mem_cluster_38_addr),
    .io_mem_cluster_38_data(MAT_io_mem_cluster_38_data),
    .io_mem_cluster_39_en(MAT_io_mem_cluster_39_en),
    .io_mem_cluster_39_addr(MAT_io_mem_cluster_39_addr),
    .io_mem_cluster_39_data(MAT_io_mem_cluster_39_data),
    .io_mem_cluster_40_en(MAT_io_mem_cluster_40_en),
    .io_mem_cluster_40_addr(MAT_io_mem_cluster_40_addr),
    .io_mem_cluster_40_data(MAT_io_mem_cluster_40_data),
    .io_mem_cluster_41_en(MAT_io_mem_cluster_41_en),
    .io_mem_cluster_41_addr(MAT_io_mem_cluster_41_addr),
    .io_mem_cluster_41_data(MAT_io_mem_cluster_41_data),
    .io_mem_cluster_42_en(MAT_io_mem_cluster_42_en),
    .io_mem_cluster_42_addr(MAT_io_mem_cluster_42_addr),
    .io_mem_cluster_42_data(MAT_io_mem_cluster_42_data),
    .io_mem_cluster_43_en(MAT_io_mem_cluster_43_en),
    .io_mem_cluster_43_addr(MAT_io_mem_cluster_43_addr),
    .io_mem_cluster_43_data(MAT_io_mem_cluster_43_data),
    .io_mem_cluster_44_en(MAT_io_mem_cluster_44_en),
    .io_mem_cluster_44_addr(MAT_io_mem_cluster_44_addr),
    .io_mem_cluster_44_data(MAT_io_mem_cluster_44_data),
    .io_mem_cluster_45_en(MAT_io_mem_cluster_45_en),
    .io_mem_cluster_45_addr(MAT_io_mem_cluster_45_addr),
    .io_mem_cluster_45_data(MAT_io_mem_cluster_45_data),
    .io_mem_cluster_46_en(MAT_io_mem_cluster_46_en),
    .io_mem_cluster_46_addr(MAT_io_mem_cluster_46_addr),
    .io_mem_cluster_46_data(MAT_io_mem_cluster_46_data),
    .io_mem_cluster_47_en(MAT_io_mem_cluster_47_en),
    .io_mem_cluster_47_addr(MAT_io_mem_cluster_47_addr),
    .io_mem_cluster_47_data(MAT_io_mem_cluster_47_data),
    .io_mem_cluster_48_en(MAT_io_mem_cluster_48_en),
    .io_mem_cluster_48_addr(MAT_io_mem_cluster_48_addr),
    .io_mem_cluster_48_data(MAT_io_mem_cluster_48_data),
    .io_mem_cluster_49_en(MAT_io_mem_cluster_49_en),
    .io_mem_cluster_49_addr(MAT_io_mem_cluster_49_addr),
    .io_mem_cluster_49_data(MAT_io_mem_cluster_49_data),
    .io_mem_cluster_50_en(MAT_io_mem_cluster_50_en),
    .io_mem_cluster_50_addr(MAT_io_mem_cluster_50_addr),
    .io_mem_cluster_50_data(MAT_io_mem_cluster_50_data),
    .io_mem_cluster_51_en(MAT_io_mem_cluster_51_en),
    .io_mem_cluster_51_addr(MAT_io_mem_cluster_51_addr),
    .io_mem_cluster_51_data(MAT_io_mem_cluster_51_data),
    .io_mem_cluster_52_en(MAT_io_mem_cluster_52_en),
    .io_mem_cluster_52_addr(MAT_io_mem_cluster_52_addr),
    .io_mem_cluster_52_data(MAT_io_mem_cluster_52_data),
    .io_mem_cluster_53_en(MAT_io_mem_cluster_53_en),
    .io_mem_cluster_53_addr(MAT_io_mem_cluster_53_addr),
    .io_mem_cluster_53_data(MAT_io_mem_cluster_53_data),
    .io_mem_cluster_54_en(MAT_io_mem_cluster_54_en),
    .io_mem_cluster_54_addr(MAT_io_mem_cluster_54_addr),
    .io_mem_cluster_54_data(MAT_io_mem_cluster_54_data),
    .io_mem_cluster_55_en(MAT_io_mem_cluster_55_en),
    .io_mem_cluster_55_addr(MAT_io_mem_cluster_55_addr),
    .io_mem_cluster_55_data(MAT_io_mem_cluster_55_data),
    .io_mem_cluster_56_en(MAT_io_mem_cluster_56_en),
    .io_mem_cluster_56_addr(MAT_io_mem_cluster_56_addr),
    .io_mem_cluster_56_data(MAT_io_mem_cluster_56_data),
    .io_mem_cluster_57_en(MAT_io_mem_cluster_57_en),
    .io_mem_cluster_57_addr(MAT_io_mem_cluster_57_addr),
    .io_mem_cluster_57_data(MAT_io_mem_cluster_57_data),
    .io_mem_cluster_58_en(MAT_io_mem_cluster_58_en),
    .io_mem_cluster_58_addr(MAT_io_mem_cluster_58_addr),
    .io_mem_cluster_58_data(MAT_io_mem_cluster_58_data),
    .io_mem_cluster_59_en(MAT_io_mem_cluster_59_en),
    .io_mem_cluster_59_addr(MAT_io_mem_cluster_59_addr),
    .io_mem_cluster_59_data(MAT_io_mem_cluster_59_data),
    .io_mem_cluster_60_en(MAT_io_mem_cluster_60_en),
    .io_mem_cluster_60_addr(MAT_io_mem_cluster_60_addr),
    .io_mem_cluster_60_data(MAT_io_mem_cluster_60_data),
    .io_mem_cluster_61_en(MAT_io_mem_cluster_61_en),
    .io_mem_cluster_61_addr(MAT_io_mem_cluster_61_addr),
    .io_mem_cluster_61_data(MAT_io_mem_cluster_61_data),
    .io_mem_cluster_62_en(MAT_io_mem_cluster_62_en),
    .io_mem_cluster_62_addr(MAT_io_mem_cluster_62_addr),
    .io_mem_cluster_62_data(MAT_io_mem_cluster_62_data),
    .io_mem_cluster_63_en(MAT_io_mem_cluster_63_en),
    .io_mem_cluster_63_addr(MAT_io_mem_cluster_63_addr),
    .io_mem_cluster_63_data(MAT_io_mem_cluster_63_data)
  );
  Executor EXE ( // @[processor.scala 15:21]
    .clock(EXE_clock),
    .io_pipe_phv_in_data_0(EXE_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(EXE_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(EXE_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(EXE_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(EXE_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(EXE_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(EXE_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(EXE_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(EXE_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(EXE_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(EXE_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(EXE_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(EXE_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(EXE_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(EXE_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(EXE_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(EXE_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(EXE_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(EXE_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(EXE_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(EXE_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(EXE_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(EXE_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(EXE_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(EXE_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(EXE_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(EXE_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(EXE_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(EXE_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(EXE_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(EXE_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(EXE_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(EXE_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(EXE_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(EXE_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(EXE_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(EXE_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(EXE_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(EXE_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(EXE_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(EXE_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(EXE_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(EXE_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(EXE_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(EXE_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(EXE_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(EXE_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(EXE_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(EXE_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(EXE_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(EXE_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(EXE_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(EXE_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(EXE_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(EXE_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(EXE_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(EXE_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(EXE_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(EXE_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(EXE_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(EXE_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(EXE_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(EXE_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(EXE_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(EXE_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(EXE_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(EXE_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(EXE_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(EXE_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(EXE_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(EXE_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(EXE_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(EXE_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(EXE_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(EXE_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(EXE_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(EXE_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(EXE_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(EXE_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(EXE_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(EXE_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(EXE_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(EXE_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(EXE_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(EXE_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(EXE_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(EXE_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(EXE_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(EXE_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(EXE_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(EXE_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(EXE_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(EXE_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(EXE_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(EXE_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(EXE_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(EXE_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(EXE_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(EXE_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(EXE_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(EXE_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(EXE_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(EXE_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(EXE_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(EXE_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(EXE_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(EXE_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(EXE_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(EXE_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(EXE_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(EXE_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(EXE_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(EXE_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(EXE_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(EXE_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(EXE_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(EXE_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(EXE_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(EXE_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(EXE_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(EXE_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(EXE_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(EXE_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(EXE_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(EXE_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(EXE_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(EXE_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(EXE_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(EXE_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(EXE_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(EXE_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(EXE_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(EXE_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(EXE_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(EXE_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(EXE_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(EXE_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(EXE_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(EXE_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(EXE_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(EXE_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(EXE_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(EXE_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(EXE_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(EXE_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(EXE_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(EXE_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(EXE_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(EXE_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(EXE_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(EXE_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(EXE_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(EXE_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(EXE_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(EXE_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(EXE_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(EXE_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(EXE_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(EXE_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(EXE_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(EXE_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(EXE_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(EXE_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(EXE_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(EXE_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(EXE_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(EXE_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(EXE_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(EXE_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(EXE_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(EXE_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(EXE_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(EXE_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(EXE_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(EXE_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(EXE_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(EXE_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(EXE_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(EXE_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(EXE_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(EXE_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(EXE_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(EXE_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(EXE_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(EXE_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(EXE_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(EXE_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(EXE_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(EXE_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(EXE_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(EXE_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(EXE_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(EXE_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(EXE_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(EXE_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(EXE_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(EXE_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(EXE_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(EXE_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(EXE_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(EXE_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(EXE_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(EXE_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(EXE_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(EXE_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(EXE_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(EXE_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(EXE_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(EXE_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(EXE_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(EXE_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(EXE_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(EXE_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(EXE_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(EXE_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(EXE_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(EXE_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(EXE_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(EXE_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(EXE_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(EXE_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(EXE_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(EXE_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(EXE_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(EXE_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(EXE_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(EXE_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(EXE_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(EXE_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(EXE_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(EXE_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(EXE_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(EXE_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(EXE_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(EXE_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(EXE_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(EXE_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(EXE_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(EXE_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(EXE_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(EXE_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(EXE_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(EXE_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(EXE_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(EXE_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(EXE_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(EXE_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(EXE_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(EXE_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(EXE_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(EXE_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(EXE_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(EXE_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(EXE_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(EXE_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(EXE_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(EXE_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(EXE_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(EXE_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(EXE_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(EXE_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(EXE_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(EXE_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(EXE_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(EXE_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(EXE_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(EXE_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(EXE_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(EXE_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(EXE_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(EXE_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(EXE_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(EXE_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(EXE_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(EXE_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(EXE_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(EXE_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(EXE_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(EXE_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(EXE_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(EXE_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(EXE_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(EXE_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(EXE_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(EXE_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(EXE_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(EXE_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(EXE_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(EXE_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(EXE_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(EXE_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(EXE_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(EXE_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(EXE_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(EXE_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(EXE_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(EXE_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(EXE_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(EXE_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(EXE_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(EXE_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(EXE_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(EXE_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(EXE_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(EXE_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(EXE_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(EXE_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(EXE_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(EXE_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(EXE_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(EXE_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(EXE_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(EXE_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(EXE_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(EXE_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(EXE_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(EXE_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(EXE_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(EXE_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(EXE_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(EXE_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(EXE_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(EXE_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(EXE_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(EXE_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(EXE_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(EXE_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(EXE_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(EXE_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(EXE_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(EXE_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(EXE_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(EXE_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(EXE_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(EXE_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(EXE_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(EXE_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(EXE_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(EXE_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(EXE_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(EXE_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(EXE_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(EXE_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(EXE_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(EXE_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(EXE_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(EXE_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(EXE_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(EXE_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(EXE_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(EXE_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(EXE_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(EXE_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(EXE_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(EXE_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(EXE_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(EXE_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(EXE_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(EXE_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(EXE_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(EXE_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(EXE_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(EXE_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(EXE_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(EXE_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(EXE_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(EXE_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(EXE_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(EXE_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(EXE_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(EXE_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(EXE_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(EXE_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(EXE_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(EXE_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(EXE_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(EXE_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(EXE_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(EXE_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(EXE_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(EXE_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(EXE_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(EXE_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(EXE_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(EXE_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(EXE_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(EXE_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(EXE_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(EXE_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(EXE_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(EXE_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(EXE_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(EXE_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(EXE_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(EXE_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(EXE_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(EXE_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(EXE_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(EXE_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(EXE_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(EXE_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(EXE_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(EXE_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(EXE_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(EXE_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(EXE_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(EXE_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(EXE_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(EXE_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(EXE_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(EXE_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(EXE_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(EXE_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(EXE_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(EXE_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(EXE_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(EXE_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(EXE_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(EXE_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(EXE_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(EXE_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(EXE_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(EXE_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(EXE_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(EXE_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(EXE_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(EXE_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(EXE_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(EXE_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(EXE_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(EXE_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(EXE_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(EXE_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(EXE_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(EXE_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(EXE_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(EXE_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(EXE_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(EXE_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(EXE_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(EXE_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(EXE_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(EXE_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(EXE_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(EXE_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(EXE_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(EXE_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(EXE_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(EXE_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(EXE_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(EXE_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(EXE_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(EXE_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(EXE_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(EXE_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(EXE_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(EXE_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(EXE_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(EXE_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(EXE_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(EXE_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(EXE_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(EXE_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(EXE_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(EXE_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(EXE_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(EXE_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(EXE_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(EXE_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(EXE_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(EXE_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(EXE_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(EXE_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(EXE_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(EXE_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(EXE_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(EXE_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(EXE_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(EXE_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(EXE_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(EXE_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(EXE_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(EXE_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(EXE_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(EXE_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(EXE_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(EXE_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(EXE_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(EXE_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(EXE_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(EXE_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(EXE_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(EXE_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(EXE_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(EXE_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(EXE_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(EXE_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(EXE_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(EXE_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(EXE_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(EXE_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(EXE_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(EXE_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(EXE_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(EXE_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(EXE_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(EXE_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(EXE_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(EXE_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(EXE_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(EXE_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(EXE_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(EXE_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(EXE_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(EXE_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(EXE_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(EXE_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(EXE_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(EXE_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(EXE_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(EXE_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(EXE_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(EXE_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(EXE_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(EXE_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(EXE_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(EXE_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(EXE_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(EXE_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(EXE_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(EXE_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(EXE_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(EXE_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(EXE_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(EXE_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(EXE_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(EXE_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(EXE_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(EXE_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(EXE_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(EXE_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(EXE_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(EXE_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(EXE_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(EXE_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(EXE_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(EXE_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(EXE_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(EXE_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(EXE_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(EXE_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(EXE_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(EXE_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(EXE_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(EXE_io_pipe_phv_out_next_config_id),
    .io_hit(EXE_io_hit),
    .io_match_value(EXE_io_match_value),
    .io_action_mod_en_0(EXE_io_action_mod_en_0),
    .io_action_mod_en_1(EXE_io_action_mod_en_1),
    .io_action_mod_addr(EXE_io_action_mod_addr),
    .io_action_mod_data_0(EXE_io_action_mod_data_0),
    .io_action_mod_data_1(EXE_io_action_mod_data_1)
  );
  assign io_pipe_phv_out_data_0 = EXE_io_pipe_phv_out_data_0; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_1 = EXE_io_pipe_phv_out_data_1; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_2 = EXE_io_pipe_phv_out_data_2; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_3 = EXE_io_pipe_phv_out_data_3; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_4 = EXE_io_pipe_phv_out_data_4; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_5 = EXE_io_pipe_phv_out_data_5; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_6 = EXE_io_pipe_phv_out_data_6; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_7 = EXE_io_pipe_phv_out_data_7; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_8 = EXE_io_pipe_phv_out_data_8; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_9 = EXE_io_pipe_phv_out_data_9; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_10 = EXE_io_pipe_phv_out_data_10; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_11 = EXE_io_pipe_phv_out_data_11; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_12 = EXE_io_pipe_phv_out_data_12; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_13 = EXE_io_pipe_phv_out_data_13; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_14 = EXE_io_pipe_phv_out_data_14; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_15 = EXE_io_pipe_phv_out_data_15; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_16 = EXE_io_pipe_phv_out_data_16; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_17 = EXE_io_pipe_phv_out_data_17; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_18 = EXE_io_pipe_phv_out_data_18; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_19 = EXE_io_pipe_phv_out_data_19; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_20 = EXE_io_pipe_phv_out_data_20; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_21 = EXE_io_pipe_phv_out_data_21; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_22 = EXE_io_pipe_phv_out_data_22; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_23 = EXE_io_pipe_phv_out_data_23; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_24 = EXE_io_pipe_phv_out_data_24; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_25 = EXE_io_pipe_phv_out_data_25; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_26 = EXE_io_pipe_phv_out_data_26; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_27 = EXE_io_pipe_phv_out_data_27; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_28 = EXE_io_pipe_phv_out_data_28; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_29 = EXE_io_pipe_phv_out_data_29; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_30 = EXE_io_pipe_phv_out_data_30; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_31 = EXE_io_pipe_phv_out_data_31; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_32 = EXE_io_pipe_phv_out_data_32; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_33 = EXE_io_pipe_phv_out_data_33; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_34 = EXE_io_pipe_phv_out_data_34; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_35 = EXE_io_pipe_phv_out_data_35; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_36 = EXE_io_pipe_phv_out_data_36; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_37 = EXE_io_pipe_phv_out_data_37; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_38 = EXE_io_pipe_phv_out_data_38; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_39 = EXE_io_pipe_phv_out_data_39; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_40 = EXE_io_pipe_phv_out_data_40; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_41 = EXE_io_pipe_phv_out_data_41; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_42 = EXE_io_pipe_phv_out_data_42; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_43 = EXE_io_pipe_phv_out_data_43; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_44 = EXE_io_pipe_phv_out_data_44; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_45 = EXE_io_pipe_phv_out_data_45; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_46 = EXE_io_pipe_phv_out_data_46; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_47 = EXE_io_pipe_phv_out_data_47; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_48 = EXE_io_pipe_phv_out_data_48; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_49 = EXE_io_pipe_phv_out_data_49; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_50 = EXE_io_pipe_phv_out_data_50; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_51 = EXE_io_pipe_phv_out_data_51; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_52 = EXE_io_pipe_phv_out_data_52; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_53 = EXE_io_pipe_phv_out_data_53; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_54 = EXE_io_pipe_phv_out_data_54; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_55 = EXE_io_pipe_phv_out_data_55; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_56 = EXE_io_pipe_phv_out_data_56; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_57 = EXE_io_pipe_phv_out_data_57; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_58 = EXE_io_pipe_phv_out_data_58; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_59 = EXE_io_pipe_phv_out_data_59; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_60 = EXE_io_pipe_phv_out_data_60; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_61 = EXE_io_pipe_phv_out_data_61; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_62 = EXE_io_pipe_phv_out_data_62; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_63 = EXE_io_pipe_phv_out_data_63; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_64 = EXE_io_pipe_phv_out_data_64; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_65 = EXE_io_pipe_phv_out_data_65; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_66 = EXE_io_pipe_phv_out_data_66; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_67 = EXE_io_pipe_phv_out_data_67; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_68 = EXE_io_pipe_phv_out_data_68; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_69 = EXE_io_pipe_phv_out_data_69; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_70 = EXE_io_pipe_phv_out_data_70; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_71 = EXE_io_pipe_phv_out_data_71; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_72 = EXE_io_pipe_phv_out_data_72; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_73 = EXE_io_pipe_phv_out_data_73; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_74 = EXE_io_pipe_phv_out_data_74; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_75 = EXE_io_pipe_phv_out_data_75; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_76 = EXE_io_pipe_phv_out_data_76; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_77 = EXE_io_pipe_phv_out_data_77; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_78 = EXE_io_pipe_phv_out_data_78; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_79 = EXE_io_pipe_phv_out_data_79; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_80 = EXE_io_pipe_phv_out_data_80; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_81 = EXE_io_pipe_phv_out_data_81; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_82 = EXE_io_pipe_phv_out_data_82; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_83 = EXE_io_pipe_phv_out_data_83; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_84 = EXE_io_pipe_phv_out_data_84; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_85 = EXE_io_pipe_phv_out_data_85; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_86 = EXE_io_pipe_phv_out_data_86; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_87 = EXE_io_pipe_phv_out_data_87; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_88 = EXE_io_pipe_phv_out_data_88; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_89 = EXE_io_pipe_phv_out_data_89; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_90 = EXE_io_pipe_phv_out_data_90; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_91 = EXE_io_pipe_phv_out_data_91; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_92 = EXE_io_pipe_phv_out_data_92; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_93 = EXE_io_pipe_phv_out_data_93; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_94 = EXE_io_pipe_phv_out_data_94; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_95 = EXE_io_pipe_phv_out_data_95; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_96 = EXE_io_pipe_phv_out_data_96; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_97 = EXE_io_pipe_phv_out_data_97; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_98 = EXE_io_pipe_phv_out_data_98; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_99 = EXE_io_pipe_phv_out_data_99; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_100 = EXE_io_pipe_phv_out_data_100; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_101 = EXE_io_pipe_phv_out_data_101; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_102 = EXE_io_pipe_phv_out_data_102; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_103 = EXE_io_pipe_phv_out_data_103; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_104 = EXE_io_pipe_phv_out_data_104; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_105 = EXE_io_pipe_phv_out_data_105; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_106 = EXE_io_pipe_phv_out_data_106; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_107 = EXE_io_pipe_phv_out_data_107; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_108 = EXE_io_pipe_phv_out_data_108; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_109 = EXE_io_pipe_phv_out_data_109; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_110 = EXE_io_pipe_phv_out_data_110; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_111 = EXE_io_pipe_phv_out_data_111; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_112 = EXE_io_pipe_phv_out_data_112; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_113 = EXE_io_pipe_phv_out_data_113; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_114 = EXE_io_pipe_phv_out_data_114; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_115 = EXE_io_pipe_phv_out_data_115; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_116 = EXE_io_pipe_phv_out_data_116; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_117 = EXE_io_pipe_phv_out_data_117; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_118 = EXE_io_pipe_phv_out_data_118; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_119 = EXE_io_pipe_phv_out_data_119; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_120 = EXE_io_pipe_phv_out_data_120; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_121 = EXE_io_pipe_phv_out_data_121; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_122 = EXE_io_pipe_phv_out_data_122; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_123 = EXE_io_pipe_phv_out_data_123; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_124 = EXE_io_pipe_phv_out_data_124; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_125 = EXE_io_pipe_phv_out_data_125; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_126 = EXE_io_pipe_phv_out_data_126; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_127 = EXE_io_pipe_phv_out_data_127; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_128 = EXE_io_pipe_phv_out_data_128; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_129 = EXE_io_pipe_phv_out_data_129; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_130 = EXE_io_pipe_phv_out_data_130; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_131 = EXE_io_pipe_phv_out_data_131; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_132 = EXE_io_pipe_phv_out_data_132; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_133 = EXE_io_pipe_phv_out_data_133; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_134 = EXE_io_pipe_phv_out_data_134; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_135 = EXE_io_pipe_phv_out_data_135; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_136 = EXE_io_pipe_phv_out_data_136; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_137 = EXE_io_pipe_phv_out_data_137; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_138 = EXE_io_pipe_phv_out_data_138; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_139 = EXE_io_pipe_phv_out_data_139; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_140 = EXE_io_pipe_phv_out_data_140; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_141 = EXE_io_pipe_phv_out_data_141; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_142 = EXE_io_pipe_phv_out_data_142; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_143 = EXE_io_pipe_phv_out_data_143; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_144 = EXE_io_pipe_phv_out_data_144; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_145 = EXE_io_pipe_phv_out_data_145; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_146 = EXE_io_pipe_phv_out_data_146; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_147 = EXE_io_pipe_phv_out_data_147; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_148 = EXE_io_pipe_phv_out_data_148; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_149 = EXE_io_pipe_phv_out_data_149; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_150 = EXE_io_pipe_phv_out_data_150; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_151 = EXE_io_pipe_phv_out_data_151; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_152 = EXE_io_pipe_phv_out_data_152; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_153 = EXE_io_pipe_phv_out_data_153; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_154 = EXE_io_pipe_phv_out_data_154; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_155 = EXE_io_pipe_phv_out_data_155; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_156 = EXE_io_pipe_phv_out_data_156; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_157 = EXE_io_pipe_phv_out_data_157; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_158 = EXE_io_pipe_phv_out_data_158; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_159 = EXE_io_pipe_phv_out_data_159; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_160 = EXE_io_pipe_phv_out_data_160; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_161 = EXE_io_pipe_phv_out_data_161; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_162 = EXE_io_pipe_phv_out_data_162; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_163 = EXE_io_pipe_phv_out_data_163; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_164 = EXE_io_pipe_phv_out_data_164; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_165 = EXE_io_pipe_phv_out_data_165; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_166 = EXE_io_pipe_phv_out_data_166; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_167 = EXE_io_pipe_phv_out_data_167; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_168 = EXE_io_pipe_phv_out_data_168; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_169 = EXE_io_pipe_phv_out_data_169; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_170 = EXE_io_pipe_phv_out_data_170; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_171 = EXE_io_pipe_phv_out_data_171; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_172 = EXE_io_pipe_phv_out_data_172; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_173 = EXE_io_pipe_phv_out_data_173; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_174 = EXE_io_pipe_phv_out_data_174; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_175 = EXE_io_pipe_phv_out_data_175; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_176 = EXE_io_pipe_phv_out_data_176; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_177 = EXE_io_pipe_phv_out_data_177; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_178 = EXE_io_pipe_phv_out_data_178; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_179 = EXE_io_pipe_phv_out_data_179; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_180 = EXE_io_pipe_phv_out_data_180; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_181 = EXE_io_pipe_phv_out_data_181; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_182 = EXE_io_pipe_phv_out_data_182; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_183 = EXE_io_pipe_phv_out_data_183; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_184 = EXE_io_pipe_phv_out_data_184; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_185 = EXE_io_pipe_phv_out_data_185; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_186 = EXE_io_pipe_phv_out_data_186; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_187 = EXE_io_pipe_phv_out_data_187; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_188 = EXE_io_pipe_phv_out_data_188; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_189 = EXE_io_pipe_phv_out_data_189; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_190 = EXE_io_pipe_phv_out_data_190; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_191 = EXE_io_pipe_phv_out_data_191; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_192 = EXE_io_pipe_phv_out_data_192; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_193 = EXE_io_pipe_phv_out_data_193; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_194 = EXE_io_pipe_phv_out_data_194; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_195 = EXE_io_pipe_phv_out_data_195; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_196 = EXE_io_pipe_phv_out_data_196; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_197 = EXE_io_pipe_phv_out_data_197; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_198 = EXE_io_pipe_phv_out_data_198; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_199 = EXE_io_pipe_phv_out_data_199; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_200 = EXE_io_pipe_phv_out_data_200; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_201 = EXE_io_pipe_phv_out_data_201; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_202 = EXE_io_pipe_phv_out_data_202; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_203 = EXE_io_pipe_phv_out_data_203; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_204 = EXE_io_pipe_phv_out_data_204; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_205 = EXE_io_pipe_phv_out_data_205; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_206 = EXE_io_pipe_phv_out_data_206; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_207 = EXE_io_pipe_phv_out_data_207; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_208 = EXE_io_pipe_phv_out_data_208; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_209 = EXE_io_pipe_phv_out_data_209; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_210 = EXE_io_pipe_phv_out_data_210; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_211 = EXE_io_pipe_phv_out_data_211; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_212 = EXE_io_pipe_phv_out_data_212; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_213 = EXE_io_pipe_phv_out_data_213; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_214 = EXE_io_pipe_phv_out_data_214; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_215 = EXE_io_pipe_phv_out_data_215; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_216 = EXE_io_pipe_phv_out_data_216; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_217 = EXE_io_pipe_phv_out_data_217; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_218 = EXE_io_pipe_phv_out_data_218; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_219 = EXE_io_pipe_phv_out_data_219; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_220 = EXE_io_pipe_phv_out_data_220; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_221 = EXE_io_pipe_phv_out_data_221; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_222 = EXE_io_pipe_phv_out_data_222; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_223 = EXE_io_pipe_phv_out_data_223; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_224 = EXE_io_pipe_phv_out_data_224; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_225 = EXE_io_pipe_phv_out_data_225; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_226 = EXE_io_pipe_phv_out_data_226; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_227 = EXE_io_pipe_phv_out_data_227; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_228 = EXE_io_pipe_phv_out_data_228; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_229 = EXE_io_pipe_phv_out_data_229; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_230 = EXE_io_pipe_phv_out_data_230; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_231 = EXE_io_pipe_phv_out_data_231; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_232 = EXE_io_pipe_phv_out_data_232; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_233 = EXE_io_pipe_phv_out_data_233; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_234 = EXE_io_pipe_phv_out_data_234; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_235 = EXE_io_pipe_phv_out_data_235; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_236 = EXE_io_pipe_phv_out_data_236; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_237 = EXE_io_pipe_phv_out_data_237; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_238 = EXE_io_pipe_phv_out_data_238; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_239 = EXE_io_pipe_phv_out_data_239; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_240 = EXE_io_pipe_phv_out_data_240; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_241 = EXE_io_pipe_phv_out_data_241; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_242 = EXE_io_pipe_phv_out_data_242; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_243 = EXE_io_pipe_phv_out_data_243; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_244 = EXE_io_pipe_phv_out_data_244; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_245 = EXE_io_pipe_phv_out_data_245; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_246 = EXE_io_pipe_phv_out_data_246; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_247 = EXE_io_pipe_phv_out_data_247; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_248 = EXE_io_pipe_phv_out_data_248; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_249 = EXE_io_pipe_phv_out_data_249; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_250 = EXE_io_pipe_phv_out_data_250; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_251 = EXE_io_pipe_phv_out_data_251; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_252 = EXE_io_pipe_phv_out_data_252; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_253 = EXE_io_pipe_phv_out_data_253; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_254 = EXE_io_pipe_phv_out_data_254; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_255 = EXE_io_pipe_phv_out_data_255; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_0 = EXE_io_pipe_phv_out_header_0; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_1 = EXE_io_pipe_phv_out_header_1; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_2 = EXE_io_pipe_phv_out_header_2; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_3 = EXE_io_pipe_phv_out_header_3; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_4 = EXE_io_pipe_phv_out_header_4; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_5 = EXE_io_pipe_phv_out_header_5; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_6 = EXE_io_pipe_phv_out_header_6; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_7 = EXE_io_pipe_phv_out_header_7; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_8 = EXE_io_pipe_phv_out_header_8; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_9 = EXE_io_pipe_phv_out_header_9; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_10 = EXE_io_pipe_phv_out_header_10; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_11 = EXE_io_pipe_phv_out_header_11; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_12 = EXE_io_pipe_phv_out_header_12; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_13 = EXE_io_pipe_phv_out_header_13; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_14 = EXE_io_pipe_phv_out_header_14; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_15 = EXE_io_pipe_phv_out_header_15; // @[processor.scala 29:24]
  assign io_pipe_phv_out_parse_current_state = EXE_io_pipe_phv_out_parse_current_state; // @[processor.scala 29:24]
  assign io_pipe_phv_out_parse_current_offset = EXE_io_pipe_phv_out_parse_current_offset; // @[processor.scala 29:24]
  assign io_pipe_phv_out_parse_transition_field = EXE_io_pipe_phv_out_parse_transition_field; // @[processor.scala 29:24]
  assign io_pipe_phv_out_next_processor_id = EXE_io_pipe_phv_out_next_processor_id; // @[processor.scala 29:24]
  assign io_pipe_phv_out_next_config_id = EXE_io_pipe_phv_out_next_config_id; // @[processor.scala 29:24]
  assign io_mem_cluster_0_en = MAT_io_mem_cluster_0_en; // @[processor.scala 22:24]
  assign io_mem_cluster_0_addr = MAT_io_mem_cluster_0_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_1_en = MAT_io_mem_cluster_1_en; // @[processor.scala 22:24]
  assign io_mem_cluster_1_addr = MAT_io_mem_cluster_1_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_2_en = MAT_io_mem_cluster_2_en; // @[processor.scala 22:24]
  assign io_mem_cluster_2_addr = MAT_io_mem_cluster_2_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_3_en = MAT_io_mem_cluster_3_en; // @[processor.scala 22:24]
  assign io_mem_cluster_3_addr = MAT_io_mem_cluster_3_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_4_en = MAT_io_mem_cluster_4_en; // @[processor.scala 22:24]
  assign io_mem_cluster_4_addr = MAT_io_mem_cluster_4_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_5_en = MAT_io_mem_cluster_5_en; // @[processor.scala 22:24]
  assign io_mem_cluster_5_addr = MAT_io_mem_cluster_5_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_6_en = MAT_io_mem_cluster_6_en; // @[processor.scala 22:24]
  assign io_mem_cluster_6_addr = MAT_io_mem_cluster_6_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_7_en = MAT_io_mem_cluster_7_en; // @[processor.scala 22:24]
  assign io_mem_cluster_7_addr = MAT_io_mem_cluster_7_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_8_en = MAT_io_mem_cluster_8_en; // @[processor.scala 22:24]
  assign io_mem_cluster_8_addr = MAT_io_mem_cluster_8_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_9_en = MAT_io_mem_cluster_9_en; // @[processor.scala 22:24]
  assign io_mem_cluster_9_addr = MAT_io_mem_cluster_9_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_10_en = MAT_io_mem_cluster_10_en; // @[processor.scala 22:24]
  assign io_mem_cluster_10_addr = MAT_io_mem_cluster_10_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_11_en = MAT_io_mem_cluster_11_en; // @[processor.scala 22:24]
  assign io_mem_cluster_11_addr = MAT_io_mem_cluster_11_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_12_en = MAT_io_mem_cluster_12_en; // @[processor.scala 22:24]
  assign io_mem_cluster_12_addr = MAT_io_mem_cluster_12_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_13_en = MAT_io_mem_cluster_13_en; // @[processor.scala 22:24]
  assign io_mem_cluster_13_addr = MAT_io_mem_cluster_13_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_14_en = MAT_io_mem_cluster_14_en; // @[processor.scala 22:24]
  assign io_mem_cluster_14_addr = MAT_io_mem_cluster_14_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_15_en = MAT_io_mem_cluster_15_en; // @[processor.scala 22:24]
  assign io_mem_cluster_15_addr = MAT_io_mem_cluster_15_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_16_en = MAT_io_mem_cluster_16_en; // @[processor.scala 22:24]
  assign io_mem_cluster_16_addr = MAT_io_mem_cluster_16_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_17_en = MAT_io_mem_cluster_17_en; // @[processor.scala 22:24]
  assign io_mem_cluster_17_addr = MAT_io_mem_cluster_17_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_18_en = MAT_io_mem_cluster_18_en; // @[processor.scala 22:24]
  assign io_mem_cluster_18_addr = MAT_io_mem_cluster_18_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_19_en = MAT_io_mem_cluster_19_en; // @[processor.scala 22:24]
  assign io_mem_cluster_19_addr = MAT_io_mem_cluster_19_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_20_en = MAT_io_mem_cluster_20_en; // @[processor.scala 22:24]
  assign io_mem_cluster_20_addr = MAT_io_mem_cluster_20_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_21_en = MAT_io_mem_cluster_21_en; // @[processor.scala 22:24]
  assign io_mem_cluster_21_addr = MAT_io_mem_cluster_21_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_22_en = MAT_io_mem_cluster_22_en; // @[processor.scala 22:24]
  assign io_mem_cluster_22_addr = MAT_io_mem_cluster_22_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_23_en = MAT_io_mem_cluster_23_en; // @[processor.scala 22:24]
  assign io_mem_cluster_23_addr = MAT_io_mem_cluster_23_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_24_en = MAT_io_mem_cluster_24_en; // @[processor.scala 22:24]
  assign io_mem_cluster_24_addr = MAT_io_mem_cluster_24_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_25_en = MAT_io_mem_cluster_25_en; // @[processor.scala 22:24]
  assign io_mem_cluster_25_addr = MAT_io_mem_cluster_25_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_26_en = MAT_io_mem_cluster_26_en; // @[processor.scala 22:24]
  assign io_mem_cluster_26_addr = MAT_io_mem_cluster_26_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_27_en = MAT_io_mem_cluster_27_en; // @[processor.scala 22:24]
  assign io_mem_cluster_27_addr = MAT_io_mem_cluster_27_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_28_en = MAT_io_mem_cluster_28_en; // @[processor.scala 22:24]
  assign io_mem_cluster_28_addr = MAT_io_mem_cluster_28_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_29_en = MAT_io_mem_cluster_29_en; // @[processor.scala 22:24]
  assign io_mem_cluster_29_addr = MAT_io_mem_cluster_29_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_30_en = MAT_io_mem_cluster_30_en; // @[processor.scala 22:24]
  assign io_mem_cluster_30_addr = MAT_io_mem_cluster_30_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_31_en = MAT_io_mem_cluster_31_en; // @[processor.scala 22:24]
  assign io_mem_cluster_31_addr = MAT_io_mem_cluster_31_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_32_en = MAT_io_mem_cluster_32_en; // @[processor.scala 22:24]
  assign io_mem_cluster_32_addr = MAT_io_mem_cluster_32_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_33_en = MAT_io_mem_cluster_33_en; // @[processor.scala 22:24]
  assign io_mem_cluster_33_addr = MAT_io_mem_cluster_33_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_34_en = MAT_io_mem_cluster_34_en; // @[processor.scala 22:24]
  assign io_mem_cluster_34_addr = MAT_io_mem_cluster_34_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_35_en = MAT_io_mem_cluster_35_en; // @[processor.scala 22:24]
  assign io_mem_cluster_35_addr = MAT_io_mem_cluster_35_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_36_en = MAT_io_mem_cluster_36_en; // @[processor.scala 22:24]
  assign io_mem_cluster_36_addr = MAT_io_mem_cluster_36_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_37_en = MAT_io_mem_cluster_37_en; // @[processor.scala 22:24]
  assign io_mem_cluster_37_addr = MAT_io_mem_cluster_37_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_38_en = MAT_io_mem_cluster_38_en; // @[processor.scala 22:24]
  assign io_mem_cluster_38_addr = MAT_io_mem_cluster_38_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_39_en = MAT_io_mem_cluster_39_en; // @[processor.scala 22:24]
  assign io_mem_cluster_39_addr = MAT_io_mem_cluster_39_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_40_en = MAT_io_mem_cluster_40_en; // @[processor.scala 22:24]
  assign io_mem_cluster_40_addr = MAT_io_mem_cluster_40_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_41_en = MAT_io_mem_cluster_41_en; // @[processor.scala 22:24]
  assign io_mem_cluster_41_addr = MAT_io_mem_cluster_41_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_42_en = MAT_io_mem_cluster_42_en; // @[processor.scala 22:24]
  assign io_mem_cluster_42_addr = MAT_io_mem_cluster_42_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_43_en = MAT_io_mem_cluster_43_en; // @[processor.scala 22:24]
  assign io_mem_cluster_43_addr = MAT_io_mem_cluster_43_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_44_en = MAT_io_mem_cluster_44_en; // @[processor.scala 22:24]
  assign io_mem_cluster_44_addr = MAT_io_mem_cluster_44_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_45_en = MAT_io_mem_cluster_45_en; // @[processor.scala 22:24]
  assign io_mem_cluster_45_addr = MAT_io_mem_cluster_45_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_46_en = MAT_io_mem_cluster_46_en; // @[processor.scala 22:24]
  assign io_mem_cluster_46_addr = MAT_io_mem_cluster_46_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_47_en = MAT_io_mem_cluster_47_en; // @[processor.scala 22:24]
  assign io_mem_cluster_47_addr = MAT_io_mem_cluster_47_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_48_en = MAT_io_mem_cluster_48_en; // @[processor.scala 22:24]
  assign io_mem_cluster_48_addr = MAT_io_mem_cluster_48_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_49_en = MAT_io_mem_cluster_49_en; // @[processor.scala 22:24]
  assign io_mem_cluster_49_addr = MAT_io_mem_cluster_49_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_50_en = MAT_io_mem_cluster_50_en; // @[processor.scala 22:24]
  assign io_mem_cluster_50_addr = MAT_io_mem_cluster_50_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_51_en = MAT_io_mem_cluster_51_en; // @[processor.scala 22:24]
  assign io_mem_cluster_51_addr = MAT_io_mem_cluster_51_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_52_en = MAT_io_mem_cluster_52_en; // @[processor.scala 22:24]
  assign io_mem_cluster_52_addr = MAT_io_mem_cluster_52_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_53_en = MAT_io_mem_cluster_53_en; // @[processor.scala 22:24]
  assign io_mem_cluster_53_addr = MAT_io_mem_cluster_53_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_54_en = MAT_io_mem_cluster_54_en; // @[processor.scala 22:24]
  assign io_mem_cluster_54_addr = MAT_io_mem_cluster_54_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_55_en = MAT_io_mem_cluster_55_en; // @[processor.scala 22:24]
  assign io_mem_cluster_55_addr = MAT_io_mem_cluster_55_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_56_en = MAT_io_mem_cluster_56_en; // @[processor.scala 22:24]
  assign io_mem_cluster_56_addr = MAT_io_mem_cluster_56_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_57_en = MAT_io_mem_cluster_57_en; // @[processor.scala 22:24]
  assign io_mem_cluster_57_addr = MAT_io_mem_cluster_57_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_58_en = MAT_io_mem_cluster_58_en; // @[processor.scala 22:24]
  assign io_mem_cluster_58_addr = MAT_io_mem_cluster_58_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_59_en = MAT_io_mem_cluster_59_en; // @[processor.scala 22:24]
  assign io_mem_cluster_59_addr = MAT_io_mem_cluster_59_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_60_en = MAT_io_mem_cluster_60_en; // @[processor.scala 22:24]
  assign io_mem_cluster_60_addr = MAT_io_mem_cluster_60_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_61_en = MAT_io_mem_cluster_61_en; // @[processor.scala 22:24]
  assign io_mem_cluster_61_addr = MAT_io_mem_cluster_61_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_62_en = MAT_io_mem_cluster_62_en; // @[processor.scala 22:24]
  assign io_mem_cluster_62_addr = MAT_io_mem_cluster_62_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_63_en = MAT_io_mem_cluster_63_en; // @[processor.scala 22:24]
  assign io_mem_cluster_63_addr = MAT_io_mem_cluster_63_addr; // @[processor.scala 22:24]
  assign PAR_clock = clock;
  assign PAR_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_96 = io_pipe_phv_in_data_96; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_97 = io_pipe_phv_in_data_97; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_98 = io_pipe_phv_in_data_98; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_99 = io_pipe_phv_in_data_99; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_100 = io_pipe_phv_in_data_100; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_101 = io_pipe_phv_in_data_101; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_102 = io_pipe_phv_in_data_102; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_103 = io_pipe_phv_in_data_103; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_104 = io_pipe_phv_in_data_104; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_105 = io_pipe_phv_in_data_105; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_106 = io_pipe_phv_in_data_106; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_107 = io_pipe_phv_in_data_107; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_108 = io_pipe_phv_in_data_108; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_109 = io_pipe_phv_in_data_109; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_110 = io_pipe_phv_in_data_110; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_111 = io_pipe_phv_in_data_111; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_112 = io_pipe_phv_in_data_112; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_113 = io_pipe_phv_in_data_113; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_114 = io_pipe_phv_in_data_114; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_115 = io_pipe_phv_in_data_115; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_116 = io_pipe_phv_in_data_116; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_117 = io_pipe_phv_in_data_117; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_118 = io_pipe_phv_in_data_118; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_119 = io_pipe_phv_in_data_119; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_120 = io_pipe_phv_in_data_120; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_121 = io_pipe_phv_in_data_121; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_122 = io_pipe_phv_in_data_122; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_123 = io_pipe_phv_in_data_123; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_124 = io_pipe_phv_in_data_124; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_125 = io_pipe_phv_in_data_125; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_126 = io_pipe_phv_in_data_126; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_127 = io_pipe_phv_in_data_127; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_128 = io_pipe_phv_in_data_128; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_129 = io_pipe_phv_in_data_129; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_130 = io_pipe_phv_in_data_130; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_131 = io_pipe_phv_in_data_131; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_132 = io_pipe_phv_in_data_132; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_133 = io_pipe_phv_in_data_133; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_134 = io_pipe_phv_in_data_134; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_135 = io_pipe_phv_in_data_135; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_136 = io_pipe_phv_in_data_136; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_137 = io_pipe_phv_in_data_137; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_138 = io_pipe_phv_in_data_138; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_139 = io_pipe_phv_in_data_139; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_140 = io_pipe_phv_in_data_140; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_141 = io_pipe_phv_in_data_141; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_142 = io_pipe_phv_in_data_142; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_143 = io_pipe_phv_in_data_143; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_144 = io_pipe_phv_in_data_144; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_145 = io_pipe_phv_in_data_145; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_146 = io_pipe_phv_in_data_146; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_147 = io_pipe_phv_in_data_147; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_148 = io_pipe_phv_in_data_148; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_149 = io_pipe_phv_in_data_149; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_150 = io_pipe_phv_in_data_150; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_151 = io_pipe_phv_in_data_151; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_152 = io_pipe_phv_in_data_152; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_153 = io_pipe_phv_in_data_153; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_154 = io_pipe_phv_in_data_154; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_155 = io_pipe_phv_in_data_155; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_156 = io_pipe_phv_in_data_156; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_157 = io_pipe_phv_in_data_157; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_158 = io_pipe_phv_in_data_158; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_159 = io_pipe_phv_in_data_159; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_160 = io_pipe_phv_in_data_160; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_161 = io_pipe_phv_in_data_161; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_162 = io_pipe_phv_in_data_162; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_163 = io_pipe_phv_in_data_163; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_164 = io_pipe_phv_in_data_164; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_165 = io_pipe_phv_in_data_165; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_166 = io_pipe_phv_in_data_166; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_167 = io_pipe_phv_in_data_167; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_168 = io_pipe_phv_in_data_168; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_169 = io_pipe_phv_in_data_169; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_170 = io_pipe_phv_in_data_170; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_171 = io_pipe_phv_in_data_171; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_172 = io_pipe_phv_in_data_172; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_173 = io_pipe_phv_in_data_173; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_174 = io_pipe_phv_in_data_174; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_175 = io_pipe_phv_in_data_175; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_176 = io_pipe_phv_in_data_176; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_177 = io_pipe_phv_in_data_177; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_178 = io_pipe_phv_in_data_178; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_179 = io_pipe_phv_in_data_179; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_180 = io_pipe_phv_in_data_180; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_181 = io_pipe_phv_in_data_181; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_182 = io_pipe_phv_in_data_182; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_183 = io_pipe_phv_in_data_183; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_184 = io_pipe_phv_in_data_184; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_185 = io_pipe_phv_in_data_185; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_186 = io_pipe_phv_in_data_186; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_187 = io_pipe_phv_in_data_187; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_188 = io_pipe_phv_in_data_188; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_189 = io_pipe_phv_in_data_189; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_190 = io_pipe_phv_in_data_190; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_191 = io_pipe_phv_in_data_191; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_192 = io_pipe_phv_in_data_192; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_193 = io_pipe_phv_in_data_193; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_194 = io_pipe_phv_in_data_194; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_195 = io_pipe_phv_in_data_195; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_196 = io_pipe_phv_in_data_196; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_197 = io_pipe_phv_in_data_197; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_198 = io_pipe_phv_in_data_198; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_199 = io_pipe_phv_in_data_199; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_200 = io_pipe_phv_in_data_200; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_201 = io_pipe_phv_in_data_201; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_202 = io_pipe_phv_in_data_202; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_203 = io_pipe_phv_in_data_203; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_204 = io_pipe_phv_in_data_204; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_205 = io_pipe_phv_in_data_205; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_206 = io_pipe_phv_in_data_206; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_207 = io_pipe_phv_in_data_207; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_208 = io_pipe_phv_in_data_208; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_209 = io_pipe_phv_in_data_209; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_210 = io_pipe_phv_in_data_210; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_211 = io_pipe_phv_in_data_211; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_212 = io_pipe_phv_in_data_212; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_213 = io_pipe_phv_in_data_213; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_214 = io_pipe_phv_in_data_214; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_215 = io_pipe_phv_in_data_215; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_216 = io_pipe_phv_in_data_216; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_217 = io_pipe_phv_in_data_217; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_218 = io_pipe_phv_in_data_218; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_219 = io_pipe_phv_in_data_219; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_220 = io_pipe_phv_in_data_220; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_221 = io_pipe_phv_in_data_221; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_222 = io_pipe_phv_in_data_222; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_223 = io_pipe_phv_in_data_223; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_224 = io_pipe_phv_in_data_224; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_225 = io_pipe_phv_in_data_225; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_226 = io_pipe_phv_in_data_226; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_227 = io_pipe_phv_in_data_227; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_228 = io_pipe_phv_in_data_228; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_229 = io_pipe_phv_in_data_229; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_230 = io_pipe_phv_in_data_230; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_231 = io_pipe_phv_in_data_231; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_232 = io_pipe_phv_in_data_232; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_233 = io_pipe_phv_in_data_233; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_234 = io_pipe_phv_in_data_234; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_235 = io_pipe_phv_in_data_235; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_236 = io_pipe_phv_in_data_236; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_237 = io_pipe_phv_in_data_237; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_238 = io_pipe_phv_in_data_238; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_239 = io_pipe_phv_in_data_239; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_240 = io_pipe_phv_in_data_240; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_241 = io_pipe_phv_in_data_241; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_242 = io_pipe_phv_in_data_242; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_243 = io_pipe_phv_in_data_243; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_244 = io_pipe_phv_in_data_244; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_245 = io_pipe_phv_in_data_245; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_246 = io_pipe_phv_in_data_246; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_247 = io_pipe_phv_in_data_247; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_248 = io_pipe_phv_in_data_248; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_249 = io_pipe_phv_in_data_249; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_250 = io_pipe_phv_in_data_250; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_251 = io_pipe_phv_in_data_251; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_252 = io_pipe_phv_in_data_252; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_253 = io_pipe_phv_in_data_253; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_254 = io_pipe_phv_in_data_254; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_255 = io_pipe_phv_in_data_255; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_0 = io_pipe_phv_in_header_0; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_1 = io_pipe_phv_in_header_1; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_2 = io_pipe_phv_in_header_2; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_3 = io_pipe_phv_in_header_3; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_4 = io_pipe_phv_in_header_4; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_5 = io_pipe_phv_in_header_5; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_6 = io_pipe_phv_in_header_6; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_7 = io_pipe_phv_in_header_7; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_8 = io_pipe_phv_in_header_8; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_9 = io_pipe_phv_in_header_9; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_10 = io_pipe_phv_in_header_10; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_11 = io_pipe_phv_in_header_11; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_12 = io_pipe_phv_in_header_12; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_13 = io_pipe_phv_in_header_13; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_14 = io_pipe_phv_in_header_14; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_15 = io_pipe_phv_in_header_15; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_parse_current_state = io_pipe_phv_in_parse_current_state; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_parse_current_offset = io_pipe_phv_in_parse_current_offset; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_parse_transition_field = io_pipe_phv_in_parse_transition_field; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_next_processor_id = io_pipe_phv_in_next_processor_id; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_next_config_id = io_pipe_phv_in_next_config_id; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_is_valid_processor = io_pipe_phv_in_is_valid_processor; // @[processor.scala 17:24]
  assign PAR_io_mod_en = io_mod_par_mod_en; // @[processor.scala 18:24]
  assign PAR_io_mod_last_mau_id_mod = io_mod_par_mod_last_mau_id_mod; // @[processor.scala 18:24]
  assign PAR_io_mod_last_mau_id = io_mod_par_mod_last_mau_id; // @[processor.scala 18:24]
  assign PAR_io_mod_cs = io_mod_par_mod_cs; // @[processor.scala 18:24]
  assign PAR_io_mod_module_mod_state_id_mod = io_mod_par_mod_module_mod_state_id_mod; // @[processor.scala 18:24]
  assign PAR_io_mod_module_mod_state_id = io_mod_par_mod_module_mod_state_id; // @[processor.scala 18:24]
  assign PAR_io_mod_module_mod_sram_w_cs = io_mod_par_mod_module_mod_sram_w_cs; // @[processor.scala 18:24]
  assign PAR_io_mod_module_mod_sram_w_en = io_mod_par_mod_module_mod_sram_w_en; // @[processor.scala 18:24]
  assign PAR_io_mod_module_mod_sram_w_addr = io_mod_par_mod_module_mod_sram_w_addr; // @[processor.scala 18:24]
  assign PAR_io_mod_module_mod_sram_w_data = io_mod_par_mod_module_mod_sram_w_data; // @[processor.scala 18:24]
  assign MAT_clock = clock;
  assign MAT_io_pipe_phv_in_data_0 = PAR_io_pipe_phv_out_data_0; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_1 = PAR_io_pipe_phv_out_data_1; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_2 = PAR_io_pipe_phv_out_data_2; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_3 = PAR_io_pipe_phv_out_data_3; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_4 = PAR_io_pipe_phv_out_data_4; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_5 = PAR_io_pipe_phv_out_data_5; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_6 = PAR_io_pipe_phv_out_data_6; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_7 = PAR_io_pipe_phv_out_data_7; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_8 = PAR_io_pipe_phv_out_data_8; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_9 = PAR_io_pipe_phv_out_data_9; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_10 = PAR_io_pipe_phv_out_data_10; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_11 = PAR_io_pipe_phv_out_data_11; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_12 = PAR_io_pipe_phv_out_data_12; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_13 = PAR_io_pipe_phv_out_data_13; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_14 = PAR_io_pipe_phv_out_data_14; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_15 = PAR_io_pipe_phv_out_data_15; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_16 = PAR_io_pipe_phv_out_data_16; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_17 = PAR_io_pipe_phv_out_data_17; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_18 = PAR_io_pipe_phv_out_data_18; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_19 = PAR_io_pipe_phv_out_data_19; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_20 = PAR_io_pipe_phv_out_data_20; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_21 = PAR_io_pipe_phv_out_data_21; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_22 = PAR_io_pipe_phv_out_data_22; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_23 = PAR_io_pipe_phv_out_data_23; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_24 = PAR_io_pipe_phv_out_data_24; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_25 = PAR_io_pipe_phv_out_data_25; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_26 = PAR_io_pipe_phv_out_data_26; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_27 = PAR_io_pipe_phv_out_data_27; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_28 = PAR_io_pipe_phv_out_data_28; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_29 = PAR_io_pipe_phv_out_data_29; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_30 = PAR_io_pipe_phv_out_data_30; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_31 = PAR_io_pipe_phv_out_data_31; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_32 = PAR_io_pipe_phv_out_data_32; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_33 = PAR_io_pipe_phv_out_data_33; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_34 = PAR_io_pipe_phv_out_data_34; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_35 = PAR_io_pipe_phv_out_data_35; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_36 = PAR_io_pipe_phv_out_data_36; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_37 = PAR_io_pipe_phv_out_data_37; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_38 = PAR_io_pipe_phv_out_data_38; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_39 = PAR_io_pipe_phv_out_data_39; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_40 = PAR_io_pipe_phv_out_data_40; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_41 = PAR_io_pipe_phv_out_data_41; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_42 = PAR_io_pipe_phv_out_data_42; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_43 = PAR_io_pipe_phv_out_data_43; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_44 = PAR_io_pipe_phv_out_data_44; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_45 = PAR_io_pipe_phv_out_data_45; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_46 = PAR_io_pipe_phv_out_data_46; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_47 = PAR_io_pipe_phv_out_data_47; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_48 = PAR_io_pipe_phv_out_data_48; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_49 = PAR_io_pipe_phv_out_data_49; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_50 = PAR_io_pipe_phv_out_data_50; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_51 = PAR_io_pipe_phv_out_data_51; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_52 = PAR_io_pipe_phv_out_data_52; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_53 = PAR_io_pipe_phv_out_data_53; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_54 = PAR_io_pipe_phv_out_data_54; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_55 = PAR_io_pipe_phv_out_data_55; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_56 = PAR_io_pipe_phv_out_data_56; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_57 = PAR_io_pipe_phv_out_data_57; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_58 = PAR_io_pipe_phv_out_data_58; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_59 = PAR_io_pipe_phv_out_data_59; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_60 = PAR_io_pipe_phv_out_data_60; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_61 = PAR_io_pipe_phv_out_data_61; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_62 = PAR_io_pipe_phv_out_data_62; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_63 = PAR_io_pipe_phv_out_data_63; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_64 = PAR_io_pipe_phv_out_data_64; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_65 = PAR_io_pipe_phv_out_data_65; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_66 = PAR_io_pipe_phv_out_data_66; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_67 = PAR_io_pipe_phv_out_data_67; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_68 = PAR_io_pipe_phv_out_data_68; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_69 = PAR_io_pipe_phv_out_data_69; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_70 = PAR_io_pipe_phv_out_data_70; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_71 = PAR_io_pipe_phv_out_data_71; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_72 = PAR_io_pipe_phv_out_data_72; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_73 = PAR_io_pipe_phv_out_data_73; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_74 = PAR_io_pipe_phv_out_data_74; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_75 = PAR_io_pipe_phv_out_data_75; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_76 = PAR_io_pipe_phv_out_data_76; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_77 = PAR_io_pipe_phv_out_data_77; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_78 = PAR_io_pipe_phv_out_data_78; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_79 = PAR_io_pipe_phv_out_data_79; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_80 = PAR_io_pipe_phv_out_data_80; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_81 = PAR_io_pipe_phv_out_data_81; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_82 = PAR_io_pipe_phv_out_data_82; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_83 = PAR_io_pipe_phv_out_data_83; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_84 = PAR_io_pipe_phv_out_data_84; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_85 = PAR_io_pipe_phv_out_data_85; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_86 = PAR_io_pipe_phv_out_data_86; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_87 = PAR_io_pipe_phv_out_data_87; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_88 = PAR_io_pipe_phv_out_data_88; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_89 = PAR_io_pipe_phv_out_data_89; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_90 = PAR_io_pipe_phv_out_data_90; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_91 = PAR_io_pipe_phv_out_data_91; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_92 = PAR_io_pipe_phv_out_data_92; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_93 = PAR_io_pipe_phv_out_data_93; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_94 = PAR_io_pipe_phv_out_data_94; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_95 = PAR_io_pipe_phv_out_data_95; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_96 = PAR_io_pipe_phv_out_data_96; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_97 = PAR_io_pipe_phv_out_data_97; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_98 = PAR_io_pipe_phv_out_data_98; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_99 = PAR_io_pipe_phv_out_data_99; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_100 = PAR_io_pipe_phv_out_data_100; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_101 = PAR_io_pipe_phv_out_data_101; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_102 = PAR_io_pipe_phv_out_data_102; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_103 = PAR_io_pipe_phv_out_data_103; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_104 = PAR_io_pipe_phv_out_data_104; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_105 = PAR_io_pipe_phv_out_data_105; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_106 = PAR_io_pipe_phv_out_data_106; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_107 = PAR_io_pipe_phv_out_data_107; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_108 = PAR_io_pipe_phv_out_data_108; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_109 = PAR_io_pipe_phv_out_data_109; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_110 = PAR_io_pipe_phv_out_data_110; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_111 = PAR_io_pipe_phv_out_data_111; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_112 = PAR_io_pipe_phv_out_data_112; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_113 = PAR_io_pipe_phv_out_data_113; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_114 = PAR_io_pipe_phv_out_data_114; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_115 = PAR_io_pipe_phv_out_data_115; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_116 = PAR_io_pipe_phv_out_data_116; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_117 = PAR_io_pipe_phv_out_data_117; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_118 = PAR_io_pipe_phv_out_data_118; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_119 = PAR_io_pipe_phv_out_data_119; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_120 = PAR_io_pipe_phv_out_data_120; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_121 = PAR_io_pipe_phv_out_data_121; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_122 = PAR_io_pipe_phv_out_data_122; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_123 = PAR_io_pipe_phv_out_data_123; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_124 = PAR_io_pipe_phv_out_data_124; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_125 = PAR_io_pipe_phv_out_data_125; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_126 = PAR_io_pipe_phv_out_data_126; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_127 = PAR_io_pipe_phv_out_data_127; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_128 = PAR_io_pipe_phv_out_data_128; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_129 = PAR_io_pipe_phv_out_data_129; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_130 = PAR_io_pipe_phv_out_data_130; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_131 = PAR_io_pipe_phv_out_data_131; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_132 = PAR_io_pipe_phv_out_data_132; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_133 = PAR_io_pipe_phv_out_data_133; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_134 = PAR_io_pipe_phv_out_data_134; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_135 = PAR_io_pipe_phv_out_data_135; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_136 = PAR_io_pipe_phv_out_data_136; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_137 = PAR_io_pipe_phv_out_data_137; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_138 = PAR_io_pipe_phv_out_data_138; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_139 = PAR_io_pipe_phv_out_data_139; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_140 = PAR_io_pipe_phv_out_data_140; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_141 = PAR_io_pipe_phv_out_data_141; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_142 = PAR_io_pipe_phv_out_data_142; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_143 = PAR_io_pipe_phv_out_data_143; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_144 = PAR_io_pipe_phv_out_data_144; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_145 = PAR_io_pipe_phv_out_data_145; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_146 = PAR_io_pipe_phv_out_data_146; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_147 = PAR_io_pipe_phv_out_data_147; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_148 = PAR_io_pipe_phv_out_data_148; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_149 = PAR_io_pipe_phv_out_data_149; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_150 = PAR_io_pipe_phv_out_data_150; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_151 = PAR_io_pipe_phv_out_data_151; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_152 = PAR_io_pipe_phv_out_data_152; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_153 = PAR_io_pipe_phv_out_data_153; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_154 = PAR_io_pipe_phv_out_data_154; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_155 = PAR_io_pipe_phv_out_data_155; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_156 = PAR_io_pipe_phv_out_data_156; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_157 = PAR_io_pipe_phv_out_data_157; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_158 = PAR_io_pipe_phv_out_data_158; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_159 = PAR_io_pipe_phv_out_data_159; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_160 = PAR_io_pipe_phv_out_data_160; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_161 = PAR_io_pipe_phv_out_data_161; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_162 = PAR_io_pipe_phv_out_data_162; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_163 = PAR_io_pipe_phv_out_data_163; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_164 = PAR_io_pipe_phv_out_data_164; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_165 = PAR_io_pipe_phv_out_data_165; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_166 = PAR_io_pipe_phv_out_data_166; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_167 = PAR_io_pipe_phv_out_data_167; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_168 = PAR_io_pipe_phv_out_data_168; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_169 = PAR_io_pipe_phv_out_data_169; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_170 = PAR_io_pipe_phv_out_data_170; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_171 = PAR_io_pipe_phv_out_data_171; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_172 = PAR_io_pipe_phv_out_data_172; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_173 = PAR_io_pipe_phv_out_data_173; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_174 = PAR_io_pipe_phv_out_data_174; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_175 = PAR_io_pipe_phv_out_data_175; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_176 = PAR_io_pipe_phv_out_data_176; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_177 = PAR_io_pipe_phv_out_data_177; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_178 = PAR_io_pipe_phv_out_data_178; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_179 = PAR_io_pipe_phv_out_data_179; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_180 = PAR_io_pipe_phv_out_data_180; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_181 = PAR_io_pipe_phv_out_data_181; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_182 = PAR_io_pipe_phv_out_data_182; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_183 = PAR_io_pipe_phv_out_data_183; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_184 = PAR_io_pipe_phv_out_data_184; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_185 = PAR_io_pipe_phv_out_data_185; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_186 = PAR_io_pipe_phv_out_data_186; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_187 = PAR_io_pipe_phv_out_data_187; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_188 = PAR_io_pipe_phv_out_data_188; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_189 = PAR_io_pipe_phv_out_data_189; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_190 = PAR_io_pipe_phv_out_data_190; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_191 = PAR_io_pipe_phv_out_data_191; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_192 = PAR_io_pipe_phv_out_data_192; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_193 = PAR_io_pipe_phv_out_data_193; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_194 = PAR_io_pipe_phv_out_data_194; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_195 = PAR_io_pipe_phv_out_data_195; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_196 = PAR_io_pipe_phv_out_data_196; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_197 = PAR_io_pipe_phv_out_data_197; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_198 = PAR_io_pipe_phv_out_data_198; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_199 = PAR_io_pipe_phv_out_data_199; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_200 = PAR_io_pipe_phv_out_data_200; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_201 = PAR_io_pipe_phv_out_data_201; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_202 = PAR_io_pipe_phv_out_data_202; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_203 = PAR_io_pipe_phv_out_data_203; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_204 = PAR_io_pipe_phv_out_data_204; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_205 = PAR_io_pipe_phv_out_data_205; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_206 = PAR_io_pipe_phv_out_data_206; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_207 = PAR_io_pipe_phv_out_data_207; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_208 = PAR_io_pipe_phv_out_data_208; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_209 = PAR_io_pipe_phv_out_data_209; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_210 = PAR_io_pipe_phv_out_data_210; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_211 = PAR_io_pipe_phv_out_data_211; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_212 = PAR_io_pipe_phv_out_data_212; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_213 = PAR_io_pipe_phv_out_data_213; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_214 = PAR_io_pipe_phv_out_data_214; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_215 = PAR_io_pipe_phv_out_data_215; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_216 = PAR_io_pipe_phv_out_data_216; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_217 = PAR_io_pipe_phv_out_data_217; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_218 = PAR_io_pipe_phv_out_data_218; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_219 = PAR_io_pipe_phv_out_data_219; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_220 = PAR_io_pipe_phv_out_data_220; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_221 = PAR_io_pipe_phv_out_data_221; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_222 = PAR_io_pipe_phv_out_data_222; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_223 = PAR_io_pipe_phv_out_data_223; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_224 = PAR_io_pipe_phv_out_data_224; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_225 = PAR_io_pipe_phv_out_data_225; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_226 = PAR_io_pipe_phv_out_data_226; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_227 = PAR_io_pipe_phv_out_data_227; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_228 = PAR_io_pipe_phv_out_data_228; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_229 = PAR_io_pipe_phv_out_data_229; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_230 = PAR_io_pipe_phv_out_data_230; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_231 = PAR_io_pipe_phv_out_data_231; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_232 = PAR_io_pipe_phv_out_data_232; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_233 = PAR_io_pipe_phv_out_data_233; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_234 = PAR_io_pipe_phv_out_data_234; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_235 = PAR_io_pipe_phv_out_data_235; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_236 = PAR_io_pipe_phv_out_data_236; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_237 = PAR_io_pipe_phv_out_data_237; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_238 = PAR_io_pipe_phv_out_data_238; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_239 = PAR_io_pipe_phv_out_data_239; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_240 = PAR_io_pipe_phv_out_data_240; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_241 = PAR_io_pipe_phv_out_data_241; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_242 = PAR_io_pipe_phv_out_data_242; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_243 = PAR_io_pipe_phv_out_data_243; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_244 = PAR_io_pipe_phv_out_data_244; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_245 = PAR_io_pipe_phv_out_data_245; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_246 = PAR_io_pipe_phv_out_data_246; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_247 = PAR_io_pipe_phv_out_data_247; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_248 = PAR_io_pipe_phv_out_data_248; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_249 = PAR_io_pipe_phv_out_data_249; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_250 = PAR_io_pipe_phv_out_data_250; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_251 = PAR_io_pipe_phv_out_data_251; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_252 = PAR_io_pipe_phv_out_data_252; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_253 = PAR_io_pipe_phv_out_data_253; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_254 = PAR_io_pipe_phv_out_data_254; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_255 = PAR_io_pipe_phv_out_data_255; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_0 = PAR_io_pipe_phv_out_header_0; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_1 = PAR_io_pipe_phv_out_header_1; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_2 = PAR_io_pipe_phv_out_header_2; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_3 = PAR_io_pipe_phv_out_header_3; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_4 = PAR_io_pipe_phv_out_header_4; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_5 = PAR_io_pipe_phv_out_header_5; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_6 = PAR_io_pipe_phv_out_header_6; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_7 = PAR_io_pipe_phv_out_header_7; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_8 = PAR_io_pipe_phv_out_header_8; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_9 = PAR_io_pipe_phv_out_header_9; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_10 = PAR_io_pipe_phv_out_header_10; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_11 = PAR_io_pipe_phv_out_header_11; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_12 = PAR_io_pipe_phv_out_header_12; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_13 = PAR_io_pipe_phv_out_header_13; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_14 = PAR_io_pipe_phv_out_header_14; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_15 = PAR_io_pipe_phv_out_header_15; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_parse_current_state = PAR_io_pipe_phv_out_parse_current_state; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_parse_current_offset = PAR_io_pipe_phv_out_parse_current_offset; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_parse_transition_field = PAR_io_pipe_phv_out_parse_transition_field; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_next_processor_id = PAR_io_pipe_phv_out_next_processor_id; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_next_config_id = PAR_io_pipe_phv_out_next_config_id; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_is_valid_processor = PAR_io_pipe_phv_out_is_valid_processor; // @[processor.scala 20:24]
  assign MAT_io_mod_en = io_mod_mat_mod_en; // @[processor.scala 21:24]
  assign MAT_io_mod_config_id = io_mod_mat_mod_config_id; // @[processor.scala 21:24]
  assign MAT_io_mod_key_mod_header_id = io_mod_mat_mod_key_mod_header_id; // @[processor.scala 21:24]
  assign MAT_io_mod_key_mod_internal_offset = io_mod_mat_mod_key_mod_internal_offset; // @[processor.scala 21:24]
  assign MAT_io_mod_key_mod_key_length = io_mod_mat_mod_key_mod_key_length; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_0 = io_mod_mat_mod_table_mod_sram_id_table_0; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_1 = io_mod_mat_mod_table_mod_sram_id_table_1; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_2 = io_mod_mat_mod_table_mod_sram_id_table_2; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_3 = io_mod_mat_mod_table_mod_sram_id_table_3; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_4 = io_mod_mat_mod_table_mod_sram_id_table_4; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_5 = io_mod_mat_mod_table_mod_sram_id_table_5; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_6 = io_mod_mat_mod_table_mod_sram_id_table_6; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_7 = io_mod_mat_mod_table_mod_sram_id_table_7; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_8 = io_mod_mat_mod_table_mod_sram_id_table_8; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_9 = io_mod_mat_mod_table_mod_sram_id_table_9; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_10 = io_mod_mat_mod_table_mod_sram_id_table_10; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_11 = io_mod_mat_mod_table_mod_sram_id_table_11; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_12 = io_mod_mat_mod_table_mod_sram_id_table_12; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_13 = io_mod_mat_mod_table_mod_sram_id_table_13; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_14 = io_mod_mat_mod_table_mod_sram_id_table_14; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_15 = io_mod_mat_mod_table_mod_sram_id_table_15; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_16 = io_mod_mat_mod_table_mod_sram_id_table_16; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_17 = io_mod_mat_mod_table_mod_sram_id_table_17; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_18 = io_mod_mat_mod_table_mod_sram_id_table_18; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_19 = io_mod_mat_mod_table_mod_sram_id_table_19; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_20 = io_mod_mat_mod_table_mod_sram_id_table_20; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_21 = io_mod_mat_mod_table_mod_sram_id_table_21; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_22 = io_mod_mat_mod_table_mod_sram_id_table_22; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_23 = io_mod_mat_mod_table_mod_sram_id_table_23; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_24 = io_mod_mat_mod_table_mod_sram_id_table_24; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_25 = io_mod_mat_mod_table_mod_sram_id_table_25; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_26 = io_mod_mat_mod_table_mod_sram_id_table_26; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_27 = io_mod_mat_mod_table_mod_sram_id_table_27; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_28 = io_mod_mat_mod_table_mod_sram_id_table_28; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_29 = io_mod_mat_mod_table_mod_sram_id_table_29; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_30 = io_mod_mat_mod_table_mod_sram_id_table_30; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_31 = io_mod_mat_mod_table_mod_sram_id_table_31; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_32 = io_mod_mat_mod_table_mod_sram_id_table_32; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_33 = io_mod_mat_mod_table_mod_sram_id_table_33; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_34 = io_mod_mat_mod_table_mod_sram_id_table_34; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_35 = io_mod_mat_mod_table_mod_sram_id_table_35; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_36 = io_mod_mat_mod_table_mod_sram_id_table_36; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_37 = io_mod_mat_mod_table_mod_sram_id_table_37; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_38 = io_mod_mat_mod_table_mod_sram_id_table_38; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_39 = io_mod_mat_mod_table_mod_sram_id_table_39; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_40 = io_mod_mat_mod_table_mod_sram_id_table_40; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_41 = io_mod_mat_mod_table_mod_sram_id_table_41; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_42 = io_mod_mat_mod_table_mod_sram_id_table_42; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_43 = io_mod_mat_mod_table_mod_sram_id_table_43; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_44 = io_mod_mat_mod_table_mod_sram_id_table_44; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_45 = io_mod_mat_mod_table_mod_sram_id_table_45; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_46 = io_mod_mat_mod_table_mod_sram_id_table_46; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_47 = io_mod_mat_mod_table_mod_sram_id_table_47; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_48 = io_mod_mat_mod_table_mod_sram_id_table_48; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_49 = io_mod_mat_mod_table_mod_sram_id_table_49; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_50 = io_mod_mat_mod_table_mod_sram_id_table_50; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_51 = io_mod_mat_mod_table_mod_sram_id_table_51; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_52 = io_mod_mat_mod_table_mod_sram_id_table_52; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_53 = io_mod_mat_mod_table_mod_sram_id_table_53; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_54 = io_mod_mat_mod_table_mod_sram_id_table_54; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_55 = io_mod_mat_mod_table_mod_sram_id_table_55; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_56 = io_mod_mat_mod_table_mod_sram_id_table_56; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_57 = io_mod_mat_mod_table_mod_sram_id_table_57; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_58 = io_mod_mat_mod_table_mod_sram_id_table_58; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_59 = io_mod_mat_mod_table_mod_sram_id_table_59; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_60 = io_mod_mat_mod_table_mod_sram_id_table_60; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_61 = io_mod_mat_mod_table_mod_sram_id_table_61; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_62 = io_mod_mat_mod_table_mod_sram_id_table_62; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_sram_id_table_63 = io_mod_mat_mod_table_mod_sram_id_table_63; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_table_width = io_mod_mat_mod_table_mod_table_width; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_table_depth = io_mod_mat_mod_table_mod_table_depth; // @[processor.scala 21:24]
  assign MAT_io_mem_cluster_0_data = io_mem_cluster_0_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_1_data = io_mem_cluster_1_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_2_data = io_mem_cluster_2_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_3_data = io_mem_cluster_3_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_4_data = io_mem_cluster_4_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_5_data = io_mem_cluster_5_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_6_data = io_mem_cluster_6_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_7_data = io_mem_cluster_7_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_8_data = io_mem_cluster_8_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_9_data = io_mem_cluster_9_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_10_data = io_mem_cluster_10_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_11_data = io_mem_cluster_11_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_12_data = io_mem_cluster_12_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_13_data = io_mem_cluster_13_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_14_data = io_mem_cluster_14_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_15_data = io_mem_cluster_15_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_16_data = io_mem_cluster_16_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_17_data = io_mem_cluster_17_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_18_data = io_mem_cluster_18_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_19_data = io_mem_cluster_19_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_20_data = io_mem_cluster_20_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_21_data = io_mem_cluster_21_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_22_data = io_mem_cluster_22_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_23_data = io_mem_cluster_23_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_24_data = io_mem_cluster_24_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_25_data = io_mem_cluster_25_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_26_data = io_mem_cluster_26_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_27_data = io_mem_cluster_27_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_28_data = io_mem_cluster_28_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_29_data = io_mem_cluster_29_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_30_data = io_mem_cluster_30_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_31_data = io_mem_cluster_31_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_32_data = io_mem_cluster_32_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_33_data = io_mem_cluster_33_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_34_data = io_mem_cluster_34_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_35_data = io_mem_cluster_35_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_36_data = io_mem_cluster_36_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_37_data = io_mem_cluster_37_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_38_data = io_mem_cluster_38_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_39_data = io_mem_cluster_39_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_40_data = io_mem_cluster_40_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_41_data = io_mem_cluster_41_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_42_data = io_mem_cluster_42_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_43_data = io_mem_cluster_43_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_44_data = io_mem_cluster_44_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_45_data = io_mem_cluster_45_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_46_data = io_mem_cluster_46_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_47_data = io_mem_cluster_47_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_48_data = io_mem_cluster_48_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_49_data = io_mem_cluster_49_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_50_data = io_mem_cluster_50_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_51_data = io_mem_cluster_51_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_52_data = io_mem_cluster_52_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_53_data = io_mem_cluster_53_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_54_data = io_mem_cluster_54_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_55_data = io_mem_cluster_55_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_56_data = io_mem_cluster_56_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_57_data = io_mem_cluster_57_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_58_data = io_mem_cluster_58_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_59_data = io_mem_cluster_59_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_60_data = io_mem_cluster_60_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_61_data = io_mem_cluster_61_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_62_data = io_mem_cluster_62_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_63_data = io_mem_cluster_63_data; // @[processor.scala 22:24]
  assign EXE_clock = clock;
  assign EXE_io_pipe_phv_in_data_0 = MAT_io_pipe_phv_out_data_0; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_1 = MAT_io_pipe_phv_out_data_1; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_2 = MAT_io_pipe_phv_out_data_2; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_3 = MAT_io_pipe_phv_out_data_3; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_4 = MAT_io_pipe_phv_out_data_4; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_5 = MAT_io_pipe_phv_out_data_5; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_6 = MAT_io_pipe_phv_out_data_6; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_7 = MAT_io_pipe_phv_out_data_7; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_8 = MAT_io_pipe_phv_out_data_8; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_9 = MAT_io_pipe_phv_out_data_9; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_10 = MAT_io_pipe_phv_out_data_10; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_11 = MAT_io_pipe_phv_out_data_11; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_12 = MAT_io_pipe_phv_out_data_12; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_13 = MAT_io_pipe_phv_out_data_13; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_14 = MAT_io_pipe_phv_out_data_14; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_15 = MAT_io_pipe_phv_out_data_15; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_16 = MAT_io_pipe_phv_out_data_16; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_17 = MAT_io_pipe_phv_out_data_17; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_18 = MAT_io_pipe_phv_out_data_18; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_19 = MAT_io_pipe_phv_out_data_19; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_20 = MAT_io_pipe_phv_out_data_20; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_21 = MAT_io_pipe_phv_out_data_21; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_22 = MAT_io_pipe_phv_out_data_22; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_23 = MAT_io_pipe_phv_out_data_23; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_24 = MAT_io_pipe_phv_out_data_24; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_25 = MAT_io_pipe_phv_out_data_25; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_26 = MAT_io_pipe_phv_out_data_26; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_27 = MAT_io_pipe_phv_out_data_27; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_28 = MAT_io_pipe_phv_out_data_28; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_29 = MAT_io_pipe_phv_out_data_29; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_30 = MAT_io_pipe_phv_out_data_30; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_31 = MAT_io_pipe_phv_out_data_31; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_32 = MAT_io_pipe_phv_out_data_32; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_33 = MAT_io_pipe_phv_out_data_33; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_34 = MAT_io_pipe_phv_out_data_34; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_35 = MAT_io_pipe_phv_out_data_35; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_36 = MAT_io_pipe_phv_out_data_36; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_37 = MAT_io_pipe_phv_out_data_37; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_38 = MAT_io_pipe_phv_out_data_38; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_39 = MAT_io_pipe_phv_out_data_39; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_40 = MAT_io_pipe_phv_out_data_40; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_41 = MAT_io_pipe_phv_out_data_41; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_42 = MAT_io_pipe_phv_out_data_42; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_43 = MAT_io_pipe_phv_out_data_43; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_44 = MAT_io_pipe_phv_out_data_44; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_45 = MAT_io_pipe_phv_out_data_45; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_46 = MAT_io_pipe_phv_out_data_46; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_47 = MAT_io_pipe_phv_out_data_47; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_48 = MAT_io_pipe_phv_out_data_48; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_49 = MAT_io_pipe_phv_out_data_49; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_50 = MAT_io_pipe_phv_out_data_50; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_51 = MAT_io_pipe_phv_out_data_51; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_52 = MAT_io_pipe_phv_out_data_52; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_53 = MAT_io_pipe_phv_out_data_53; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_54 = MAT_io_pipe_phv_out_data_54; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_55 = MAT_io_pipe_phv_out_data_55; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_56 = MAT_io_pipe_phv_out_data_56; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_57 = MAT_io_pipe_phv_out_data_57; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_58 = MAT_io_pipe_phv_out_data_58; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_59 = MAT_io_pipe_phv_out_data_59; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_60 = MAT_io_pipe_phv_out_data_60; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_61 = MAT_io_pipe_phv_out_data_61; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_62 = MAT_io_pipe_phv_out_data_62; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_63 = MAT_io_pipe_phv_out_data_63; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_64 = MAT_io_pipe_phv_out_data_64; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_65 = MAT_io_pipe_phv_out_data_65; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_66 = MAT_io_pipe_phv_out_data_66; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_67 = MAT_io_pipe_phv_out_data_67; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_68 = MAT_io_pipe_phv_out_data_68; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_69 = MAT_io_pipe_phv_out_data_69; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_70 = MAT_io_pipe_phv_out_data_70; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_71 = MAT_io_pipe_phv_out_data_71; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_72 = MAT_io_pipe_phv_out_data_72; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_73 = MAT_io_pipe_phv_out_data_73; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_74 = MAT_io_pipe_phv_out_data_74; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_75 = MAT_io_pipe_phv_out_data_75; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_76 = MAT_io_pipe_phv_out_data_76; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_77 = MAT_io_pipe_phv_out_data_77; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_78 = MAT_io_pipe_phv_out_data_78; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_79 = MAT_io_pipe_phv_out_data_79; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_80 = MAT_io_pipe_phv_out_data_80; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_81 = MAT_io_pipe_phv_out_data_81; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_82 = MAT_io_pipe_phv_out_data_82; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_83 = MAT_io_pipe_phv_out_data_83; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_84 = MAT_io_pipe_phv_out_data_84; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_85 = MAT_io_pipe_phv_out_data_85; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_86 = MAT_io_pipe_phv_out_data_86; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_87 = MAT_io_pipe_phv_out_data_87; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_88 = MAT_io_pipe_phv_out_data_88; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_89 = MAT_io_pipe_phv_out_data_89; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_90 = MAT_io_pipe_phv_out_data_90; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_91 = MAT_io_pipe_phv_out_data_91; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_92 = MAT_io_pipe_phv_out_data_92; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_93 = MAT_io_pipe_phv_out_data_93; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_94 = MAT_io_pipe_phv_out_data_94; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_95 = MAT_io_pipe_phv_out_data_95; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_96 = MAT_io_pipe_phv_out_data_96; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_97 = MAT_io_pipe_phv_out_data_97; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_98 = MAT_io_pipe_phv_out_data_98; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_99 = MAT_io_pipe_phv_out_data_99; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_100 = MAT_io_pipe_phv_out_data_100; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_101 = MAT_io_pipe_phv_out_data_101; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_102 = MAT_io_pipe_phv_out_data_102; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_103 = MAT_io_pipe_phv_out_data_103; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_104 = MAT_io_pipe_phv_out_data_104; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_105 = MAT_io_pipe_phv_out_data_105; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_106 = MAT_io_pipe_phv_out_data_106; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_107 = MAT_io_pipe_phv_out_data_107; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_108 = MAT_io_pipe_phv_out_data_108; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_109 = MAT_io_pipe_phv_out_data_109; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_110 = MAT_io_pipe_phv_out_data_110; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_111 = MAT_io_pipe_phv_out_data_111; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_112 = MAT_io_pipe_phv_out_data_112; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_113 = MAT_io_pipe_phv_out_data_113; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_114 = MAT_io_pipe_phv_out_data_114; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_115 = MAT_io_pipe_phv_out_data_115; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_116 = MAT_io_pipe_phv_out_data_116; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_117 = MAT_io_pipe_phv_out_data_117; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_118 = MAT_io_pipe_phv_out_data_118; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_119 = MAT_io_pipe_phv_out_data_119; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_120 = MAT_io_pipe_phv_out_data_120; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_121 = MAT_io_pipe_phv_out_data_121; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_122 = MAT_io_pipe_phv_out_data_122; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_123 = MAT_io_pipe_phv_out_data_123; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_124 = MAT_io_pipe_phv_out_data_124; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_125 = MAT_io_pipe_phv_out_data_125; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_126 = MAT_io_pipe_phv_out_data_126; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_127 = MAT_io_pipe_phv_out_data_127; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_128 = MAT_io_pipe_phv_out_data_128; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_129 = MAT_io_pipe_phv_out_data_129; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_130 = MAT_io_pipe_phv_out_data_130; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_131 = MAT_io_pipe_phv_out_data_131; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_132 = MAT_io_pipe_phv_out_data_132; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_133 = MAT_io_pipe_phv_out_data_133; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_134 = MAT_io_pipe_phv_out_data_134; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_135 = MAT_io_pipe_phv_out_data_135; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_136 = MAT_io_pipe_phv_out_data_136; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_137 = MAT_io_pipe_phv_out_data_137; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_138 = MAT_io_pipe_phv_out_data_138; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_139 = MAT_io_pipe_phv_out_data_139; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_140 = MAT_io_pipe_phv_out_data_140; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_141 = MAT_io_pipe_phv_out_data_141; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_142 = MAT_io_pipe_phv_out_data_142; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_143 = MAT_io_pipe_phv_out_data_143; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_144 = MAT_io_pipe_phv_out_data_144; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_145 = MAT_io_pipe_phv_out_data_145; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_146 = MAT_io_pipe_phv_out_data_146; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_147 = MAT_io_pipe_phv_out_data_147; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_148 = MAT_io_pipe_phv_out_data_148; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_149 = MAT_io_pipe_phv_out_data_149; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_150 = MAT_io_pipe_phv_out_data_150; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_151 = MAT_io_pipe_phv_out_data_151; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_152 = MAT_io_pipe_phv_out_data_152; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_153 = MAT_io_pipe_phv_out_data_153; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_154 = MAT_io_pipe_phv_out_data_154; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_155 = MAT_io_pipe_phv_out_data_155; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_156 = MAT_io_pipe_phv_out_data_156; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_157 = MAT_io_pipe_phv_out_data_157; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_158 = MAT_io_pipe_phv_out_data_158; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_159 = MAT_io_pipe_phv_out_data_159; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_160 = MAT_io_pipe_phv_out_data_160; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_161 = MAT_io_pipe_phv_out_data_161; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_162 = MAT_io_pipe_phv_out_data_162; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_163 = MAT_io_pipe_phv_out_data_163; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_164 = MAT_io_pipe_phv_out_data_164; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_165 = MAT_io_pipe_phv_out_data_165; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_166 = MAT_io_pipe_phv_out_data_166; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_167 = MAT_io_pipe_phv_out_data_167; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_168 = MAT_io_pipe_phv_out_data_168; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_169 = MAT_io_pipe_phv_out_data_169; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_170 = MAT_io_pipe_phv_out_data_170; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_171 = MAT_io_pipe_phv_out_data_171; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_172 = MAT_io_pipe_phv_out_data_172; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_173 = MAT_io_pipe_phv_out_data_173; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_174 = MAT_io_pipe_phv_out_data_174; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_175 = MAT_io_pipe_phv_out_data_175; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_176 = MAT_io_pipe_phv_out_data_176; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_177 = MAT_io_pipe_phv_out_data_177; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_178 = MAT_io_pipe_phv_out_data_178; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_179 = MAT_io_pipe_phv_out_data_179; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_180 = MAT_io_pipe_phv_out_data_180; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_181 = MAT_io_pipe_phv_out_data_181; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_182 = MAT_io_pipe_phv_out_data_182; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_183 = MAT_io_pipe_phv_out_data_183; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_184 = MAT_io_pipe_phv_out_data_184; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_185 = MAT_io_pipe_phv_out_data_185; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_186 = MAT_io_pipe_phv_out_data_186; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_187 = MAT_io_pipe_phv_out_data_187; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_188 = MAT_io_pipe_phv_out_data_188; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_189 = MAT_io_pipe_phv_out_data_189; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_190 = MAT_io_pipe_phv_out_data_190; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_191 = MAT_io_pipe_phv_out_data_191; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_192 = MAT_io_pipe_phv_out_data_192; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_193 = MAT_io_pipe_phv_out_data_193; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_194 = MAT_io_pipe_phv_out_data_194; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_195 = MAT_io_pipe_phv_out_data_195; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_196 = MAT_io_pipe_phv_out_data_196; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_197 = MAT_io_pipe_phv_out_data_197; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_198 = MAT_io_pipe_phv_out_data_198; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_199 = MAT_io_pipe_phv_out_data_199; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_200 = MAT_io_pipe_phv_out_data_200; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_201 = MAT_io_pipe_phv_out_data_201; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_202 = MAT_io_pipe_phv_out_data_202; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_203 = MAT_io_pipe_phv_out_data_203; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_204 = MAT_io_pipe_phv_out_data_204; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_205 = MAT_io_pipe_phv_out_data_205; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_206 = MAT_io_pipe_phv_out_data_206; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_207 = MAT_io_pipe_phv_out_data_207; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_208 = MAT_io_pipe_phv_out_data_208; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_209 = MAT_io_pipe_phv_out_data_209; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_210 = MAT_io_pipe_phv_out_data_210; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_211 = MAT_io_pipe_phv_out_data_211; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_212 = MAT_io_pipe_phv_out_data_212; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_213 = MAT_io_pipe_phv_out_data_213; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_214 = MAT_io_pipe_phv_out_data_214; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_215 = MAT_io_pipe_phv_out_data_215; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_216 = MAT_io_pipe_phv_out_data_216; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_217 = MAT_io_pipe_phv_out_data_217; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_218 = MAT_io_pipe_phv_out_data_218; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_219 = MAT_io_pipe_phv_out_data_219; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_220 = MAT_io_pipe_phv_out_data_220; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_221 = MAT_io_pipe_phv_out_data_221; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_222 = MAT_io_pipe_phv_out_data_222; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_223 = MAT_io_pipe_phv_out_data_223; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_224 = MAT_io_pipe_phv_out_data_224; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_225 = MAT_io_pipe_phv_out_data_225; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_226 = MAT_io_pipe_phv_out_data_226; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_227 = MAT_io_pipe_phv_out_data_227; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_228 = MAT_io_pipe_phv_out_data_228; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_229 = MAT_io_pipe_phv_out_data_229; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_230 = MAT_io_pipe_phv_out_data_230; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_231 = MAT_io_pipe_phv_out_data_231; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_232 = MAT_io_pipe_phv_out_data_232; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_233 = MAT_io_pipe_phv_out_data_233; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_234 = MAT_io_pipe_phv_out_data_234; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_235 = MAT_io_pipe_phv_out_data_235; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_236 = MAT_io_pipe_phv_out_data_236; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_237 = MAT_io_pipe_phv_out_data_237; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_238 = MAT_io_pipe_phv_out_data_238; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_239 = MAT_io_pipe_phv_out_data_239; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_240 = MAT_io_pipe_phv_out_data_240; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_241 = MAT_io_pipe_phv_out_data_241; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_242 = MAT_io_pipe_phv_out_data_242; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_243 = MAT_io_pipe_phv_out_data_243; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_244 = MAT_io_pipe_phv_out_data_244; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_245 = MAT_io_pipe_phv_out_data_245; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_246 = MAT_io_pipe_phv_out_data_246; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_247 = MAT_io_pipe_phv_out_data_247; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_248 = MAT_io_pipe_phv_out_data_248; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_249 = MAT_io_pipe_phv_out_data_249; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_250 = MAT_io_pipe_phv_out_data_250; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_251 = MAT_io_pipe_phv_out_data_251; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_252 = MAT_io_pipe_phv_out_data_252; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_253 = MAT_io_pipe_phv_out_data_253; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_254 = MAT_io_pipe_phv_out_data_254; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_255 = MAT_io_pipe_phv_out_data_255; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_0 = MAT_io_pipe_phv_out_header_0; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_1 = MAT_io_pipe_phv_out_header_1; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_2 = MAT_io_pipe_phv_out_header_2; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_3 = MAT_io_pipe_phv_out_header_3; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_4 = MAT_io_pipe_phv_out_header_4; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_5 = MAT_io_pipe_phv_out_header_5; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_6 = MAT_io_pipe_phv_out_header_6; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_7 = MAT_io_pipe_phv_out_header_7; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_8 = MAT_io_pipe_phv_out_header_8; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_9 = MAT_io_pipe_phv_out_header_9; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_10 = MAT_io_pipe_phv_out_header_10; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_11 = MAT_io_pipe_phv_out_header_11; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_12 = MAT_io_pipe_phv_out_header_12; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_13 = MAT_io_pipe_phv_out_header_13; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_14 = MAT_io_pipe_phv_out_header_14; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_15 = MAT_io_pipe_phv_out_header_15; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_parse_current_state = MAT_io_pipe_phv_out_parse_current_state; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_parse_current_offset = MAT_io_pipe_phv_out_parse_current_offset; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_parse_transition_field = MAT_io_pipe_phv_out_parse_transition_field; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_next_processor_id = MAT_io_pipe_phv_out_next_processor_id; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_next_config_id = MAT_io_pipe_phv_out_next_config_id; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_is_valid_processor = MAT_io_pipe_phv_out_is_valid_processor; // @[processor.scala 24:24]
  assign EXE_io_hit = MAT_io_hit; // @[processor.scala 25:24]
  assign EXE_io_match_value = MAT_io_match_value; // @[processor.scala 26:24]
  assign EXE_io_action_mod_en_0 = io_mod_act_mod_en_0; // @[processor.scala 27:24]
  assign EXE_io_action_mod_en_1 = io_mod_act_mod_en_1; // @[processor.scala 27:24]
  assign EXE_io_action_mod_addr = io_mod_act_mod_addr; // @[processor.scala 27:24]
  assign EXE_io_action_mod_data_0 = io_mod_act_mod_data_0; // @[processor.scala 27:24]
  assign EXE_io_action_mod_data_1 = io_mod_act_mod_data_1; // @[processor.scala 27:24]
endmodule
