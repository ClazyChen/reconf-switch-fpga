module MatchGetKey(
  input          clock,
  input  [7:0]   io_pipe_phv_in_data_0,
  input  [7:0]   io_pipe_phv_in_data_1,
  input  [7:0]   io_pipe_phv_in_data_2,
  input  [7:0]   io_pipe_phv_in_data_3,
  input  [7:0]   io_pipe_phv_in_data_4,
  input  [7:0]   io_pipe_phv_in_data_5,
  input  [7:0]   io_pipe_phv_in_data_6,
  input  [7:0]   io_pipe_phv_in_data_7,
  input  [7:0]   io_pipe_phv_in_data_8,
  input  [7:0]   io_pipe_phv_in_data_9,
  input  [7:0]   io_pipe_phv_in_data_10,
  input  [7:0]   io_pipe_phv_in_data_11,
  input  [7:0]   io_pipe_phv_in_data_12,
  input  [7:0]   io_pipe_phv_in_data_13,
  input  [7:0]   io_pipe_phv_in_data_14,
  input  [7:0]   io_pipe_phv_in_data_15,
  input  [7:0]   io_pipe_phv_in_data_16,
  input  [7:0]   io_pipe_phv_in_data_17,
  input  [7:0]   io_pipe_phv_in_data_18,
  input  [7:0]   io_pipe_phv_in_data_19,
  input  [7:0]   io_pipe_phv_in_data_20,
  input  [7:0]   io_pipe_phv_in_data_21,
  input  [7:0]   io_pipe_phv_in_data_22,
  input  [7:0]   io_pipe_phv_in_data_23,
  input  [7:0]   io_pipe_phv_in_data_24,
  input  [7:0]   io_pipe_phv_in_data_25,
  input  [7:0]   io_pipe_phv_in_data_26,
  input  [7:0]   io_pipe_phv_in_data_27,
  input  [7:0]   io_pipe_phv_in_data_28,
  input  [7:0]   io_pipe_phv_in_data_29,
  input  [7:0]   io_pipe_phv_in_data_30,
  input  [7:0]   io_pipe_phv_in_data_31,
  input  [7:0]   io_pipe_phv_in_data_32,
  input  [7:0]   io_pipe_phv_in_data_33,
  input  [7:0]   io_pipe_phv_in_data_34,
  input  [7:0]   io_pipe_phv_in_data_35,
  input  [7:0]   io_pipe_phv_in_data_36,
  input  [7:0]   io_pipe_phv_in_data_37,
  input  [7:0]   io_pipe_phv_in_data_38,
  input  [7:0]   io_pipe_phv_in_data_39,
  input  [7:0]   io_pipe_phv_in_data_40,
  input  [7:0]   io_pipe_phv_in_data_41,
  input  [7:0]   io_pipe_phv_in_data_42,
  input  [7:0]   io_pipe_phv_in_data_43,
  input  [7:0]   io_pipe_phv_in_data_44,
  input  [7:0]   io_pipe_phv_in_data_45,
  input  [7:0]   io_pipe_phv_in_data_46,
  input  [7:0]   io_pipe_phv_in_data_47,
  input  [7:0]   io_pipe_phv_in_data_48,
  input  [7:0]   io_pipe_phv_in_data_49,
  input  [7:0]   io_pipe_phv_in_data_50,
  input  [7:0]   io_pipe_phv_in_data_51,
  input  [7:0]   io_pipe_phv_in_data_52,
  input  [7:0]   io_pipe_phv_in_data_53,
  input  [7:0]   io_pipe_phv_in_data_54,
  input  [7:0]   io_pipe_phv_in_data_55,
  input  [7:0]   io_pipe_phv_in_data_56,
  input  [7:0]   io_pipe_phv_in_data_57,
  input  [7:0]   io_pipe_phv_in_data_58,
  input  [7:0]   io_pipe_phv_in_data_59,
  input  [7:0]   io_pipe_phv_in_data_60,
  input  [7:0]   io_pipe_phv_in_data_61,
  input  [7:0]   io_pipe_phv_in_data_62,
  input  [7:0]   io_pipe_phv_in_data_63,
  input  [7:0]   io_pipe_phv_in_data_64,
  input  [7:0]   io_pipe_phv_in_data_65,
  input  [7:0]   io_pipe_phv_in_data_66,
  input  [7:0]   io_pipe_phv_in_data_67,
  input  [7:0]   io_pipe_phv_in_data_68,
  input  [7:0]   io_pipe_phv_in_data_69,
  input  [7:0]   io_pipe_phv_in_data_70,
  input  [7:0]   io_pipe_phv_in_data_71,
  input  [7:0]   io_pipe_phv_in_data_72,
  input  [7:0]   io_pipe_phv_in_data_73,
  input  [7:0]   io_pipe_phv_in_data_74,
  input  [7:0]   io_pipe_phv_in_data_75,
  input  [7:0]   io_pipe_phv_in_data_76,
  input  [7:0]   io_pipe_phv_in_data_77,
  input  [7:0]   io_pipe_phv_in_data_78,
  input  [7:0]   io_pipe_phv_in_data_79,
  input  [7:0]   io_pipe_phv_in_data_80,
  input  [7:0]   io_pipe_phv_in_data_81,
  input  [7:0]   io_pipe_phv_in_data_82,
  input  [7:0]   io_pipe_phv_in_data_83,
  input  [7:0]   io_pipe_phv_in_data_84,
  input  [7:0]   io_pipe_phv_in_data_85,
  input  [7:0]   io_pipe_phv_in_data_86,
  input  [7:0]   io_pipe_phv_in_data_87,
  input  [7:0]   io_pipe_phv_in_data_88,
  input  [7:0]   io_pipe_phv_in_data_89,
  input  [7:0]   io_pipe_phv_in_data_90,
  input  [7:0]   io_pipe_phv_in_data_91,
  input  [7:0]   io_pipe_phv_in_data_92,
  input  [7:0]   io_pipe_phv_in_data_93,
  input  [7:0]   io_pipe_phv_in_data_94,
  input  [7:0]   io_pipe_phv_in_data_95,
  input  [7:0]   io_pipe_phv_in_data_96,
  input  [7:0]   io_pipe_phv_in_data_97,
  input  [7:0]   io_pipe_phv_in_data_98,
  input  [7:0]   io_pipe_phv_in_data_99,
  input  [7:0]   io_pipe_phv_in_data_100,
  input  [7:0]   io_pipe_phv_in_data_101,
  input  [7:0]   io_pipe_phv_in_data_102,
  input  [7:0]   io_pipe_phv_in_data_103,
  input  [7:0]   io_pipe_phv_in_data_104,
  input  [7:0]   io_pipe_phv_in_data_105,
  input  [7:0]   io_pipe_phv_in_data_106,
  input  [7:0]   io_pipe_phv_in_data_107,
  input  [7:0]   io_pipe_phv_in_data_108,
  input  [7:0]   io_pipe_phv_in_data_109,
  input  [7:0]   io_pipe_phv_in_data_110,
  input  [7:0]   io_pipe_phv_in_data_111,
  input  [7:0]   io_pipe_phv_in_data_112,
  input  [7:0]   io_pipe_phv_in_data_113,
  input  [7:0]   io_pipe_phv_in_data_114,
  input  [7:0]   io_pipe_phv_in_data_115,
  input  [7:0]   io_pipe_phv_in_data_116,
  input  [7:0]   io_pipe_phv_in_data_117,
  input  [7:0]   io_pipe_phv_in_data_118,
  input  [7:0]   io_pipe_phv_in_data_119,
  input  [7:0]   io_pipe_phv_in_data_120,
  input  [7:0]   io_pipe_phv_in_data_121,
  input  [7:0]   io_pipe_phv_in_data_122,
  input  [7:0]   io_pipe_phv_in_data_123,
  input  [7:0]   io_pipe_phv_in_data_124,
  input  [7:0]   io_pipe_phv_in_data_125,
  input  [7:0]   io_pipe_phv_in_data_126,
  input  [7:0]   io_pipe_phv_in_data_127,
  input  [7:0]   io_pipe_phv_in_data_128,
  input  [7:0]   io_pipe_phv_in_data_129,
  input  [7:0]   io_pipe_phv_in_data_130,
  input  [7:0]   io_pipe_phv_in_data_131,
  input  [7:0]   io_pipe_phv_in_data_132,
  input  [7:0]   io_pipe_phv_in_data_133,
  input  [7:0]   io_pipe_phv_in_data_134,
  input  [7:0]   io_pipe_phv_in_data_135,
  input  [7:0]   io_pipe_phv_in_data_136,
  input  [7:0]   io_pipe_phv_in_data_137,
  input  [7:0]   io_pipe_phv_in_data_138,
  input  [7:0]   io_pipe_phv_in_data_139,
  input  [7:0]   io_pipe_phv_in_data_140,
  input  [7:0]   io_pipe_phv_in_data_141,
  input  [7:0]   io_pipe_phv_in_data_142,
  input  [7:0]   io_pipe_phv_in_data_143,
  input  [7:0]   io_pipe_phv_in_data_144,
  input  [7:0]   io_pipe_phv_in_data_145,
  input  [7:0]   io_pipe_phv_in_data_146,
  input  [7:0]   io_pipe_phv_in_data_147,
  input  [7:0]   io_pipe_phv_in_data_148,
  input  [7:0]   io_pipe_phv_in_data_149,
  input  [7:0]   io_pipe_phv_in_data_150,
  input  [7:0]   io_pipe_phv_in_data_151,
  input  [7:0]   io_pipe_phv_in_data_152,
  input  [7:0]   io_pipe_phv_in_data_153,
  input  [7:0]   io_pipe_phv_in_data_154,
  input  [7:0]   io_pipe_phv_in_data_155,
  input  [7:0]   io_pipe_phv_in_data_156,
  input  [7:0]   io_pipe_phv_in_data_157,
  input  [7:0]   io_pipe_phv_in_data_158,
  input  [7:0]   io_pipe_phv_in_data_159,
  input  [15:0]  io_pipe_phv_in_header_0,
  input  [15:0]  io_pipe_phv_in_header_1,
  input  [15:0]  io_pipe_phv_in_header_2,
  input  [15:0]  io_pipe_phv_in_header_3,
  input  [15:0]  io_pipe_phv_in_header_4,
  input  [15:0]  io_pipe_phv_in_header_5,
  input  [15:0]  io_pipe_phv_in_header_6,
  input  [15:0]  io_pipe_phv_in_header_7,
  input  [15:0]  io_pipe_phv_in_header_8,
  input  [15:0]  io_pipe_phv_in_header_9,
  input  [15:0]  io_pipe_phv_in_header_10,
  input  [15:0]  io_pipe_phv_in_header_11,
  input  [15:0]  io_pipe_phv_in_header_12,
  input  [15:0]  io_pipe_phv_in_header_13,
  input  [15:0]  io_pipe_phv_in_header_14,
  input  [15:0]  io_pipe_phv_in_header_15,
  input  [7:0]   io_pipe_phv_in_parse_current_state,
  input  [7:0]   io_pipe_phv_in_parse_current_offset,
  input  [15:0]  io_pipe_phv_in_parse_transition_field,
  input  [3:0]   io_pipe_phv_in_next_processor_id,
  input          io_pipe_phv_in_next_config_id,
  input          io_pipe_phv_in_is_valid_processor,
  output [7:0]   io_pipe_phv_out_data_0,
  output [7:0]   io_pipe_phv_out_data_1,
  output [7:0]   io_pipe_phv_out_data_2,
  output [7:0]   io_pipe_phv_out_data_3,
  output [7:0]   io_pipe_phv_out_data_4,
  output [7:0]   io_pipe_phv_out_data_5,
  output [7:0]   io_pipe_phv_out_data_6,
  output [7:0]   io_pipe_phv_out_data_7,
  output [7:0]   io_pipe_phv_out_data_8,
  output [7:0]   io_pipe_phv_out_data_9,
  output [7:0]   io_pipe_phv_out_data_10,
  output [7:0]   io_pipe_phv_out_data_11,
  output [7:0]   io_pipe_phv_out_data_12,
  output [7:0]   io_pipe_phv_out_data_13,
  output [7:0]   io_pipe_phv_out_data_14,
  output [7:0]   io_pipe_phv_out_data_15,
  output [7:0]   io_pipe_phv_out_data_16,
  output [7:0]   io_pipe_phv_out_data_17,
  output [7:0]   io_pipe_phv_out_data_18,
  output [7:0]   io_pipe_phv_out_data_19,
  output [7:0]   io_pipe_phv_out_data_20,
  output [7:0]   io_pipe_phv_out_data_21,
  output [7:0]   io_pipe_phv_out_data_22,
  output [7:0]   io_pipe_phv_out_data_23,
  output [7:0]   io_pipe_phv_out_data_24,
  output [7:0]   io_pipe_phv_out_data_25,
  output [7:0]   io_pipe_phv_out_data_26,
  output [7:0]   io_pipe_phv_out_data_27,
  output [7:0]   io_pipe_phv_out_data_28,
  output [7:0]   io_pipe_phv_out_data_29,
  output [7:0]   io_pipe_phv_out_data_30,
  output [7:0]   io_pipe_phv_out_data_31,
  output [7:0]   io_pipe_phv_out_data_32,
  output [7:0]   io_pipe_phv_out_data_33,
  output [7:0]   io_pipe_phv_out_data_34,
  output [7:0]   io_pipe_phv_out_data_35,
  output [7:0]   io_pipe_phv_out_data_36,
  output [7:0]   io_pipe_phv_out_data_37,
  output [7:0]   io_pipe_phv_out_data_38,
  output [7:0]   io_pipe_phv_out_data_39,
  output [7:0]   io_pipe_phv_out_data_40,
  output [7:0]   io_pipe_phv_out_data_41,
  output [7:0]   io_pipe_phv_out_data_42,
  output [7:0]   io_pipe_phv_out_data_43,
  output [7:0]   io_pipe_phv_out_data_44,
  output [7:0]   io_pipe_phv_out_data_45,
  output [7:0]   io_pipe_phv_out_data_46,
  output [7:0]   io_pipe_phv_out_data_47,
  output [7:0]   io_pipe_phv_out_data_48,
  output [7:0]   io_pipe_phv_out_data_49,
  output [7:0]   io_pipe_phv_out_data_50,
  output [7:0]   io_pipe_phv_out_data_51,
  output [7:0]   io_pipe_phv_out_data_52,
  output [7:0]   io_pipe_phv_out_data_53,
  output [7:0]   io_pipe_phv_out_data_54,
  output [7:0]   io_pipe_phv_out_data_55,
  output [7:0]   io_pipe_phv_out_data_56,
  output [7:0]   io_pipe_phv_out_data_57,
  output [7:0]   io_pipe_phv_out_data_58,
  output [7:0]   io_pipe_phv_out_data_59,
  output [7:0]   io_pipe_phv_out_data_60,
  output [7:0]   io_pipe_phv_out_data_61,
  output [7:0]   io_pipe_phv_out_data_62,
  output [7:0]   io_pipe_phv_out_data_63,
  output [7:0]   io_pipe_phv_out_data_64,
  output [7:0]   io_pipe_phv_out_data_65,
  output [7:0]   io_pipe_phv_out_data_66,
  output [7:0]   io_pipe_phv_out_data_67,
  output [7:0]   io_pipe_phv_out_data_68,
  output [7:0]   io_pipe_phv_out_data_69,
  output [7:0]   io_pipe_phv_out_data_70,
  output [7:0]   io_pipe_phv_out_data_71,
  output [7:0]   io_pipe_phv_out_data_72,
  output [7:0]   io_pipe_phv_out_data_73,
  output [7:0]   io_pipe_phv_out_data_74,
  output [7:0]   io_pipe_phv_out_data_75,
  output [7:0]   io_pipe_phv_out_data_76,
  output [7:0]   io_pipe_phv_out_data_77,
  output [7:0]   io_pipe_phv_out_data_78,
  output [7:0]   io_pipe_phv_out_data_79,
  output [7:0]   io_pipe_phv_out_data_80,
  output [7:0]   io_pipe_phv_out_data_81,
  output [7:0]   io_pipe_phv_out_data_82,
  output [7:0]   io_pipe_phv_out_data_83,
  output [7:0]   io_pipe_phv_out_data_84,
  output [7:0]   io_pipe_phv_out_data_85,
  output [7:0]   io_pipe_phv_out_data_86,
  output [7:0]   io_pipe_phv_out_data_87,
  output [7:0]   io_pipe_phv_out_data_88,
  output [7:0]   io_pipe_phv_out_data_89,
  output [7:0]   io_pipe_phv_out_data_90,
  output [7:0]   io_pipe_phv_out_data_91,
  output [7:0]   io_pipe_phv_out_data_92,
  output [7:0]   io_pipe_phv_out_data_93,
  output [7:0]   io_pipe_phv_out_data_94,
  output [7:0]   io_pipe_phv_out_data_95,
  output [7:0]   io_pipe_phv_out_data_96,
  output [7:0]   io_pipe_phv_out_data_97,
  output [7:0]   io_pipe_phv_out_data_98,
  output [7:0]   io_pipe_phv_out_data_99,
  output [7:0]   io_pipe_phv_out_data_100,
  output [7:0]   io_pipe_phv_out_data_101,
  output [7:0]   io_pipe_phv_out_data_102,
  output [7:0]   io_pipe_phv_out_data_103,
  output [7:0]   io_pipe_phv_out_data_104,
  output [7:0]   io_pipe_phv_out_data_105,
  output [7:0]   io_pipe_phv_out_data_106,
  output [7:0]   io_pipe_phv_out_data_107,
  output [7:0]   io_pipe_phv_out_data_108,
  output [7:0]   io_pipe_phv_out_data_109,
  output [7:0]   io_pipe_phv_out_data_110,
  output [7:0]   io_pipe_phv_out_data_111,
  output [7:0]   io_pipe_phv_out_data_112,
  output [7:0]   io_pipe_phv_out_data_113,
  output [7:0]   io_pipe_phv_out_data_114,
  output [7:0]   io_pipe_phv_out_data_115,
  output [7:0]   io_pipe_phv_out_data_116,
  output [7:0]   io_pipe_phv_out_data_117,
  output [7:0]   io_pipe_phv_out_data_118,
  output [7:0]   io_pipe_phv_out_data_119,
  output [7:0]   io_pipe_phv_out_data_120,
  output [7:0]   io_pipe_phv_out_data_121,
  output [7:0]   io_pipe_phv_out_data_122,
  output [7:0]   io_pipe_phv_out_data_123,
  output [7:0]   io_pipe_phv_out_data_124,
  output [7:0]   io_pipe_phv_out_data_125,
  output [7:0]   io_pipe_phv_out_data_126,
  output [7:0]   io_pipe_phv_out_data_127,
  output [7:0]   io_pipe_phv_out_data_128,
  output [7:0]   io_pipe_phv_out_data_129,
  output [7:0]   io_pipe_phv_out_data_130,
  output [7:0]   io_pipe_phv_out_data_131,
  output [7:0]   io_pipe_phv_out_data_132,
  output [7:0]   io_pipe_phv_out_data_133,
  output [7:0]   io_pipe_phv_out_data_134,
  output [7:0]   io_pipe_phv_out_data_135,
  output [7:0]   io_pipe_phv_out_data_136,
  output [7:0]   io_pipe_phv_out_data_137,
  output [7:0]   io_pipe_phv_out_data_138,
  output [7:0]   io_pipe_phv_out_data_139,
  output [7:0]   io_pipe_phv_out_data_140,
  output [7:0]   io_pipe_phv_out_data_141,
  output [7:0]   io_pipe_phv_out_data_142,
  output [7:0]   io_pipe_phv_out_data_143,
  output [7:0]   io_pipe_phv_out_data_144,
  output [7:0]   io_pipe_phv_out_data_145,
  output [7:0]   io_pipe_phv_out_data_146,
  output [7:0]   io_pipe_phv_out_data_147,
  output [7:0]   io_pipe_phv_out_data_148,
  output [7:0]   io_pipe_phv_out_data_149,
  output [7:0]   io_pipe_phv_out_data_150,
  output [7:0]   io_pipe_phv_out_data_151,
  output [7:0]   io_pipe_phv_out_data_152,
  output [7:0]   io_pipe_phv_out_data_153,
  output [7:0]   io_pipe_phv_out_data_154,
  output [7:0]   io_pipe_phv_out_data_155,
  output [7:0]   io_pipe_phv_out_data_156,
  output [7:0]   io_pipe_phv_out_data_157,
  output [7:0]   io_pipe_phv_out_data_158,
  output [7:0]   io_pipe_phv_out_data_159,
  output [15:0]  io_pipe_phv_out_header_0,
  output [15:0]  io_pipe_phv_out_header_1,
  output [15:0]  io_pipe_phv_out_header_2,
  output [15:0]  io_pipe_phv_out_header_3,
  output [15:0]  io_pipe_phv_out_header_4,
  output [15:0]  io_pipe_phv_out_header_5,
  output [15:0]  io_pipe_phv_out_header_6,
  output [15:0]  io_pipe_phv_out_header_7,
  output [15:0]  io_pipe_phv_out_header_8,
  output [15:0]  io_pipe_phv_out_header_9,
  output [15:0]  io_pipe_phv_out_header_10,
  output [15:0]  io_pipe_phv_out_header_11,
  output [15:0]  io_pipe_phv_out_header_12,
  output [15:0]  io_pipe_phv_out_header_13,
  output [15:0]  io_pipe_phv_out_header_14,
  output [15:0]  io_pipe_phv_out_header_15,
  output [7:0]   io_pipe_phv_out_parse_current_state,
  output [7:0]   io_pipe_phv_out_parse_current_offset,
  output [15:0]  io_pipe_phv_out_parse_transition_field,
  output [3:0]   io_pipe_phv_out_next_processor_id,
  output         io_pipe_phv_out_next_config_id,
  output         io_pipe_phv_out_is_valid_processor,
  input  [7:0]   io_key_config_0_key_length,
  input  [7:0]   io_key_config_1_key_length,
  input  [7:0]   io_key_offset,
  output [191:0] io_match_key
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[matcher.scala 58:22]
  reg [7:0] phv_data_1; // @[matcher.scala 58:22]
  reg [7:0] phv_data_2; // @[matcher.scala 58:22]
  reg [7:0] phv_data_3; // @[matcher.scala 58:22]
  reg [7:0] phv_data_4; // @[matcher.scala 58:22]
  reg [7:0] phv_data_5; // @[matcher.scala 58:22]
  reg [7:0] phv_data_6; // @[matcher.scala 58:22]
  reg [7:0] phv_data_7; // @[matcher.scala 58:22]
  reg [7:0] phv_data_8; // @[matcher.scala 58:22]
  reg [7:0] phv_data_9; // @[matcher.scala 58:22]
  reg [7:0] phv_data_10; // @[matcher.scala 58:22]
  reg [7:0] phv_data_11; // @[matcher.scala 58:22]
  reg [7:0] phv_data_12; // @[matcher.scala 58:22]
  reg [7:0] phv_data_13; // @[matcher.scala 58:22]
  reg [7:0] phv_data_14; // @[matcher.scala 58:22]
  reg [7:0] phv_data_15; // @[matcher.scala 58:22]
  reg [7:0] phv_data_16; // @[matcher.scala 58:22]
  reg [7:0] phv_data_17; // @[matcher.scala 58:22]
  reg [7:0] phv_data_18; // @[matcher.scala 58:22]
  reg [7:0] phv_data_19; // @[matcher.scala 58:22]
  reg [7:0] phv_data_20; // @[matcher.scala 58:22]
  reg [7:0] phv_data_21; // @[matcher.scala 58:22]
  reg [7:0] phv_data_22; // @[matcher.scala 58:22]
  reg [7:0] phv_data_23; // @[matcher.scala 58:22]
  reg [7:0] phv_data_24; // @[matcher.scala 58:22]
  reg [7:0] phv_data_25; // @[matcher.scala 58:22]
  reg [7:0] phv_data_26; // @[matcher.scala 58:22]
  reg [7:0] phv_data_27; // @[matcher.scala 58:22]
  reg [7:0] phv_data_28; // @[matcher.scala 58:22]
  reg [7:0] phv_data_29; // @[matcher.scala 58:22]
  reg [7:0] phv_data_30; // @[matcher.scala 58:22]
  reg [7:0] phv_data_31; // @[matcher.scala 58:22]
  reg [7:0] phv_data_32; // @[matcher.scala 58:22]
  reg [7:0] phv_data_33; // @[matcher.scala 58:22]
  reg [7:0] phv_data_34; // @[matcher.scala 58:22]
  reg [7:0] phv_data_35; // @[matcher.scala 58:22]
  reg [7:0] phv_data_36; // @[matcher.scala 58:22]
  reg [7:0] phv_data_37; // @[matcher.scala 58:22]
  reg [7:0] phv_data_38; // @[matcher.scala 58:22]
  reg [7:0] phv_data_39; // @[matcher.scala 58:22]
  reg [7:0] phv_data_40; // @[matcher.scala 58:22]
  reg [7:0] phv_data_41; // @[matcher.scala 58:22]
  reg [7:0] phv_data_42; // @[matcher.scala 58:22]
  reg [7:0] phv_data_43; // @[matcher.scala 58:22]
  reg [7:0] phv_data_44; // @[matcher.scala 58:22]
  reg [7:0] phv_data_45; // @[matcher.scala 58:22]
  reg [7:0] phv_data_46; // @[matcher.scala 58:22]
  reg [7:0] phv_data_47; // @[matcher.scala 58:22]
  reg [7:0] phv_data_48; // @[matcher.scala 58:22]
  reg [7:0] phv_data_49; // @[matcher.scala 58:22]
  reg [7:0] phv_data_50; // @[matcher.scala 58:22]
  reg [7:0] phv_data_51; // @[matcher.scala 58:22]
  reg [7:0] phv_data_52; // @[matcher.scala 58:22]
  reg [7:0] phv_data_53; // @[matcher.scala 58:22]
  reg [7:0] phv_data_54; // @[matcher.scala 58:22]
  reg [7:0] phv_data_55; // @[matcher.scala 58:22]
  reg [7:0] phv_data_56; // @[matcher.scala 58:22]
  reg [7:0] phv_data_57; // @[matcher.scala 58:22]
  reg [7:0] phv_data_58; // @[matcher.scala 58:22]
  reg [7:0] phv_data_59; // @[matcher.scala 58:22]
  reg [7:0] phv_data_60; // @[matcher.scala 58:22]
  reg [7:0] phv_data_61; // @[matcher.scala 58:22]
  reg [7:0] phv_data_62; // @[matcher.scala 58:22]
  reg [7:0] phv_data_63; // @[matcher.scala 58:22]
  reg [7:0] phv_data_64; // @[matcher.scala 58:22]
  reg [7:0] phv_data_65; // @[matcher.scala 58:22]
  reg [7:0] phv_data_66; // @[matcher.scala 58:22]
  reg [7:0] phv_data_67; // @[matcher.scala 58:22]
  reg [7:0] phv_data_68; // @[matcher.scala 58:22]
  reg [7:0] phv_data_69; // @[matcher.scala 58:22]
  reg [7:0] phv_data_70; // @[matcher.scala 58:22]
  reg [7:0] phv_data_71; // @[matcher.scala 58:22]
  reg [7:0] phv_data_72; // @[matcher.scala 58:22]
  reg [7:0] phv_data_73; // @[matcher.scala 58:22]
  reg [7:0] phv_data_74; // @[matcher.scala 58:22]
  reg [7:0] phv_data_75; // @[matcher.scala 58:22]
  reg [7:0] phv_data_76; // @[matcher.scala 58:22]
  reg [7:0] phv_data_77; // @[matcher.scala 58:22]
  reg [7:0] phv_data_78; // @[matcher.scala 58:22]
  reg [7:0] phv_data_79; // @[matcher.scala 58:22]
  reg [7:0] phv_data_80; // @[matcher.scala 58:22]
  reg [7:0] phv_data_81; // @[matcher.scala 58:22]
  reg [7:0] phv_data_82; // @[matcher.scala 58:22]
  reg [7:0] phv_data_83; // @[matcher.scala 58:22]
  reg [7:0] phv_data_84; // @[matcher.scala 58:22]
  reg [7:0] phv_data_85; // @[matcher.scala 58:22]
  reg [7:0] phv_data_86; // @[matcher.scala 58:22]
  reg [7:0] phv_data_87; // @[matcher.scala 58:22]
  reg [7:0] phv_data_88; // @[matcher.scala 58:22]
  reg [7:0] phv_data_89; // @[matcher.scala 58:22]
  reg [7:0] phv_data_90; // @[matcher.scala 58:22]
  reg [7:0] phv_data_91; // @[matcher.scala 58:22]
  reg [7:0] phv_data_92; // @[matcher.scala 58:22]
  reg [7:0] phv_data_93; // @[matcher.scala 58:22]
  reg [7:0] phv_data_94; // @[matcher.scala 58:22]
  reg [7:0] phv_data_95; // @[matcher.scala 58:22]
  reg [7:0] phv_data_96; // @[matcher.scala 58:22]
  reg [7:0] phv_data_97; // @[matcher.scala 58:22]
  reg [7:0] phv_data_98; // @[matcher.scala 58:22]
  reg [7:0] phv_data_99; // @[matcher.scala 58:22]
  reg [7:0] phv_data_100; // @[matcher.scala 58:22]
  reg [7:0] phv_data_101; // @[matcher.scala 58:22]
  reg [7:0] phv_data_102; // @[matcher.scala 58:22]
  reg [7:0] phv_data_103; // @[matcher.scala 58:22]
  reg [7:0] phv_data_104; // @[matcher.scala 58:22]
  reg [7:0] phv_data_105; // @[matcher.scala 58:22]
  reg [7:0] phv_data_106; // @[matcher.scala 58:22]
  reg [7:0] phv_data_107; // @[matcher.scala 58:22]
  reg [7:0] phv_data_108; // @[matcher.scala 58:22]
  reg [7:0] phv_data_109; // @[matcher.scala 58:22]
  reg [7:0] phv_data_110; // @[matcher.scala 58:22]
  reg [7:0] phv_data_111; // @[matcher.scala 58:22]
  reg [7:0] phv_data_112; // @[matcher.scala 58:22]
  reg [7:0] phv_data_113; // @[matcher.scala 58:22]
  reg [7:0] phv_data_114; // @[matcher.scala 58:22]
  reg [7:0] phv_data_115; // @[matcher.scala 58:22]
  reg [7:0] phv_data_116; // @[matcher.scala 58:22]
  reg [7:0] phv_data_117; // @[matcher.scala 58:22]
  reg [7:0] phv_data_118; // @[matcher.scala 58:22]
  reg [7:0] phv_data_119; // @[matcher.scala 58:22]
  reg [7:0] phv_data_120; // @[matcher.scala 58:22]
  reg [7:0] phv_data_121; // @[matcher.scala 58:22]
  reg [7:0] phv_data_122; // @[matcher.scala 58:22]
  reg [7:0] phv_data_123; // @[matcher.scala 58:22]
  reg [7:0] phv_data_124; // @[matcher.scala 58:22]
  reg [7:0] phv_data_125; // @[matcher.scala 58:22]
  reg [7:0] phv_data_126; // @[matcher.scala 58:22]
  reg [7:0] phv_data_127; // @[matcher.scala 58:22]
  reg [7:0] phv_data_128; // @[matcher.scala 58:22]
  reg [7:0] phv_data_129; // @[matcher.scala 58:22]
  reg [7:0] phv_data_130; // @[matcher.scala 58:22]
  reg [7:0] phv_data_131; // @[matcher.scala 58:22]
  reg [7:0] phv_data_132; // @[matcher.scala 58:22]
  reg [7:0] phv_data_133; // @[matcher.scala 58:22]
  reg [7:0] phv_data_134; // @[matcher.scala 58:22]
  reg [7:0] phv_data_135; // @[matcher.scala 58:22]
  reg [7:0] phv_data_136; // @[matcher.scala 58:22]
  reg [7:0] phv_data_137; // @[matcher.scala 58:22]
  reg [7:0] phv_data_138; // @[matcher.scala 58:22]
  reg [7:0] phv_data_139; // @[matcher.scala 58:22]
  reg [7:0] phv_data_140; // @[matcher.scala 58:22]
  reg [7:0] phv_data_141; // @[matcher.scala 58:22]
  reg [7:0] phv_data_142; // @[matcher.scala 58:22]
  reg [7:0] phv_data_143; // @[matcher.scala 58:22]
  reg [7:0] phv_data_144; // @[matcher.scala 58:22]
  reg [7:0] phv_data_145; // @[matcher.scala 58:22]
  reg [7:0] phv_data_146; // @[matcher.scala 58:22]
  reg [7:0] phv_data_147; // @[matcher.scala 58:22]
  reg [7:0] phv_data_148; // @[matcher.scala 58:22]
  reg [7:0] phv_data_149; // @[matcher.scala 58:22]
  reg [7:0] phv_data_150; // @[matcher.scala 58:22]
  reg [7:0] phv_data_151; // @[matcher.scala 58:22]
  reg [7:0] phv_data_152; // @[matcher.scala 58:22]
  reg [7:0] phv_data_153; // @[matcher.scala 58:22]
  reg [7:0] phv_data_154; // @[matcher.scala 58:22]
  reg [7:0] phv_data_155; // @[matcher.scala 58:22]
  reg [7:0] phv_data_156; // @[matcher.scala 58:22]
  reg [7:0] phv_data_157; // @[matcher.scala 58:22]
  reg [7:0] phv_data_158; // @[matcher.scala 58:22]
  reg [7:0] phv_data_159; // @[matcher.scala 58:22]
  reg [15:0] phv_header_0; // @[matcher.scala 58:22]
  reg [15:0] phv_header_1; // @[matcher.scala 58:22]
  reg [15:0] phv_header_2; // @[matcher.scala 58:22]
  reg [15:0] phv_header_3; // @[matcher.scala 58:22]
  reg [15:0] phv_header_4; // @[matcher.scala 58:22]
  reg [15:0] phv_header_5; // @[matcher.scala 58:22]
  reg [15:0] phv_header_6; // @[matcher.scala 58:22]
  reg [15:0] phv_header_7; // @[matcher.scala 58:22]
  reg [15:0] phv_header_8; // @[matcher.scala 58:22]
  reg [15:0] phv_header_9; // @[matcher.scala 58:22]
  reg [15:0] phv_header_10; // @[matcher.scala 58:22]
  reg [15:0] phv_header_11; // @[matcher.scala 58:22]
  reg [15:0] phv_header_12; // @[matcher.scala 58:22]
  reg [15:0] phv_header_13; // @[matcher.scala 58:22]
  reg [15:0] phv_header_14; // @[matcher.scala 58:22]
  reg [15:0] phv_header_15; // @[matcher.scala 58:22]
  reg [7:0] phv_parse_current_state; // @[matcher.scala 58:22]
  reg [7:0] phv_parse_current_offset; // @[matcher.scala 58:22]
  reg [15:0] phv_parse_transition_field; // @[matcher.scala 58:22]
  reg [3:0] phv_next_processor_id; // @[matcher.scala 58:22]
  reg  phv_next_config_id; // @[matcher.scala 58:22]
  reg  phv_is_valid_processor; // @[matcher.scala 58:22]
  reg [7:0] key_offset; // @[matcher.scala 62:29]
  wire [7:0] _GEN_6 = phv_next_config_id ? io_key_config_1_key_length : io_key_config_0_key_length; // @[matcher.scala 71:36 matcher.scala 71:36]
  wire [8:0] _match_key_bytes_23_T = {{1'd0}, key_offset}; // @[matcher.scala 72:98]
  wire [7:0] _GEN_9 = 8'h1 == _match_key_bytes_23_T[7:0] ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_10 = 8'h2 == _match_key_bytes_23_T[7:0] ? phv_data_2 : _GEN_9; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_11 = 8'h3 == _match_key_bytes_23_T[7:0] ? phv_data_3 : _GEN_10; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_12 = 8'h4 == _match_key_bytes_23_T[7:0] ? phv_data_4 : _GEN_11; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_13 = 8'h5 == _match_key_bytes_23_T[7:0] ? phv_data_5 : _GEN_12; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_14 = 8'h6 == _match_key_bytes_23_T[7:0] ? phv_data_6 : _GEN_13; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_15 = 8'h7 == _match_key_bytes_23_T[7:0] ? phv_data_7 : _GEN_14; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_16 = 8'h8 == _match_key_bytes_23_T[7:0] ? phv_data_8 : _GEN_15; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_17 = 8'h9 == _match_key_bytes_23_T[7:0] ? phv_data_9 : _GEN_16; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_18 = 8'ha == _match_key_bytes_23_T[7:0] ? phv_data_10 : _GEN_17; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_19 = 8'hb == _match_key_bytes_23_T[7:0] ? phv_data_11 : _GEN_18; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_20 = 8'hc == _match_key_bytes_23_T[7:0] ? phv_data_12 : _GEN_19; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_21 = 8'hd == _match_key_bytes_23_T[7:0] ? phv_data_13 : _GEN_20; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_22 = 8'he == _match_key_bytes_23_T[7:0] ? phv_data_14 : _GEN_21; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_23 = 8'hf == _match_key_bytes_23_T[7:0] ? phv_data_15 : _GEN_22; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_24 = 8'h10 == _match_key_bytes_23_T[7:0] ? phv_data_16 : _GEN_23; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_25 = 8'h11 == _match_key_bytes_23_T[7:0] ? phv_data_17 : _GEN_24; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_26 = 8'h12 == _match_key_bytes_23_T[7:0] ? phv_data_18 : _GEN_25; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_27 = 8'h13 == _match_key_bytes_23_T[7:0] ? phv_data_19 : _GEN_26; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_28 = 8'h14 == _match_key_bytes_23_T[7:0] ? phv_data_20 : _GEN_27; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_29 = 8'h15 == _match_key_bytes_23_T[7:0] ? phv_data_21 : _GEN_28; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_30 = 8'h16 == _match_key_bytes_23_T[7:0] ? phv_data_22 : _GEN_29; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_31 = 8'h17 == _match_key_bytes_23_T[7:0] ? phv_data_23 : _GEN_30; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_32 = 8'h18 == _match_key_bytes_23_T[7:0] ? phv_data_24 : _GEN_31; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_33 = 8'h19 == _match_key_bytes_23_T[7:0] ? phv_data_25 : _GEN_32; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_34 = 8'h1a == _match_key_bytes_23_T[7:0] ? phv_data_26 : _GEN_33; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_35 = 8'h1b == _match_key_bytes_23_T[7:0] ? phv_data_27 : _GEN_34; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_36 = 8'h1c == _match_key_bytes_23_T[7:0] ? phv_data_28 : _GEN_35; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_37 = 8'h1d == _match_key_bytes_23_T[7:0] ? phv_data_29 : _GEN_36; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_38 = 8'h1e == _match_key_bytes_23_T[7:0] ? phv_data_30 : _GEN_37; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_39 = 8'h1f == _match_key_bytes_23_T[7:0] ? phv_data_31 : _GEN_38; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_40 = 8'h20 == _match_key_bytes_23_T[7:0] ? phv_data_32 : _GEN_39; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_41 = 8'h21 == _match_key_bytes_23_T[7:0] ? phv_data_33 : _GEN_40; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_42 = 8'h22 == _match_key_bytes_23_T[7:0] ? phv_data_34 : _GEN_41; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_43 = 8'h23 == _match_key_bytes_23_T[7:0] ? phv_data_35 : _GEN_42; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_44 = 8'h24 == _match_key_bytes_23_T[7:0] ? phv_data_36 : _GEN_43; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_45 = 8'h25 == _match_key_bytes_23_T[7:0] ? phv_data_37 : _GEN_44; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_46 = 8'h26 == _match_key_bytes_23_T[7:0] ? phv_data_38 : _GEN_45; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_47 = 8'h27 == _match_key_bytes_23_T[7:0] ? phv_data_39 : _GEN_46; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_48 = 8'h28 == _match_key_bytes_23_T[7:0] ? phv_data_40 : _GEN_47; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_49 = 8'h29 == _match_key_bytes_23_T[7:0] ? phv_data_41 : _GEN_48; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_50 = 8'h2a == _match_key_bytes_23_T[7:0] ? phv_data_42 : _GEN_49; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_51 = 8'h2b == _match_key_bytes_23_T[7:0] ? phv_data_43 : _GEN_50; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_52 = 8'h2c == _match_key_bytes_23_T[7:0] ? phv_data_44 : _GEN_51; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_53 = 8'h2d == _match_key_bytes_23_T[7:0] ? phv_data_45 : _GEN_52; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_54 = 8'h2e == _match_key_bytes_23_T[7:0] ? phv_data_46 : _GEN_53; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_55 = 8'h2f == _match_key_bytes_23_T[7:0] ? phv_data_47 : _GEN_54; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_56 = 8'h30 == _match_key_bytes_23_T[7:0] ? phv_data_48 : _GEN_55; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_57 = 8'h31 == _match_key_bytes_23_T[7:0] ? phv_data_49 : _GEN_56; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_58 = 8'h32 == _match_key_bytes_23_T[7:0] ? phv_data_50 : _GEN_57; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_59 = 8'h33 == _match_key_bytes_23_T[7:0] ? phv_data_51 : _GEN_58; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_60 = 8'h34 == _match_key_bytes_23_T[7:0] ? phv_data_52 : _GEN_59; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_61 = 8'h35 == _match_key_bytes_23_T[7:0] ? phv_data_53 : _GEN_60; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_62 = 8'h36 == _match_key_bytes_23_T[7:0] ? phv_data_54 : _GEN_61; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_63 = 8'h37 == _match_key_bytes_23_T[7:0] ? phv_data_55 : _GEN_62; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_64 = 8'h38 == _match_key_bytes_23_T[7:0] ? phv_data_56 : _GEN_63; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_65 = 8'h39 == _match_key_bytes_23_T[7:0] ? phv_data_57 : _GEN_64; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_66 = 8'h3a == _match_key_bytes_23_T[7:0] ? phv_data_58 : _GEN_65; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_67 = 8'h3b == _match_key_bytes_23_T[7:0] ? phv_data_59 : _GEN_66; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_68 = 8'h3c == _match_key_bytes_23_T[7:0] ? phv_data_60 : _GEN_67; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_69 = 8'h3d == _match_key_bytes_23_T[7:0] ? phv_data_61 : _GEN_68; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_70 = 8'h3e == _match_key_bytes_23_T[7:0] ? phv_data_62 : _GEN_69; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_71 = 8'h3f == _match_key_bytes_23_T[7:0] ? phv_data_63 : _GEN_70; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_72 = 8'h40 == _match_key_bytes_23_T[7:0] ? phv_data_64 : _GEN_71; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_73 = 8'h41 == _match_key_bytes_23_T[7:0] ? phv_data_65 : _GEN_72; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_74 = 8'h42 == _match_key_bytes_23_T[7:0] ? phv_data_66 : _GEN_73; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_75 = 8'h43 == _match_key_bytes_23_T[7:0] ? phv_data_67 : _GEN_74; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_76 = 8'h44 == _match_key_bytes_23_T[7:0] ? phv_data_68 : _GEN_75; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_77 = 8'h45 == _match_key_bytes_23_T[7:0] ? phv_data_69 : _GEN_76; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_78 = 8'h46 == _match_key_bytes_23_T[7:0] ? phv_data_70 : _GEN_77; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_79 = 8'h47 == _match_key_bytes_23_T[7:0] ? phv_data_71 : _GEN_78; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_80 = 8'h48 == _match_key_bytes_23_T[7:0] ? phv_data_72 : _GEN_79; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_81 = 8'h49 == _match_key_bytes_23_T[7:0] ? phv_data_73 : _GEN_80; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_82 = 8'h4a == _match_key_bytes_23_T[7:0] ? phv_data_74 : _GEN_81; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_83 = 8'h4b == _match_key_bytes_23_T[7:0] ? phv_data_75 : _GEN_82; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_84 = 8'h4c == _match_key_bytes_23_T[7:0] ? phv_data_76 : _GEN_83; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_85 = 8'h4d == _match_key_bytes_23_T[7:0] ? phv_data_77 : _GEN_84; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_86 = 8'h4e == _match_key_bytes_23_T[7:0] ? phv_data_78 : _GEN_85; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_87 = 8'h4f == _match_key_bytes_23_T[7:0] ? phv_data_79 : _GEN_86; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_88 = 8'h50 == _match_key_bytes_23_T[7:0] ? phv_data_80 : _GEN_87; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_89 = 8'h51 == _match_key_bytes_23_T[7:0] ? phv_data_81 : _GEN_88; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_90 = 8'h52 == _match_key_bytes_23_T[7:0] ? phv_data_82 : _GEN_89; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_91 = 8'h53 == _match_key_bytes_23_T[7:0] ? phv_data_83 : _GEN_90; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_92 = 8'h54 == _match_key_bytes_23_T[7:0] ? phv_data_84 : _GEN_91; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_93 = 8'h55 == _match_key_bytes_23_T[7:0] ? phv_data_85 : _GEN_92; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_94 = 8'h56 == _match_key_bytes_23_T[7:0] ? phv_data_86 : _GEN_93; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_95 = 8'h57 == _match_key_bytes_23_T[7:0] ? phv_data_87 : _GEN_94; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_96 = 8'h58 == _match_key_bytes_23_T[7:0] ? phv_data_88 : _GEN_95; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_97 = 8'h59 == _match_key_bytes_23_T[7:0] ? phv_data_89 : _GEN_96; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_98 = 8'h5a == _match_key_bytes_23_T[7:0] ? phv_data_90 : _GEN_97; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_99 = 8'h5b == _match_key_bytes_23_T[7:0] ? phv_data_91 : _GEN_98; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_100 = 8'h5c == _match_key_bytes_23_T[7:0] ? phv_data_92 : _GEN_99; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_101 = 8'h5d == _match_key_bytes_23_T[7:0] ? phv_data_93 : _GEN_100; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_102 = 8'h5e == _match_key_bytes_23_T[7:0] ? phv_data_94 : _GEN_101; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_103 = 8'h5f == _match_key_bytes_23_T[7:0] ? phv_data_95 : _GEN_102; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_104 = 8'h60 == _match_key_bytes_23_T[7:0] ? phv_data_96 : _GEN_103; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_105 = 8'h61 == _match_key_bytes_23_T[7:0] ? phv_data_97 : _GEN_104; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_106 = 8'h62 == _match_key_bytes_23_T[7:0] ? phv_data_98 : _GEN_105; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_107 = 8'h63 == _match_key_bytes_23_T[7:0] ? phv_data_99 : _GEN_106; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_108 = 8'h64 == _match_key_bytes_23_T[7:0] ? phv_data_100 : _GEN_107; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_109 = 8'h65 == _match_key_bytes_23_T[7:0] ? phv_data_101 : _GEN_108; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_110 = 8'h66 == _match_key_bytes_23_T[7:0] ? phv_data_102 : _GEN_109; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_111 = 8'h67 == _match_key_bytes_23_T[7:0] ? phv_data_103 : _GEN_110; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_112 = 8'h68 == _match_key_bytes_23_T[7:0] ? phv_data_104 : _GEN_111; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_113 = 8'h69 == _match_key_bytes_23_T[7:0] ? phv_data_105 : _GEN_112; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_114 = 8'h6a == _match_key_bytes_23_T[7:0] ? phv_data_106 : _GEN_113; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_115 = 8'h6b == _match_key_bytes_23_T[7:0] ? phv_data_107 : _GEN_114; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_116 = 8'h6c == _match_key_bytes_23_T[7:0] ? phv_data_108 : _GEN_115; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_117 = 8'h6d == _match_key_bytes_23_T[7:0] ? phv_data_109 : _GEN_116; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_118 = 8'h6e == _match_key_bytes_23_T[7:0] ? phv_data_110 : _GEN_117; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_119 = 8'h6f == _match_key_bytes_23_T[7:0] ? phv_data_111 : _GEN_118; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_120 = 8'h70 == _match_key_bytes_23_T[7:0] ? phv_data_112 : _GEN_119; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_121 = 8'h71 == _match_key_bytes_23_T[7:0] ? phv_data_113 : _GEN_120; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_122 = 8'h72 == _match_key_bytes_23_T[7:0] ? phv_data_114 : _GEN_121; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_123 = 8'h73 == _match_key_bytes_23_T[7:0] ? phv_data_115 : _GEN_122; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_124 = 8'h74 == _match_key_bytes_23_T[7:0] ? phv_data_116 : _GEN_123; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_125 = 8'h75 == _match_key_bytes_23_T[7:0] ? phv_data_117 : _GEN_124; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_126 = 8'h76 == _match_key_bytes_23_T[7:0] ? phv_data_118 : _GEN_125; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_127 = 8'h77 == _match_key_bytes_23_T[7:0] ? phv_data_119 : _GEN_126; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_128 = 8'h78 == _match_key_bytes_23_T[7:0] ? phv_data_120 : _GEN_127; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_129 = 8'h79 == _match_key_bytes_23_T[7:0] ? phv_data_121 : _GEN_128; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_130 = 8'h7a == _match_key_bytes_23_T[7:0] ? phv_data_122 : _GEN_129; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_131 = 8'h7b == _match_key_bytes_23_T[7:0] ? phv_data_123 : _GEN_130; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_132 = 8'h7c == _match_key_bytes_23_T[7:0] ? phv_data_124 : _GEN_131; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_133 = 8'h7d == _match_key_bytes_23_T[7:0] ? phv_data_125 : _GEN_132; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_134 = 8'h7e == _match_key_bytes_23_T[7:0] ? phv_data_126 : _GEN_133; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_135 = 8'h7f == _match_key_bytes_23_T[7:0] ? phv_data_127 : _GEN_134; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_136 = 8'h80 == _match_key_bytes_23_T[7:0] ? phv_data_128 : _GEN_135; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_137 = 8'h81 == _match_key_bytes_23_T[7:0] ? phv_data_129 : _GEN_136; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_138 = 8'h82 == _match_key_bytes_23_T[7:0] ? phv_data_130 : _GEN_137; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_139 = 8'h83 == _match_key_bytes_23_T[7:0] ? phv_data_131 : _GEN_138; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_140 = 8'h84 == _match_key_bytes_23_T[7:0] ? phv_data_132 : _GEN_139; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_141 = 8'h85 == _match_key_bytes_23_T[7:0] ? phv_data_133 : _GEN_140; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_142 = 8'h86 == _match_key_bytes_23_T[7:0] ? phv_data_134 : _GEN_141; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_143 = 8'h87 == _match_key_bytes_23_T[7:0] ? phv_data_135 : _GEN_142; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_144 = 8'h88 == _match_key_bytes_23_T[7:0] ? phv_data_136 : _GEN_143; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_145 = 8'h89 == _match_key_bytes_23_T[7:0] ? phv_data_137 : _GEN_144; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_146 = 8'h8a == _match_key_bytes_23_T[7:0] ? phv_data_138 : _GEN_145; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_147 = 8'h8b == _match_key_bytes_23_T[7:0] ? phv_data_139 : _GEN_146; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_148 = 8'h8c == _match_key_bytes_23_T[7:0] ? phv_data_140 : _GEN_147; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_149 = 8'h8d == _match_key_bytes_23_T[7:0] ? phv_data_141 : _GEN_148; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_150 = 8'h8e == _match_key_bytes_23_T[7:0] ? phv_data_142 : _GEN_149; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_151 = 8'h8f == _match_key_bytes_23_T[7:0] ? phv_data_143 : _GEN_150; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_152 = 8'h90 == _match_key_bytes_23_T[7:0] ? phv_data_144 : _GEN_151; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_153 = 8'h91 == _match_key_bytes_23_T[7:0] ? phv_data_145 : _GEN_152; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_154 = 8'h92 == _match_key_bytes_23_T[7:0] ? phv_data_146 : _GEN_153; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_155 = 8'h93 == _match_key_bytes_23_T[7:0] ? phv_data_147 : _GEN_154; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_156 = 8'h94 == _match_key_bytes_23_T[7:0] ? phv_data_148 : _GEN_155; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_157 = 8'h95 == _match_key_bytes_23_T[7:0] ? phv_data_149 : _GEN_156; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_158 = 8'h96 == _match_key_bytes_23_T[7:0] ? phv_data_150 : _GEN_157; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_159 = 8'h97 == _match_key_bytes_23_T[7:0] ? phv_data_151 : _GEN_158; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_160 = 8'h98 == _match_key_bytes_23_T[7:0] ? phv_data_152 : _GEN_159; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_161 = 8'h99 == _match_key_bytes_23_T[7:0] ? phv_data_153 : _GEN_160; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_162 = 8'h9a == _match_key_bytes_23_T[7:0] ? phv_data_154 : _GEN_161; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_163 = 8'h9b == _match_key_bytes_23_T[7:0] ? phv_data_155 : _GEN_162; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_164 = 8'h9c == _match_key_bytes_23_T[7:0] ? phv_data_156 : _GEN_163; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_165 = 8'h9d == _match_key_bytes_23_T[7:0] ? phv_data_157 : _GEN_164; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_166 = 8'h9e == _match_key_bytes_23_T[7:0] ? phv_data_158 : _GEN_165; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_167 = 8'h9f == _match_key_bytes_23_T[7:0] ? phv_data_159 : _GEN_166; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_23 = 8'h0 < _GEN_6 ? _GEN_167 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_22_T_1 = key_offset + 8'h1; // @[matcher.scala 72:98]
  wire [7:0] _GEN_170 = 8'h1 == _match_key_bytes_22_T_1 ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_171 = 8'h2 == _match_key_bytes_22_T_1 ? phv_data_2 : _GEN_170; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_172 = 8'h3 == _match_key_bytes_22_T_1 ? phv_data_3 : _GEN_171; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_173 = 8'h4 == _match_key_bytes_22_T_1 ? phv_data_4 : _GEN_172; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_174 = 8'h5 == _match_key_bytes_22_T_1 ? phv_data_5 : _GEN_173; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_175 = 8'h6 == _match_key_bytes_22_T_1 ? phv_data_6 : _GEN_174; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_176 = 8'h7 == _match_key_bytes_22_T_1 ? phv_data_7 : _GEN_175; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_177 = 8'h8 == _match_key_bytes_22_T_1 ? phv_data_8 : _GEN_176; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_178 = 8'h9 == _match_key_bytes_22_T_1 ? phv_data_9 : _GEN_177; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_179 = 8'ha == _match_key_bytes_22_T_1 ? phv_data_10 : _GEN_178; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_180 = 8'hb == _match_key_bytes_22_T_1 ? phv_data_11 : _GEN_179; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_181 = 8'hc == _match_key_bytes_22_T_1 ? phv_data_12 : _GEN_180; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_182 = 8'hd == _match_key_bytes_22_T_1 ? phv_data_13 : _GEN_181; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_183 = 8'he == _match_key_bytes_22_T_1 ? phv_data_14 : _GEN_182; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_184 = 8'hf == _match_key_bytes_22_T_1 ? phv_data_15 : _GEN_183; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_185 = 8'h10 == _match_key_bytes_22_T_1 ? phv_data_16 : _GEN_184; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_186 = 8'h11 == _match_key_bytes_22_T_1 ? phv_data_17 : _GEN_185; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_187 = 8'h12 == _match_key_bytes_22_T_1 ? phv_data_18 : _GEN_186; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_188 = 8'h13 == _match_key_bytes_22_T_1 ? phv_data_19 : _GEN_187; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_189 = 8'h14 == _match_key_bytes_22_T_1 ? phv_data_20 : _GEN_188; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_190 = 8'h15 == _match_key_bytes_22_T_1 ? phv_data_21 : _GEN_189; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_191 = 8'h16 == _match_key_bytes_22_T_1 ? phv_data_22 : _GEN_190; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_192 = 8'h17 == _match_key_bytes_22_T_1 ? phv_data_23 : _GEN_191; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_193 = 8'h18 == _match_key_bytes_22_T_1 ? phv_data_24 : _GEN_192; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_194 = 8'h19 == _match_key_bytes_22_T_1 ? phv_data_25 : _GEN_193; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_195 = 8'h1a == _match_key_bytes_22_T_1 ? phv_data_26 : _GEN_194; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_196 = 8'h1b == _match_key_bytes_22_T_1 ? phv_data_27 : _GEN_195; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_197 = 8'h1c == _match_key_bytes_22_T_1 ? phv_data_28 : _GEN_196; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_198 = 8'h1d == _match_key_bytes_22_T_1 ? phv_data_29 : _GEN_197; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_199 = 8'h1e == _match_key_bytes_22_T_1 ? phv_data_30 : _GEN_198; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_200 = 8'h1f == _match_key_bytes_22_T_1 ? phv_data_31 : _GEN_199; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_201 = 8'h20 == _match_key_bytes_22_T_1 ? phv_data_32 : _GEN_200; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_202 = 8'h21 == _match_key_bytes_22_T_1 ? phv_data_33 : _GEN_201; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_203 = 8'h22 == _match_key_bytes_22_T_1 ? phv_data_34 : _GEN_202; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_204 = 8'h23 == _match_key_bytes_22_T_1 ? phv_data_35 : _GEN_203; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_205 = 8'h24 == _match_key_bytes_22_T_1 ? phv_data_36 : _GEN_204; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_206 = 8'h25 == _match_key_bytes_22_T_1 ? phv_data_37 : _GEN_205; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_207 = 8'h26 == _match_key_bytes_22_T_1 ? phv_data_38 : _GEN_206; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_208 = 8'h27 == _match_key_bytes_22_T_1 ? phv_data_39 : _GEN_207; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_209 = 8'h28 == _match_key_bytes_22_T_1 ? phv_data_40 : _GEN_208; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_210 = 8'h29 == _match_key_bytes_22_T_1 ? phv_data_41 : _GEN_209; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_211 = 8'h2a == _match_key_bytes_22_T_1 ? phv_data_42 : _GEN_210; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_212 = 8'h2b == _match_key_bytes_22_T_1 ? phv_data_43 : _GEN_211; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_213 = 8'h2c == _match_key_bytes_22_T_1 ? phv_data_44 : _GEN_212; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_214 = 8'h2d == _match_key_bytes_22_T_1 ? phv_data_45 : _GEN_213; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_215 = 8'h2e == _match_key_bytes_22_T_1 ? phv_data_46 : _GEN_214; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_216 = 8'h2f == _match_key_bytes_22_T_1 ? phv_data_47 : _GEN_215; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_217 = 8'h30 == _match_key_bytes_22_T_1 ? phv_data_48 : _GEN_216; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_218 = 8'h31 == _match_key_bytes_22_T_1 ? phv_data_49 : _GEN_217; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_219 = 8'h32 == _match_key_bytes_22_T_1 ? phv_data_50 : _GEN_218; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_220 = 8'h33 == _match_key_bytes_22_T_1 ? phv_data_51 : _GEN_219; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_221 = 8'h34 == _match_key_bytes_22_T_1 ? phv_data_52 : _GEN_220; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_222 = 8'h35 == _match_key_bytes_22_T_1 ? phv_data_53 : _GEN_221; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_223 = 8'h36 == _match_key_bytes_22_T_1 ? phv_data_54 : _GEN_222; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_224 = 8'h37 == _match_key_bytes_22_T_1 ? phv_data_55 : _GEN_223; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_225 = 8'h38 == _match_key_bytes_22_T_1 ? phv_data_56 : _GEN_224; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_226 = 8'h39 == _match_key_bytes_22_T_1 ? phv_data_57 : _GEN_225; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_227 = 8'h3a == _match_key_bytes_22_T_1 ? phv_data_58 : _GEN_226; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_228 = 8'h3b == _match_key_bytes_22_T_1 ? phv_data_59 : _GEN_227; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_229 = 8'h3c == _match_key_bytes_22_T_1 ? phv_data_60 : _GEN_228; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_230 = 8'h3d == _match_key_bytes_22_T_1 ? phv_data_61 : _GEN_229; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_231 = 8'h3e == _match_key_bytes_22_T_1 ? phv_data_62 : _GEN_230; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_232 = 8'h3f == _match_key_bytes_22_T_1 ? phv_data_63 : _GEN_231; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_233 = 8'h40 == _match_key_bytes_22_T_1 ? phv_data_64 : _GEN_232; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_234 = 8'h41 == _match_key_bytes_22_T_1 ? phv_data_65 : _GEN_233; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_235 = 8'h42 == _match_key_bytes_22_T_1 ? phv_data_66 : _GEN_234; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_236 = 8'h43 == _match_key_bytes_22_T_1 ? phv_data_67 : _GEN_235; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_237 = 8'h44 == _match_key_bytes_22_T_1 ? phv_data_68 : _GEN_236; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_238 = 8'h45 == _match_key_bytes_22_T_1 ? phv_data_69 : _GEN_237; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_239 = 8'h46 == _match_key_bytes_22_T_1 ? phv_data_70 : _GEN_238; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_240 = 8'h47 == _match_key_bytes_22_T_1 ? phv_data_71 : _GEN_239; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_241 = 8'h48 == _match_key_bytes_22_T_1 ? phv_data_72 : _GEN_240; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_242 = 8'h49 == _match_key_bytes_22_T_1 ? phv_data_73 : _GEN_241; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_243 = 8'h4a == _match_key_bytes_22_T_1 ? phv_data_74 : _GEN_242; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_244 = 8'h4b == _match_key_bytes_22_T_1 ? phv_data_75 : _GEN_243; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_245 = 8'h4c == _match_key_bytes_22_T_1 ? phv_data_76 : _GEN_244; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_246 = 8'h4d == _match_key_bytes_22_T_1 ? phv_data_77 : _GEN_245; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_247 = 8'h4e == _match_key_bytes_22_T_1 ? phv_data_78 : _GEN_246; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_248 = 8'h4f == _match_key_bytes_22_T_1 ? phv_data_79 : _GEN_247; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_249 = 8'h50 == _match_key_bytes_22_T_1 ? phv_data_80 : _GEN_248; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_250 = 8'h51 == _match_key_bytes_22_T_1 ? phv_data_81 : _GEN_249; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_251 = 8'h52 == _match_key_bytes_22_T_1 ? phv_data_82 : _GEN_250; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_252 = 8'h53 == _match_key_bytes_22_T_1 ? phv_data_83 : _GEN_251; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_253 = 8'h54 == _match_key_bytes_22_T_1 ? phv_data_84 : _GEN_252; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_254 = 8'h55 == _match_key_bytes_22_T_1 ? phv_data_85 : _GEN_253; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_255 = 8'h56 == _match_key_bytes_22_T_1 ? phv_data_86 : _GEN_254; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_256 = 8'h57 == _match_key_bytes_22_T_1 ? phv_data_87 : _GEN_255; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_257 = 8'h58 == _match_key_bytes_22_T_1 ? phv_data_88 : _GEN_256; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_258 = 8'h59 == _match_key_bytes_22_T_1 ? phv_data_89 : _GEN_257; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_259 = 8'h5a == _match_key_bytes_22_T_1 ? phv_data_90 : _GEN_258; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_260 = 8'h5b == _match_key_bytes_22_T_1 ? phv_data_91 : _GEN_259; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_261 = 8'h5c == _match_key_bytes_22_T_1 ? phv_data_92 : _GEN_260; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_262 = 8'h5d == _match_key_bytes_22_T_1 ? phv_data_93 : _GEN_261; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_263 = 8'h5e == _match_key_bytes_22_T_1 ? phv_data_94 : _GEN_262; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_264 = 8'h5f == _match_key_bytes_22_T_1 ? phv_data_95 : _GEN_263; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_265 = 8'h60 == _match_key_bytes_22_T_1 ? phv_data_96 : _GEN_264; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_266 = 8'h61 == _match_key_bytes_22_T_1 ? phv_data_97 : _GEN_265; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_267 = 8'h62 == _match_key_bytes_22_T_1 ? phv_data_98 : _GEN_266; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_268 = 8'h63 == _match_key_bytes_22_T_1 ? phv_data_99 : _GEN_267; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_269 = 8'h64 == _match_key_bytes_22_T_1 ? phv_data_100 : _GEN_268; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_270 = 8'h65 == _match_key_bytes_22_T_1 ? phv_data_101 : _GEN_269; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_271 = 8'h66 == _match_key_bytes_22_T_1 ? phv_data_102 : _GEN_270; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_272 = 8'h67 == _match_key_bytes_22_T_1 ? phv_data_103 : _GEN_271; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_273 = 8'h68 == _match_key_bytes_22_T_1 ? phv_data_104 : _GEN_272; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_274 = 8'h69 == _match_key_bytes_22_T_1 ? phv_data_105 : _GEN_273; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_275 = 8'h6a == _match_key_bytes_22_T_1 ? phv_data_106 : _GEN_274; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_276 = 8'h6b == _match_key_bytes_22_T_1 ? phv_data_107 : _GEN_275; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_277 = 8'h6c == _match_key_bytes_22_T_1 ? phv_data_108 : _GEN_276; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_278 = 8'h6d == _match_key_bytes_22_T_1 ? phv_data_109 : _GEN_277; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_279 = 8'h6e == _match_key_bytes_22_T_1 ? phv_data_110 : _GEN_278; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_280 = 8'h6f == _match_key_bytes_22_T_1 ? phv_data_111 : _GEN_279; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_281 = 8'h70 == _match_key_bytes_22_T_1 ? phv_data_112 : _GEN_280; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_282 = 8'h71 == _match_key_bytes_22_T_1 ? phv_data_113 : _GEN_281; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_283 = 8'h72 == _match_key_bytes_22_T_1 ? phv_data_114 : _GEN_282; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_284 = 8'h73 == _match_key_bytes_22_T_1 ? phv_data_115 : _GEN_283; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_285 = 8'h74 == _match_key_bytes_22_T_1 ? phv_data_116 : _GEN_284; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_286 = 8'h75 == _match_key_bytes_22_T_1 ? phv_data_117 : _GEN_285; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_287 = 8'h76 == _match_key_bytes_22_T_1 ? phv_data_118 : _GEN_286; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_288 = 8'h77 == _match_key_bytes_22_T_1 ? phv_data_119 : _GEN_287; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_289 = 8'h78 == _match_key_bytes_22_T_1 ? phv_data_120 : _GEN_288; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_290 = 8'h79 == _match_key_bytes_22_T_1 ? phv_data_121 : _GEN_289; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_291 = 8'h7a == _match_key_bytes_22_T_1 ? phv_data_122 : _GEN_290; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_292 = 8'h7b == _match_key_bytes_22_T_1 ? phv_data_123 : _GEN_291; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_293 = 8'h7c == _match_key_bytes_22_T_1 ? phv_data_124 : _GEN_292; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_294 = 8'h7d == _match_key_bytes_22_T_1 ? phv_data_125 : _GEN_293; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_295 = 8'h7e == _match_key_bytes_22_T_1 ? phv_data_126 : _GEN_294; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_296 = 8'h7f == _match_key_bytes_22_T_1 ? phv_data_127 : _GEN_295; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_297 = 8'h80 == _match_key_bytes_22_T_1 ? phv_data_128 : _GEN_296; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_298 = 8'h81 == _match_key_bytes_22_T_1 ? phv_data_129 : _GEN_297; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_299 = 8'h82 == _match_key_bytes_22_T_1 ? phv_data_130 : _GEN_298; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_300 = 8'h83 == _match_key_bytes_22_T_1 ? phv_data_131 : _GEN_299; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_301 = 8'h84 == _match_key_bytes_22_T_1 ? phv_data_132 : _GEN_300; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_302 = 8'h85 == _match_key_bytes_22_T_1 ? phv_data_133 : _GEN_301; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_303 = 8'h86 == _match_key_bytes_22_T_1 ? phv_data_134 : _GEN_302; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_304 = 8'h87 == _match_key_bytes_22_T_1 ? phv_data_135 : _GEN_303; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_305 = 8'h88 == _match_key_bytes_22_T_1 ? phv_data_136 : _GEN_304; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_306 = 8'h89 == _match_key_bytes_22_T_1 ? phv_data_137 : _GEN_305; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_307 = 8'h8a == _match_key_bytes_22_T_1 ? phv_data_138 : _GEN_306; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_308 = 8'h8b == _match_key_bytes_22_T_1 ? phv_data_139 : _GEN_307; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_309 = 8'h8c == _match_key_bytes_22_T_1 ? phv_data_140 : _GEN_308; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_310 = 8'h8d == _match_key_bytes_22_T_1 ? phv_data_141 : _GEN_309; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_311 = 8'h8e == _match_key_bytes_22_T_1 ? phv_data_142 : _GEN_310; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_312 = 8'h8f == _match_key_bytes_22_T_1 ? phv_data_143 : _GEN_311; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_313 = 8'h90 == _match_key_bytes_22_T_1 ? phv_data_144 : _GEN_312; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_314 = 8'h91 == _match_key_bytes_22_T_1 ? phv_data_145 : _GEN_313; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_315 = 8'h92 == _match_key_bytes_22_T_1 ? phv_data_146 : _GEN_314; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_316 = 8'h93 == _match_key_bytes_22_T_1 ? phv_data_147 : _GEN_315; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_317 = 8'h94 == _match_key_bytes_22_T_1 ? phv_data_148 : _GEN_316; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_318 = 8'h95 == _match_key_bytes_22_T_1 ? phv_data_149 : _GEN_317; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_319 = 8'h96 == _match_key_bytes_22_T_1 ? phv_data_150 : _GEN_318; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_320 = 8'h97 == _match_key_bytes_22_T_1 ? phv_data_151 : _GEN_319; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_321 = 8'h98 == _match_key_bytes_22_T_1 ? phv_data_152 : _GEN_320; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_322 = 8'h99 == _match_key_bytes_22_T_1 ? phv_data_153 : _GEN_321; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_323 = 8'h9a == _match_key_bytes_22_T_1 ? phv_data_154 : _GEN_322; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_324 = 8'h9b == _match_key_bytes_22_T_1 ? phv_data_155 : _GEN_323; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_325 = 8'h9c == _match_key_bytes_22_T_1 ? phv_data_156 : _GEN_324; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_326 = 8'h9d == _match_key_bytes_22_T_1 ? phv_data_157 : _GEN_325; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_327 = 8'h9e == _match_key_bytes_22_T_1 ? phv_data_158 : _GEN_326; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_328 = 8'h9f == _match_key_bytes_22_T_1 ? phv_data_159 : _GEN_327; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_22 = 8'h1 < _GEN_6 ? _GEN_328 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_21_T_1 = key_offset + 8'h2; // @[matcher.scala 72:98]
  wire [7:0] _GEN_331 = 8'h1 == _match_key_bytes_21_T_1 ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_332 = 8'h2 == _match_key_bytes_21_T_1 ? phv_data_2 : _GEN_331; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_333 = 8'h3 == _match_key_bytes_21_T_1 ? phv_data_3 : _GEN_332; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_334 = 8'h4 == _match_key_bytes_21_T_1 ? phv_data_4 : _GEN_333; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_335 = 8'h5 == _match_key_bytes_21_T_1 ? phv_data_5 : _GEN_334; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_336 = 8'h6 == _match_key_bytes_21_T_1 ? phv_data_6 : _GEN_335; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_337 = 8'h7 == _match_key_bytes_21_T_1 ? phv_data_7 : _GEN_336; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_338 = 8'h8 == _match_key_bytes_21_T_1 ? phv_data_8 : _GEN_337; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_339 = 8'h9 == _match_key_bytes_21_T_1 ? phv_data_9 : _GEN_338; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_340 = 8'ha == _match_key_bytes_21_T_1 ? phv_data_10 : _GEN_339; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_341 = 8'hb == _match_key_bytes_21_T_1 ? phv_data_11 : _GEN_340; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_342 = 8'hc == _match_key_bytes_21_T_1 ? phv_data_12 : _GEN_341; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_343 = 8'hd == _match_key_bytes_21_T_1 ? phv_data_13 : _GEN_342; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_344 = 8'he == _match_key_bytes_21_T_1 ? phv_data_14 : _GEN_343; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_345 = 8'hf == _match_key_bytes_21_T_1 ? phv_data_15 : _GEN_344; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_346 = 8'h10 == _match_key_bytes_21_T_1 ? phv_data_16 : _GEN_345; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_347 = 8'h11 == _match_key_bytes_21_T_1 ? phv_data_17 : _GEN_346; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_348 = 8'h12 == _match_key_bytes_21_T_1 ? phv_data_18 : _GEN_347; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_349 = 8'h13 == _match_key_bytes_21_T_1 ? phv_data_19 : _GEN_348; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_350 = 8'h14 == _match_key_bytes_21_T_1 ? phv_data_20 : _GEN_349; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_351 = 8'h15 == _match_key_bytes_21_T_1 ? phv_data_21 : _GEN_350; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_352 = 8'h16 == _match_key_bytes_21_T_1 ? phv_data_22 : _GEN_351; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_353 = 8'h17 == _match_key_bytes_21_T_1 ? phv_data_23 : _GEN_352; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_354 = 8'h18 == _match_key_bytes_21_T_1 ? phv_data_24 : _GEN_353; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_355 = 8'h19 == _match_key_bytes_21_T_1 ? phv_data_25 : _GEN_354; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_356 = 8'h1a == _match_key_bytes_21_T_1 ? phv_data_26 : _GEN_355; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_357 = 8'h1b == _match_key_bytes_21_T_1 ? phv_data_27 : _GEN_356; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_358 = 8'h1c == _match_key_bytes_21_T_1 ? phv_data_28 : _GEN_357; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_359 = 8'h1d == _match_key_bytes_21_T_1 ? phv_data_29 : _GEN_358; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_360 = 8'h1e == _match_key_bytes_21_T_1 ? phv_data_30 : _GEN_359; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_361 = 8'h1f == _match_key_bytes_21_T_1 ? phv_data_31 : _GEN_360; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_362 = 8'h20 == _match_key_bytes_21_T_1 ? phv_data_32 : _GEN_361; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_363 = 8'h21 == _match_key_bytes_21_T_1 ? phv_data_33 : _GEN_362; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_364 = 8'h22 == _match_key_bytes_21_T_1 ? phv_data_34 : _GEN_363; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_365 = 8'h23 == _match_key_bytes_21_T_1 ? phv_data_35 : _GEN_364; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_366 = 8'h24 == _match_key_bytes_21_T_1 ? phv_data_36 : _GEN_365; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_367 = 8'h25 == _match_key_bytes_21_T_1 ? phv_data_37 : _GEN_366; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_368 = 8'h26 == _match_key_bytes_21_T_1 ? phv_data_38 : _GEN_367; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_369 = 8'h27 == _match_key_bytes_21_T_1 ? phv_data_39 : _GEN_368; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_370 = 8'h28 == _match_key_bytes_21_T_1 ? phv_data_40 : _GEN_369; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_371 = 8'h29 == _match_key_bytes_21_T_1 ? phv_data_41 : _GEN_370; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_372 = 8'h2a == _match_key_bytes_21_T_1 ? phv_data_42 : _GEN_371; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_373 = 8'h2b == _match_key_bytes_21_T_1 ? phv_data_43 : _GEN_372; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_374 = 8'h2c == _match_key_bytes_21_T_1 ? phv_data_44 : _GEN_373; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_375 = 8'h2d == _match_key_bytes_21_T_1 ? phv_data_45 : _GEN_374; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_376 = 8'h2e == _match_key_bytes_21_T_1 ? phv_data_46 : _GEN_375; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_377 = 8'h2f == _match_key_bytes_21_T_1 ? phv_data_47 : _GEN_376; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_378 = 8'h30 == _match_key_bytes_21_T_1 ? phv_data_48 : _GEN_377; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_379 = 8'h31 == _match_key_bytes_21_T_1 ? phv_data_49 : _GEN_378; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_380 = 8'h32 == _match_key_bytes_21_T_1 ? phv_data_50 : _GEN_379; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_381 = 8'h33 == _match_key_bytes_21_T_1 ? phv_data_51 : _GEN_380; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_382 = 8'h34 == _match_key_bytes_21_T_1 ? phv_data_52 : _GEN_381; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_383 = 8'h35 == _match_key_bytes_21_T_1 ? phv_data_53 : _GEN_382; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_384 = 8'h36 == _match_key_bytes_21_T_1 ? phv_data_54 : _GEN_383; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_385 = 8'h37 == _match_key_bytes_21_T_1 ? phv_data_55 : _GEN_384; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_386 = 8'h38 == _match_key_bytes_21_T_1 ? phv_data_56 : _GEN_385; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_387 = 8'h39 == _match_key_bytes_21_T_1 ? phv_data_57 : _GEN_386; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_388 = 8'h3a == _match_key_bytes_21_T_1 ? phv_data_58 : _GEN_387; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_389 = 8'h3b == _match_key_bytes_21_T_1 ? phv_data_59 : _GEN_388; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_390 = 8'h3c == _match_key_bytes_21_T_1 ? phv_data_60 : _GEN_389; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_391 = 8'h3d == _match_key_bytes_21_T_1 ? phv_data_61 : _GEN_390; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_392 = 8'h3e == _match_key_bytes_21_T_1 ? phv_data_62 : _GEN_391; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_393 = 8'h3f == _match_key_bytes_21_T_1 ? phv_data_63 : _GEN_392; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_394 = 8'h40 == _match_key_bytes_21_T_1 ? phv_data_64 : _GEN_393; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_395 = 8'h41 == _match_key_bytes_21_T_1 ? phv_data_65 : _GEN_394; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_396 = 8'h42 == _match_key_bytes_21_T_1 ? phv_data_66 : _GEN_395; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_397 = 8'h43 == _match_key_bytes_21_T_1 ? phv_data_67 : _GEN_396; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_398 = 8'h44 == _match_key_bytes_21_T_1 ? phv_data_68 : _GEN_397; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_399 = 8'h45 == _match_key_bytes_21_T_1 ? phv_data_69 : _GEN_398; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_400 = 8'h46 == _match_key_bytes_21_T_1 ? phv_data_70 : _GEN_399; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_401 = 8'h47 == _match_key_bytes_21_T_1 ? phv_data_71 : _GEN_400; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_402 = 8'h48 == _match_key_bytes_21_T_1 ? phv_data_72 : _GEN_401; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_403 = 8'h49 == _match_key_bytes_21_T_1 ? phv_data_73 : _GEN_402; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_404 = 8'h4a == _match_key_bytes_21_T_1 ? phv_data_74 : _GEN_403; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_405 = 8'h4b == _match_key_bytes_21_T_1 ? phv_data_75 : _GEN_404; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_406 = 8'h4c == _match_key_bytes_21_T_1 ? phv_data_76 : _GEN_405; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_407 = 8'h4d == _match_key_bytes_21_T_1 ? phv_data_77 : _GEN_406; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_408 = 8'h4e == _match_key_bytes_21_T_1 ? phv_data_78 : _GEN_407; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_409 = 8'h4f == _match_key_bytes_21_T_1 ? phv_data_79 : _GEN_408; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_410 = 8'h50 == _match_key_bytes_21_T_1 ? phv_data_80 : _GEN_409; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_411 = 8'h51 == _match_key_bytes_21_T_1 ? phv_data_81 : _GEN_410; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_412 = 8'h52 == _match_key_bytes_21_T_1 ? phv_data_82 : _GEN_411; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_413 = 8'h53 == _match_key_bytes_21_T_1 ? phv_data_83 : _GEN_412; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_414 = 8'h54 == _match_key_bytes_21_T_1 ? phv_data_84 : _GEN_413; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_415 = 8'h55 == _match_key_bytes_21_T_1 ? phv_data_85 : _GEN_414; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_416 = 8'h56 == _match_key_bytes_21_T_1 ? phv_data_86 : _GEN_415; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_417 = 8'h57 == _match_key_bytes_21_T_1 ? phv_data_87 : _GEN_416; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_418 = 8'h58 == _match_key_bytes_21_T_1 ? phv_data_88 : _GEN_417; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_419 = 8'h59 == _match_key_bytes_21_T_1 ? phv_data_89 : _GEN_418; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_420 = 8'h5a == _match_key_bytes_21_T_1 ? phv_data_90 : _GEN_419; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_421 = 8'h5b == _match_key_bytes_21_T_1 ? phv_data_91 : _GEN_420; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_422 = 8'h5c == _match_key_bytes_21_T_1 ? phv_data_92 : _GEN_421; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_423 = 8'h5d == _match_key_bytes_21_T_1 ? phv_data_93 : _GEN_422; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_424 = 8'h5e == _match_key_bytes_21_T_1 ? phv_data_94 : _GEN_423; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_425 = 8'h5f == _match_key_bytes_21_T_1 ? phv_data_95 : _GEN_424; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_426 = 8'h60 == _match_key_bytes_21_T_1 ? phv_data_96 : _GEN_425; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_427 = 8'h61 == _match_key_bytes_21_T_1 ? phv_data_97 : _GEN_426; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_428 = 8'h62 == _match_key_bytes_21_T_1 ? phv_data_98 : _GEN_427; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_429 = 8'h63 == _match_key_bytes_21_T_1 ? phv_data_99 : _GEN_428; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_430 = 8'h64 == _match_key_bytes_21_T_1 ? phv_data_100 : _GEN_429; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_431 = 8'h65 == _match_key_bytes_21_T_1 ? phv_data_101 : _GEN_430; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_432 = 8'h66 == _match_key_bytes_21_T_1 ? phv_data_102 : _GEN_431; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_433 = 8'h67 == _match_key_bytes_21_T_1 ? phv_data_103 : _GEN_432; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_434 = 8'h68 == _match_key_bytes_21_T_1 ? phv_data_104 : _GEN_433; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_435 = 8'h69 == _match_key_bytes_21_T_1 ? phv_data_105 : _GEN_434; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_436 = 8'h6a == _match_key_bytes_21_T_1 ? phv_data_106 : _GEN_435; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_437 = 8'h6b == _match_key_bytes_21_T_1 ? phv_data_107 : _GEN_436; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_438 = 8'h6c == _match_key_bytes_21_T_1 ? phv_data_108 : _GEN_437; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_439 = 8'h6d == _match_key_bytes_21_T_1 ? phv_data_109 : _GEN_438; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_440 = 8'h6e == _match_key_bytes_21_T_1 ? phv_data_110 : _GEN_439; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_441 = 8'h6f == _match_key_bytes_21_T_1 ? phv_data_111 : _GEN_440; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_442 = 8'h70 == _match_key_bytes_21_T_1 ? phv_data_112 : _GEN_441; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_443 = 8'h71 == _match_key_bytes_21_T_1 ? phv_data_113 : _GEN_442; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_444 = 8'h72 == _match_key_bytes_21_T_1 ? phv_data_114 : _GEN_443; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_445 = 8'h73 == _match_key_bytes_21_T_1 ? phv_data_115 : _GEN_444; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_446 = 8'h74 == _match_key_bytes_21_T_1 ? phv_data_116 : _GEN_445; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_447 = 8'h75 == _match_key_bytes_21_T_1 ? phv_data_117 : _GEN_446; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_448 = 8'h76 == _match_key_bytes_21_T_1 ? phv_data_118 : _GEN_447; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_449 = 8'h77 == _match_key_bytes_21_T_1 ? phv_data_119 : _GEN_448; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_450 = 8'h78 == _match_key_bytes_21_T_1 ? phv_data_120 : _GEN_449; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_451 = 8'h79 == _match_key_bytes_21_T_1 ? phv_data_121 : _GEN_450; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_452 = 8'h7a == _match_key_bytes_21_T_1 ? phv_data_122 : _GEN_451; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_453 = 8'h7b == _match_key_bytes_21_T_1 ? phv_data_123 : _GEN_452; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_454 = 8'h7c == _match_key_bytes_21_T_1 ? phv_data_124 : _GEN_453; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_455 = 8'h7d == _match_key_bytes_21_T_1 ? phv_data_125 : _GEN_454; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_456 = 8'h7e == _match_key_bytes_21_T_1 ? phv_data_126 : _GEN_455; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_457 = 8'h7f == _match_key_bytes_21_T_1 ? phv_data_127 : _GEN_456; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_458 = 8'h80 == _match_key_bytes_21_T_1 ? phv_data_128 : _GEN_457; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_459 = 8'h81 == _match_key_bytes_21_T_1 ? phv_data_129 : _GEN_458; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_460 = 8'h82 == _match_key_bytes_21_T_1 ? phv_data_130 : _GEN_459; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_461 = 8'h83 == _match_key_bytes_21_T_1 ? phv_data_131 : _GEN_460; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_462 = 8'h84 == _match_key_bytes_21_T_1 ? phv_data_132 : _GEN_461; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_463 = 8'h85 == _match_key_bytes_21_T_1 ? phv_data_133 : _GEN_462; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_464 = 8'h86 == _match_key_bytes_21_T_1 ? phv_data_134 : _GEN_463; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_465 = 8'h87 == _match_key_bytes_21_T_1 ? phv_data_135 : _GEN_464; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_466 = 8'h88 == _match_key_bytes_21_T_1 ? phv_data_136 : _GEN_465; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_467 = 8'h89 == _match_key_bytes_21_T_1 ? phv_data_137 : _GEN_466; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_468 = 8'h8a == _match_key_bytes_21_T_1 ? phv_data_138 : _GEN_467; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_469 = 8'h8b == _match_key_bytes_21_T_1 ? phv_data_139 : _GEN_468; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_470 = 8'h8c == _match_key_bytes_21_T_1 ? phv_data_140 : _GEN_469; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_471 = 8'h8d == _match_key_bytes_21_T_1 ? phv_data_141 : _GEN_470; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_472 = 8'h8e == _match_key_bytes_21_T_1 ? phv_data_142 : _GEN_471; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_473 = 8'h8f == _match_key_bytes_21_T_1 ? phv_data_143 : _GEN_472; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_474 = 8'h90 == _match_key_bytes_21_T_1 ? phv_data_144 : _GEN_473; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_475 = 8'h91 == _match_key_bytes_21_T_1 ? phv_data_145 : _GEN_474; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_476 = 8'h92 == _match_key_bytes_21_T_1 ? phv_data_146 : _GEN_475; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_477 = 8'h93 == _match_key_bytes_21_T_1 ? phv_data_147 : _GEN_476; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_478 = 8'h94 == _match_key_bytes_21_T_1 ? phv_data_148 : _GEN_477; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_479 = 8'h95 == _match_key_bytes_21_T_1 ? phv_data_149 : _GEN_478; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_480 = 8'h96 == _match_key_bytes_21_T_1 ? phv_data_150 : _GEN_479; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_481 = 8'h97 == _match_key_bytes_21_T_1 ? phv_data_151 : _GEN_480; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_482 = 8'h98 == _match_key_bytes_21_T_1 ? phv_data_152 : _GEN_481; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_483 = 8'h99 == _match_key_bytes_21_T_1 ? phv_data_153 : _GEN_482; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_484 = 8'h9a == _match_key_bytes_21_T_1 ? phv_data_154 : _GEN_483; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_485 = 8'h9b == _match_key_bytes_21_T_1 ? phv_data_155 : _GEN_484; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_486 = 8'h9c == _match_key_bytes_21_T_1 ? phv_data_156 : _GEN_485; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_487 = 8'h9d == _match_key_bytes_21_T_1 ? phv_data_157 : _GEN_486; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_488 = 8'h9e == _match_key_bytes_21_T_1 ? phv_data_158 : _GEN_487; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_489 = 8'h9f == _match_key_bytes_21_T_1 ? phv_data_159 : _GEN_488; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_21 = 8'h2 < _GEN_6 ? _GEN_489 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_20_T_1 = key_offset + 8'h3; // @[matcher.scala 72:98]
  wire [7:0] _GEN_492 = 8'h1 == _match_key_bytes_20_T_1 ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_493 = 8'h2 == _match_key_bytes_20_T_1 ? phv_data_2 : _GEN_492; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_494 = 8'h3 == _match_key_bytes_20_T_1 ? phv_data_3 : _GEN_493; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_495 = 8'h4 == _match_key_bytes_20_T_1 ? phv_data_4 : _GEN_494; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_496 = 8'h5 == _match_key_bytes_20_T_1 ? phv_data_5 : _GEN_495; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_497 = 8'h6 == _match_key_bytes_20_T_1 ? phv_data_6 : _GEN_496; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_498 = 8'h7 == _match_key_bytes_20_T_1 ? phv_data_7 : _GEN_497; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_499 = 8'h8 == _match_key_bytes_20_T_1 ? phv_data_8 : _GEN_498; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_500 = 8'h9 == _match_key_bytes_20_T_1 ? phv_data_9 : _GEN_499; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_501 = 8'ha == _match_key_bytes_20_T_1 ? phv_data_10 : _GEN_500; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_502 = 8'hb == _match_key_bytes_20_T_1 ? phv_data_11 : _GEN_501; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_503 = 8'hc == _match_key_bytes_20_T_1 ? phv_data_12 : _GEN_502; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_504 = 8'hd == _match_key_bytes_20_T_1 ? phv_data_13 : _GEN_503; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_505 = 8'he == _match_key_bytes_20_T_1 ? phv_data_14 : _GEN_504; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_506 = 8'hf == _match_key_bytes_20_T_1 ? phv_data_15 : _GEN_505; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_507 = 8'h10 == _match_key_bytes_20_T_1 ? phv_data_16 : _GEN_506; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_508 = 8'h11 == _match_key_bytes_20_T_1 ? phv_data_17 : _GEN_507; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_509 = 8'h12 == _match_key_bytes_20_T_1 ? phv_data_18 : _GEN_508; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_510 = 8'h13 == _match_key_bytes_20_T_1 ? phv_data_19 : _GEN_509; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_511 = 8'h14 == _match_key_bytes_20_T_1 ? phv_data_20 : _GEN_510; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_512 = 8'h15 == _match_key_bytes_20_T_1 ? phv_data_21 : _GEN_511; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_513 = 8'h16 == _match_key_bytes_20_T_1 ? phv_data_22 : _GEN_512; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_514 = 8'h17 == _match_key_bytes_20_T_1 ? phv_data_23 : _GEN_513; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_515 = 8'h18 == _match_key_bytes_20_T_1 ? phv_data_24 : _GEN_514; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_516 = 8'h19 == _match_key_bytes_20_T_1 ? phv_data_25 : _GEN_515; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_517 = 8'h1a == _match_key_bytes_20_T_1 ? phv_data_26 : _GEN_516; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_518 = 8'h1b == _match_key_bytes_20_T_1 ? phv_data_27 : _GEN_517; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_519 = 8'h1c == _match_key_bytes_20_T_1 ? phv_data_28 : _GEN_518; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_520 = 8'h1d == _match_key_bytes_20_T_1 ? phv_data_29 : _GEN_519; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_521 = 8'h1e == _match_key_bytes_20_T_1 ? phv_data_30 : _GEN_520; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_522 = 8'h1f == _match_key_bytes_20_T_1 ? phv_data_31 : _GEN_521; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_523 = 8'h20 == _match_key_bytes_20_T_1 ? phv_data_32 : _GEN_522; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_524 = 8'h21 == _match_key_bytes_20_T_1 ? phv_data_33 : _GEN_523; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_525 = 8'h22 == _match_key_bytes_20_T_1 ? phv_data_34 : _GEN_524; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_526 = 8'h23 == _match_key_bytes_20_T_1 ? phv_data_35 : _GEN_525; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_527 = 8'h24 == _match_key_bytes_20_T_1 ? phv_data_36 : _GEN_526; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_528 = 8'h25 == _match_key_bytes_20_T_1 ? phv_data_37 : _GEN_527; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_529 = 8'h26 == _match_key_bytes_20_T_1 ? phv_data_38 : _GEN_528; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_530 = 8'h27 == _match_key_bytes_20_T_1 ? phv_data_39 : _GEN_529; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_531 = 8'h28 == _match_key_bytes_20_T_1 ? phv_data_40 : _GEN_530; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_532 = 8'h29 == _match_key_bytes_20_T_1 ? phv_data_41 : _GEN_531; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_533 = 8'h2a == _match_key_bytes_20_T_1 ? phv_data_42 : _GEN_532; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_534 = 8'h2b == _match_key_bytes_20_T_1 ? phv_data_43 : _GEN_533; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_535 = 8'h2c == _match_key_bytes_20_T_1 ? phv_data_44 : _GEN_534; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_536 = 8'h2d == _match_key_bytes_20_T_1 ? phv_data_45 : _GEN_535; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_537 = 8'h2e == _match_key_bytes_20_T_1 ? phv_data_46 : _GEN_536; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_538 = 8'h2f == _match_key_bytes_20_T_1 ? phv_data_47 : _GEN_537; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_539 = 8'h30 == _match_key_bytes_20_T_1 ? phv_data_48 : _GEN_538; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_540 = 8'h31 == _match_key_bytes_20_T_1 ? phv_data_49 : _GEN_539; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_541 = 8'h32 == _match_key_bytes_20_T_1 ? phv_data_50 : _GEN_540; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_542 = 8'h33 == _match_key_bytes_20_T_1 ? phv_data_51 : _GEN_541; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_543 = 8'h34 == _match_key_bytes_20_T_1 ? phv_data_52 : _GEN_542; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_544 = 8'h35 == _match_key_bytes_20_T_1 ? phv_data_53 : _GEN_543; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_545 = 8'h36 == _match_key_bytes_20_T_1 ? phv_data_54 : _GEN_544; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_546 = 8'h37 == _match_key_bytes_20_T_1 ? phv_data_55 : _GEN_545; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_547 = 8'h38 == _match_key_bytes_20_T_1 ? phv_data_56 : _GEN_546; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_548 = 8'h39 == _match_key_bytes_20_T_1 ? phv_data_57 : _GEN_547; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_549 = 8'h3a == _match_key_bytes_20_T_1 ? phv_data_58 : _GEN_548; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_550 = 8'h3b == _match_key_bytes_20_T_1 ? phv_data_59 : _GEN_549; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_551 = 8'h3c == _match_key_bytes_20_T_1 ? phv_data_60 : _GEN_550; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_552 = 8'h3d == _match_key_bytes_20_T_1 ? phv_data_61 : _GEN_551; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_553 = 8'h3e == _match_key_bytes_20_T_1 ? phv_data_62 : _GEN_552; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_554 = 8'h3f == _match_key_bytes_20_T_1 ? phv_data_63 : _GEN_553; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_555 = 8'h40 == _match_key_bytes_20_T_1 ? phv_data_64 : _GEN_554; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_556 = 8'h41 == _match_key_bytes_20_T_1 ? phv_data_65 : _GEN_555; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_557 = 8'h42 == _match_key_bytes_20_T_1 ? phv_data_66 : _GEN_556; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_558 = 8'h43 == _match_key_bytes_20_T_1 ? phv_data_67 : _GEN_557; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_559 = 8'h44 == _match_key_bytes_20_T_1 ? phv_data_68 : _GEN_558; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_560 = 8'h45 == _match_key_bytes_20_T_1 ? phv_data_69 : _GEN_559; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_561 = 8'h46 == _match_key_bytes_20_T_1 ? phv_data_70 : _GEN_560; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_562 = 8'h47 == _match_key_bytes_20_T_1 ? phv_data_71 : _GEN_561; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_563 = 8'h48 == _match_key_bytes_20_T_1 ? phv_data_72 : _GEN_562; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_564 = 8'h49 == _match_key_bytes_20_T_1 ? phv_data_73 : _GEN_563; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_565 = 8'h4a == _match_key_bytes_20_T_1 ? phv_data_74 : _GEN_564; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_566 = 8'h4b == _match_key_bytes_20_T_1 ? phv_data_75 : _GEN_565; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_567 = 8'h4c == _match_key_bytes_20_T_1 ? phv_data_76 : _GEN_566; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_568 = 8'h4d == _match_key_bytes_20_T_1 ? phv_data_77 : _GEN_567; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_569 = 8'h4e == _match_key_bytes_20_T_1 ? phv_data_78 : _GEN_568; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_570 = 8'h4f == _match_key_bytes_20_T_1 ? phv_data_79 : _GEN_569; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_571 = 8'h50 == _match_key_bytes_20_T_1 ? phv_data_80 : _GEN_570; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_572 = 8'h51 == _match_key_bytes_20_T_1 ? phv_data_81 : _GEN_571; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_573 = 8'h52 == _match_key_bytes_20_T_1 ? phv_data_82 : _GEN_572; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_574 = 8'h53 == _match_key_bytes_20_T_1 ? phv_data_83 : _GEN_573; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_575 = 8'h54 == _match_key_bytes_20_T_1 ? phv_data_84 : _GEN_574; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_576 = 8'h55 == _match_key_bytes_20_T_1 ? phv_data_85 : _GEN_575; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_577 = 8'h56 == _match_key_bytes_20_T_1 ? phv_data_86 : _GEN_576; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_578 = 8'h57 == _match_key_bytes_20_T_1 ? phv_data_87 : _GEN_577; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_579 = 8'h58 == _match_key_bytes_20_T_1 ? phv_data_88 : _GEN_578; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_580 = 8'h59 == _match_key_bytes_20_T_1 ? phv_data_89 : _GEN_579; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_581 = 8'h5a == _match_key_bytes_20_T_1 ? phv_data_90 : _GEN_580; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_582 = 8'h5b == _match_key_bytes_20_T_1 ? phv_data_91 : _GEN_581; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_583 = 8'h5c == _match_key_bytes_20_T_1 ? phv_data_92 : _GEN_582; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_584 = 8'h5d == _match_key_bytes_20_T_1 ? phv_data_93 : _GEN_583; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_585 = 8'h5e == _match_key_bytes_20_T_1 ? phv_data_94 : _GEN_584; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_586 = 8'h5f == _match_key_bytes_20_T_1 ? phv_data_95 : _GEN_585; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_587 = 8'h60 == _match_key_bytes_20_T_1 ? phv_data_96 : _GEN_586; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_588 = 8'h61 == _match_key_bytes_20_T_1 ? phv_data_97 : _GEN_587; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_589 = 8'h62 == _match_key_bytes_20_T_1 ? phv_data_98 : _GEN_588; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_590 = 8'h63 == _match_key_bytes_20_T_1 ? phv_data_99 : _GEN_589; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_591 = 8'h64 == _match_key_bytes_20_T_1 ? phv_data_100 : _GEN_590; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_592 = 8'h65 == _match_key_bytes_20_T_1 ? phv_data_101 : _GEN_591; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_593 = 8'h66 == _match_key_bytes_20_T_1 ? phv_data_102 : _GEN_592; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_594 = 8'h67 == _match_key_bytes_20_T_1 ? phv_data_103 : _GEN_593; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_595 = 8'h68 == _match_key_bytes_20_T_1 ? phv_data_104 : _GEN_594; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_596 = 8'h69 == _match_key_bytes_20_T_1 ? phv_data_105 : _GEN_595; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_597 = 8'h6a == _match_key_bytes_20_T_1 ? phv_data_106 : _GEN_596; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_598 = 8'h6b == _match_key_bytes_20_T_1 ? phv_data_107 : _GEN_597; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_599 = 8'h6c == _match_key_bytes_20_T_1 ? phv_data_108 : _GEN_598; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_600 = 8'h6d == _match_key_bytes_20_T_1 ? phv_data_109 : _GEN_599; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_601 = 8'h6e == _match_key_bytes_20_T_1 ? phv_data_110 : _GEN_600; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_602 = 8'h6f == _match_key_bytes_20_T_1 ? phv_data_111 : _GEN_601; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_603 = 8'h70 == _match_key_bytes_20_T_1 ? phv_data_112 : _GEN_602; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_604 = 8'h71 == _match_key_bytes_20_T_1 ? phv_data_113 : _GEN_603; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_605 = 8'h72 == _match_key_bytes_20_T_1 ? phv_data_114 : _GEN_604; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_606 = 8'h73 == _match_key_bytes_20_T_1 ? phv_data_115 : _GEN_605; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_607 = 8'h74 == _match_key_bytes_20_T_1 ? phv_data_116 : _GEN_606; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_608 = 8'h75 == _match_key_bytes_20_T_1 ? phv_data_117 : _GEN_607; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_609 = 8'h76 == _match_key_bytes_20_T_1 ? phv_data_118 : _GEN_608; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_610 = 8'h77 == _match_key_bytes_20_T_1 ? phv_data_119 : _GEN_609; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_611 = 8'h78 == _match_key_bytes_20_T_1 ? phv_data_120 : _GEN_610; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_612 = 8'h79 == _match_key_bytes_20_T_1 ? phv_data_121 : _GEN_611; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_613 = 8'h7a == _match_key_bytes_20_T_1 ? phv_data_122 : _GEN_612; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_614 = 8'h7b == _match_key_bytes_20_T_1 ? phv_data_123 : _GEN_613; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_615 = 8'h7c == _match_key_bytes_20_T_1 ? phv_data_124 : _GEN_614; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_616 = 8'h7d == _match_key_bytes_20_T_1 ? phv_data_125 : _GEN_615; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_617 = 8'h7e == _match_key_bytes_20_T_1 ? phv_data_126 : _GEN_616; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_618 = 8'h7f == _match_key_bytes_20_T_1 ? phv_data_127 : _GEN_617; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_619 = 8'h80 == _match_key_bytes_20_T_1 ? phv_data_128 : _GEN_618; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_620 = 8'h81 == _match_key_bytes_20_T_1 ? phv_data_129 : _GEN_619; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_621 = 8'h82 == _match_key_bytes_20_T_1 ? phv_data_130 : _GEN_620; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_622 = 8'h83 == _match_key_bytes_20_T_1 ? phv_data_131 : _GEN_621; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_623 = 8'h84 == _match_key_bytes_20_T_1 ? phv_data_132 : _GEN_622; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_624 = 8'h85 == _match_key_bytes_20_T_1 ? phv_data_133 : _GEN_623; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_625 = 8'h86 == _match_key_bytes_20_T_1 ? phv_data_134 : _GEN_624; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_626 = 8'h87 == _match_key_bytes_20_T_1 ? phv_data_135 : _GEN_625; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_627 = 8'h88 == _match_key_bytes_20_T_1 ? phv_data_136 : _GEN_626; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_628 = 8'h89 == _match_key_bytes_20_T_1 ? phv_data_137 : _GEN_627; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_629 = 8'h8a == _match_key_bytes_20_T_1 ? phv_data_138 : _GEN_628; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_630 = 8'h8b == _match_key_bytes_20_T_1 ? phv_data_139 : _GEN_629; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_631 = 8'h8c == _match_key_bytes_20_T_1 ? phv_data_140 : _GEN_630; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_632 = 8'h8d == _match_key_bytes_20_T_1 ? phv_data_141 : _GEN_631; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_633 = 8'h8e == _match_key_bytes_20_T_1 ? phv_data_142 : _GEN_632; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_634 = 8'h8f == _match_key_bytes_20_T_1 ? phv_data_143 : _GEN_633; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_635 = 8'h90 == _match_key_bytes_20_T_1 ? phv_data_144 : _GEN_634; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_636 = 8'h91 == _match_key_bytes_20_T_1 ? phv_data_145 : _GEN_635; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_637 = 8'h92 == _match_key_bytes_20_T_1 ? phv_data_146 : _GEN_636; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_638 = 8'h93 == _match_key_bytes_20_T_1 ? phv_data_147 : _GEN_637; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_639 = 8'h94 == _match_key_bytes_20_T_1 ? phv_data_148 : _GEN_638; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_640 = 8'h95 == _match_key_bytes_20_T_1 ? phv_data_149 : _GEN_639; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_641 = 8'h96 == _match_key_bytes_20_T_1 ? phv_data_150 : _GEN_640; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_642 = 8'h97 == _match_key_bytes_20_T_1 ? phv_data_151 : _GEN_641; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_643 = 8'h98 == _match_key_bytes_20_T_1 ? phv_data_152 : _GEN_642; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_644 = 8'h99 == _match_key_bytes_20_T_1 ? phv_data_153 : _GEN_643; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_645 = 8'h9a == _match_key_bytes_20_T_1 ? phv_data_154 : _GEN_644; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_646 = 8'h9b == _match_key_bytes_20_T_1 ? phv_data_155 : _GEN_645; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_647 = 8'h9c == _match_key_bytes_20_T_1 ? phv_data_156 : _GEN_646; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_648 = 8'h9d == _match_key_bytes_20_T_1 ? phv_data_157 : _GEN_647; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_649 = 8'h9e == _match_key_bytes_20_T_1 ? phv_data_158 : _GEN_648; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_650 = 8'h9f == _match_key_bytes_20_T_1 ? phv_data_159 : _GEN_649; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_20 = 8'h3 < _GEN_6 ? _GEN_650 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_19_T_1 = key_offset + 8'h4; // @[matcher.scala 72:98]
  wire [7:0] _GEN_653 = 8'h1 == _match_key_bytes_19_T_1 ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_654 = 8'h2 == _match_key_bytes_19_T_1 ? phv_data_2 : _GEN_653; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_655 = 8'h3 == _match_key_bytes_19_T_1 ? phv_data_3 : _GEN_654; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_656 = 8'h4 == _match_key_bytes_19_T_1 ? phv_data_4 : _GEN_655; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_657 = 8'h5 == _match_key_bytes_19_T_1 ? phv_data_5 : _GEN_656; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_658 = 8'h6 == _match_key_bytes_19_T_1 ? phv_data_6 : _GEN_657; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_659 = 8'h7 == _match_key_bytes_19_T_1 ? phv_data_7 : _GEN_658; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_660 = 8'h8 == _match_key_bytes_19_T_1 ? phv_data_8 : _GEN_659; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_661 = 8'h9 == _match_key_bytes_19_T_1 ? phv_data_9 : _GEN_660; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_662 = 8'ha == _match_key_bytes_19_T_1 ? phv_data_10 : _GEN_661; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_663 = 8'hb == _match_key_bytes_19_T_1 ? phv_data_11 : _GEN_662; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_664 = 8'hc == _match_key_bytes_19_T_1 ? phv_data_12 : _GEN_663; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_665 = 8'hd == _match_key_bytes_19_T_1 ? phv_data_13 : _GEN_664; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_666 = 8'he == _match_key_bytes_19_T_1 ? phv_data_14 : _GEN_665; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_667 = 8'hf == _match_key_bytes_19_T_1 ? phv_data_15 : _GEN_666; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_668 = 8'h10 == _match_key_bytes_19_T_1 ? phv_data_16 : _GEN_667; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_669 = 8'h11 == _match_key_bytes_19_T_1 ? phv_data_17 : _GEN_668; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_670 = 8'h12 == _match_key_bytes_19_T_1 ? phv_data_18 : _GEN_669; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_671 = 8'h13 == _match_key_bytes_19_T_1 ? phv_data_19 : _GEN_670; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_672 = 8'h14 == _match_key_bytes_19_T_1 ? phv_data_20 : _GEN_671; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_673 = 8'h15 == _match_key_bytes_19_T_1 ? phv_data_21 : _GEN_672; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_674 = 8'h16 == _match_key_bytes_19_T_1 ? phv_data_22 : _GEN_673; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_675 = 8'h17 == _match_key_bytes_19_T_1 ? phv_data_23 : _GEN_674; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_676 = 8'h18 == _match_key_bytes_19_T_1 ? phv_data_24 : _GEN_675; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_677 = 8'h19 == _match_key_bytes_19_T_1 ? phv_data_25 : _GEN_676; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_678 = 8'h1a == _match_key_bytes_19_T_1 ? phv_data_26 : _GEN_677; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_679 = 8'h1b == _match_key_bytes_19_T_1 ? phv_data_27 : _GEN_678; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_680 = 8'h1c == _match_key_bytes_19_T_1 ? phv_data_28 : _GEN_679; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_681 = 8'h1d == _match_key_bytes_19_T_1 ? phv_data_29 : _GEN_680; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_682 = 8'h1e == _match_key_bytes_19_T_1 ? phv_data_30 : _GEN_681; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_683 = 8'h1f == _match_key_bytes_19_T_1 ? phv_data_31 : _GEN_682; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_684 = 8'h20 == _match_key_bytes_19_T_1 ? phv_data_32 : _GEN_683; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_685 = 8'h21 == _match_key_bytes_19_T_1 ? phv_data_33 : _GEN_684; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_686 = 8'h22 == _match_key_bytes_19_T_1 ? phv_data_34 : _GEN_685; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_687 = 8'h23 == _match_key_bytes_19_T_1 ? phv_data_35 : _GEN_686; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_688 = 8'h24 == _match_key_bytes_19_T_1 ? phv_data_36 : _GEN_687; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_689 = 8'h25 == _match_key_bytes_19_T_1 ? phv_data_37 : _GEN_688; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_690 = 8'h26 == _match_key_bytes_19_T_1 ? phv_data_38 : _GEN_689; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_691 = 8'h27 == _match_key_bytes_19_T_1 ? phv_data_39 : _GEN_690; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_692 = 8'h28 == _match_key_bytes_19_T_1 ? phv_data_40 : _GEN_691; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_693 = 8'h29 == _match_key_bytes_19_T_1 ? phv_data_41 : _GEN_692; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_694 = 8'h2a == _match_key_bytes_19_T_1 ? phv_data_42 : _GEN_693; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_695 = 8'h2b == _match_key_bytes_19_T_1 ? phv_data_43 : _GEN_694; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_696 = 8'h2c == _match_key_bytes_19_T_1 ? phv_data_44 : _GEN_695; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_697 = 8'h2d == _match_key_bytes_19_T_1 ? phv_data_45 : _GEN_696; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_698 = 8'h2e == _match_key_bytes_19_T_1 ? phv_data_46 : _GEN_697; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_699 = 8'h2f == _match_key_bytes_19_T_1 ? phv_data_47 : _GEN_698; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_700 = 8'h30 == _match_key_bytes_19_T_1 ? phv_data_48 : _GEN_699; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_701 = 8'h31 == _match_key_bytes_19_T_1 ? phv_data_49 : _GEN_700; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_702 = 8'h32 == _match_key_bytes_19_T_1 ? phv_data_50 : _GEN_701; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_703 = 8'h33 == _match_key_bytes_19_T_1 ? phv_data_51 : _GEN_702; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_704 = 8'h34 == _match_key_bytes_19_T_1 ? phv_data_52 : _GEN_703; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_705 = 8'h35 == _match_key_bytes_19_T_1 ? phv_data_53 : _GEN_704; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_706 = 8'h36 == _match_key_bytes_19_T_1 ? phv_data_54 : _GEN_705; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_707 = 8'h37 == _match_key_bytes_19_T_1 ? phv_data_55 : _GEN_706; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_708 = 8'h38 == _match_key_bytes_19_T_1 ? phv_data_56 : _GEN_707; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_709 = 8'h39 == _match_key_bytes_19_T_1 ? phv_data_57 : _GEN_708; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_710 = 8'h3a == _match_key_bytes_19_T_1 ? phv_data_58 : _GEN_709; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_711 = 8'h3b == _match_key_bytes_19_T_1 ? phv_data_59 : _GEN_710; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_712 = 8'h3c == _match_key_bytes_19_T_1 ? phv_data_60 : _GEN_711; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_713 = 8'h3d == _match_key_bytes_19_T_1 ? phv_data_61 : _GEN_712; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_714 = 8'h3e == _match_key_bytes_19_T_1 ? phv_data_62 : _GEN_713; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_715 = 8'h3f == _match_key_bytes_19_T_1 ? phv_data_63 : _GEN_714; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_716 = 8'h40 == _match_key_bytes_19_T_1 ? phv_data_64 : _GEN_715; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_717 = 8'h41 == _match_key_bytes_19_T_1 ? phv_data_65 : _GEN_716; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_718 = 8'h42 == _match_key_bytes_19_T_1 ? phv_data_66 : _GEN_717; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_719 = 8'h43 == _match_key_bytes_19_T_1 ? phv_data_67 : _GEN_718; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_720 = 8'h44 == _match_key_bytes_19_T_1 ? phv_data_68 : _GEN_719; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_721 = 8'h45 == _match_key_bytes_19_T_1 ? phv_data_69 : _GEN_720; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_722 = 8'h46 == _match_key_bytes_19_T_1 ? phv_data_70 : _GEN_721; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_723 = 8'h47 == _match_key_bytes_19_T_1 ? phv_data_71 : _GEN_722; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_724 = 8'h48 == _match_key_bytes_19_T_1 ? phv_data_72 : _GEN_723; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_725 = 8'h49 == _match_key_bytes_19_T_1 ? phv_data_73 : _GEN_724; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_726 = 8'h4a == _match_key_bytes_19_T_1 ? phv_data_74 : _GEN_725; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_727 = 8'h4b == _match_key_bytes_19_T_1 ? phv_data_75 : _GEN_726; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_728 = 8'h4c == _match_key_bytes_19_T_1 ? phv_data_76 : _GEN_727; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_729 = 8'h4d == _match_key_bytes_19_T_1 ? phv_data_77 : _GEN_728; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_730 = 8'h4e == _match_key_bytes_19_T_1 ? phv_data_78 : _GEN_729; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_731 = 8'h4f == _match_key_bytes_19_T_1 ? phv_data_79 : _GEN_730; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_732 = 8'h50 == _match_key_bytes_19_T_1 ? phv_data_80 : _GEN_731; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_733 = 8'h51 == _match_key_bytes_19_T_1 ? phv_data_81 : _GEN_732; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_734 = 8'h52 == _match_key_bytes_19_T_1 ? phv_data_82 : _GEN_733; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_735 = 8'h53 == _match_key_bytes_19_T_1 ? phv_data_83 : _GEN_734; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_736 = 8'h54 == _match_key_bytes_19_T_1 ? phv_data_84 : _GEN_735; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_737 = 8'h55 == _match_key_bytes_19_T_1 ? phv_data_85 : _GEN_736; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_738 = 8'h56 == _match_key_bytes_19_T_1 ? phv_data_86 : _GEN_737; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_739 = 8'h57 == _match_key_bytes_19_T_1 ? phv_data_87 : _GEN_738; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_740 = 8'h58 == _match_key_bytes_19_T_1 ? phv_data_88 : _GEN_739; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_741 = 8'h59 == _match_key_bytes_19_T_1 ? phv_data_89 : _GEN_740; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_742 = 8'h5a == _match_key_bytes_19_T_1 ? phv_data_90 : _GEN_741; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_743 = 8'h5b == _match_key_bytes_19_T_1 ? phv_data_91 : _GEN_742; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_744 = 8'h5c == _match_key_bytes_19_T_1 ? phv_data_92 : _GEN_743; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_745 = 8'h5d == _match_key_bytes_19_T_1 ? phv_data_93 : _GEN_744; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_746 = 8'h5e == _match_key_bytes_19_T_1 ? phv_data_94 : _GEN_745; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_747 = 8'h5f == _match_key_bytes_19_T_1 ? phv_data_95 : _GEN_746; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_748 = 8'h60 == _match_key_bytes_19_T_1 ? phv_data_96 : _GEN_747; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_749 = 8'h61 == _match_key_bytes_19_T_1 ? phv_data_97 : _GEN_748; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_750 = 8'h62 == _match_key_bytes_19_T_1 ? phv_data_98 : _GEN_749; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_751 = 8'h63 == _match_key_bytes_19_T_1 ? phv_data_99 : _GEN_750; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_752 = 8'h64 == _match_key_bytes_19_T_1 ? phv_data_100 : _GEN_751; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_753 = 8'h65 == _match_key_bytes_19_T_1 ? phv_data_101 : _GEN_752; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_754 = 8'h66 == _match_key_bytes_19_T_1 ? phv_data_102 : _GEN_753; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_755 = 8'h67 == _match_key_bytes_19_T_1 ? phv_data_103 : _GEN_754; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_756 = 8'h68 == _match_key_bytes_19_T_1 ? phv_data_104 : _GEN_755; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_757 = 8'h69 == _match_key_bytes_19_T_1 ? phv_data_105 : _GEN_756; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_758 = 8'h6a == _match_key_bytes_19_T_1 ? phv_data_106 : _GEN_757; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_759 = 8'h6b == _match_key_bytes_19_T_1 ? phv_data_107 : _GEN_758; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_760 = 8'h6c == _match_key_bytes_19_T_1 ? phv_data_108 : _GEN_759; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_761 = 8'h6d == _match_key_bytes_19_T_1 ? phv_data_109 : _GEN_760; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_762 = 8'h6e == _match_key_bytes_19_T_1 ? phv_data_110 : _GEN_761; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_763 = 8'h6f == _match_key_bytes_19_T_1 ? phv_data_111 : _GEN_762; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_764 = 8'h70 == _match_key_bytes_19_T_1 ? phv_data_112 : _GEN_763; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_765 = 8'h71 == _match_key_bytes_19_T_1 ? phv_data_113 : _GEN_764; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_766 = 8'h72 == _match_key_bytes_19_T_1 ? phv_data_114 : _GEN_765; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_767 = 8'h73 == _match_key_bytes_19_T_1 ? phv_data_115 : _GEN_766; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_768 = 8'h74 == _match_key_bytes_19_T_1 ? phv_data_116 : _GEN_767; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_769 = 8'h75 == _match_key_bytes_19_T_1 ? phv_data_117 : _GEN_768; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_770 = 8'h76 == _match_key_bytes_19_T_1 ? phv_data_118 : _GEN_769; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_771 = 8'h77 == _match_key_bytes_19_T_1 ? phv_data_119 : _GEN_770; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_772 = 8'h78 == _match_key_bytes_19_T_1 ? phv_data_120 : _GEN_771; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_773 = 8'h79 == _match_key_bytes_19_T_1 ? phv_data_121 : _GEN_772; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_774 = 8'h7a == _match_key_bytes_19_T_1 ? phv_data_122 : _GEN_773; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_775 = 8'h7b == _match_key_bytes_19_T_1 ? phv_data_123 : _GEN_774; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_776 = 8'h7c == _match_key_bytes_19_T_1 ? phv_data_124 : _GEN_775; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_777 = 8'h7d == _match_key_bytes_19_T_1 ? phv_data_125 : _GEN_776; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_778 = 8'h7e == _match_key_bytes_19_T_1 ? phv_data_126 : _GEN_777; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_779 = 8'h7f == _match_key_bytes_19_T_1 ? phv_data_127 : _GEN_778; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_780 = 8'h80 == _match_key_bytes_19_T_1 ? phv_data_128 : _GEN_779; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_781 = 8'h81 == _match_key_bytes_19_T_1 ? phv_data_129 : _GEN_780; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_782 = 8'h82 == _match_key_bytes_19_T_1 ? phv_data_130 : _GEN_781; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_783 = 8'h83 == _match_key_bytes_19_T_1 ? phv_data_131 : _GEN_782; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_784 = 8'h84 == _match_key_bytes_19_T_1 ? phv_data_132 : _GEN_783; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_785 = 8'h85 == _match_key_bytes_19_T_1 ? phv_data_133 : _GEN_784; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_786 = 8'h86 == _match_key_bytes_19_T_1 ? phv_data_134 : _GEN_785; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_787 = 8'h87 == _match_key_bytes_19_T_1 ? phv_data_135 : _GEN_786; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_788 = 8'h88 == _match_key_bytes_19_T_1 ? phv_data_136 : _GEN_787; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_789 = 8'h89 == _match_key_bytes_19_T_1 ? phv_data_137 : _GEN_788; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_790 = 8'h8a == _match_key_bytes_19_T_1 ? phv_data_138 : _GEN_789; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_791 = 8'h8b == _match_key_bytes_19_T_1 ? phv_data_139 : _GEN_790; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_792 = 8'h8c == _match_key_bytes_19_T_1 ? phv_data_140 : _GEN_791; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_793 = 8'h8d == _match_key_bytes_19_T_1 ? phv_data_141 : _GEN_792; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_794 = 8'h8e == _match_key_bytes_19_T_1 ? phv_data_142 : _GEN_793; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_795 = 8'h8f == _match_key_bytes_19_T_1 ? phv_data_143 : _GEN_794; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_796 = 8'h90 == _match_key_bytes_19_T_1 ? phv_data_144 : _GEN_795; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_797 = 8'h91 == _match_key_bytes_19_T_1 ? phv_data_145 : _GEN_796; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_798 = 8'h92 == _match_key_bytes_19_T_1 ? phv_data_146 : _GEN_797; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_799 = 8'h93 == _match_key_bytes_19_T_1 ? phv_data_147 : _GEN_798; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_800 = 8'h94 == _match_key_bytes_19_T_1 ? phv_data_148 : _GEN_799; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_801 = 8'h95 == _match_key_bytes_19_T_1 ? phv_data_149 : _GEN_800; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_802 = 8'h96 == _match_key_bytes_19_T_1 ? phv_data_150 : _GEN_801; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_803 = 8'h97 == _match_key_bytes_19_T_1 ? phv_data_151 : _GEN_802; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_804 = 8'h98 == _match_key_bytes_19_T_1 ? phv_data_152 : _GEN_803; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_805 = 8'h99 == _match_key_bytes_19_T_1 ? phv_data_153 : _GEN_804; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_806 = 8'h9a == _match_key_bytes_19_T_1 ? phv_data_154 : _GEN_805; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_807 = 8'h9b == _match_key_bytes_19_T_1 ? phv_data_155 : _GEN_806; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_808 = 8'h9c == _match_key_bytes_19_T_1 ? phv_data_156 : _GEN_807; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_809 = 8'h9d == _match_key_bytes_19_T_1 ? phv_data_157 : _GEN_808; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_810 = 8'h9e == _match_key_bytes_19_T_1 ? phv_data_158 : _GEN_809; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_811 = 8'h9f == _match_key_bytes_19_T_1 ? phv_data_159 : _GEN_810; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_19 = 8'h4 < _GEN_6 ? _GEN_811 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_18_T_1 = key_offset + 8'h5; // @[matcher.scala 72:98]
  wire [7:0] _GEN_814 = 8'h1 == _match_key_bytes_18_T_1 ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_815 = 8'h2 == _match_key_bytes_18_T_1 ? phv_data_2 : _GEN_814; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_816 = 8'h3 == _match_key_bytes_18_T_1 ? phv_data_3 : _GEN_815; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_817 = 8'h4 == _match_key_bytes_18_T_1 ? phv_data_4 : _GEN_816; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_818 = 8'h5 == _match_key_bytes_18_T_1 ? phv_data_5 : _GEN_817; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_819 = 8'h6 == _match_key_bytes_18_T_1 ? phv_data_6 : _GEN_818; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_820 = 8'h7 == _match_key_bytes_18_T_1 ? phv_data_7 : _GEN_819; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_821 = 8'h8 == _match_key_bytes_18_T_1 ? phv_data_8 : _GEN_820; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_822 = 8'h9 == _match_key_bytes_18_T_1 ? phv_data_9 : _GEN_821; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_823 = 8'ha == _match_key_bytes_18_T_1 ? phv_data_10 : _GEN_822; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_824 = 8'hb == _match_key_bytes_18_T_1 ? phv_data_11 : _GEN_823; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_825 = 8'hc == _match_key_bytes_18_T_1 ? phv_data_12 : _GEN_824; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_826 = 8'hd == _match_key_bytes_18_T_1 ? phv_data_13 : _GEN_825; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_827 = 8'he == _match_key_bytes_18_T_1 ? phv_data_14 : _GEN_826; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_828 = 8'hf == _match_key_bytes_18_T_1 ? phv_data_15 : _GEN_827; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_829 = 8'h10 == _match_key_bytes_18_T_1 ? phv_data_16 : _GEN_828; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_830 = 8'h11 == _match_key_bytes_18_T_1 ? phv_data_17 : _GEN_829; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_831 = 8'h12 == _match_key_bytes_18_T_1 ? phv_data_18 : _GEN_830; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_832 = 8'h13 == _match_key_bytes_18_T_1 ? phv_data_19 : _GEN_831; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_833 = 8'h14 == _match_key_bytes_18_T_1 ? phv_data_20 : _GEN_832; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_834 = 8'h15 == _match_key_bytes_18_T_1 ? phv_data_21 : _GEN_833; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_835 = 8'h16 == _match_key_bytes_18_T_1 ? phv_data_22 : _GEN_834; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_836 = 8'h17 == _match_key_bytes_18_T_1 ? phv_data_23 : _GEN_835; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_837 = 8'h18 == _match_key_bytes_18_T_1 ? phv_data_24 : _GEN_836; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_838 = 8'h19 == _match_key_bytes_18_T_1 ? phv_data_25 : _GEN_837; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_839 = 8'h1a == _match_key_bytes_18_T_1 ? phv_data_26 : _GEN_838; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_840 = 8'h1b == _match_key_bytes_18_T_1 ? phv_data_27 : _GEN_839; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_841 = 8'h1c == _match_key_bytes_18_T_1 ? phv_data_28 : _GEN_840; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_842 = 8'h1d == _match_key_bytes_18_T_1 ? phv_data_29 : _GEN_841; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_843 = 8'h1e == _match_key_bytes_18_T_1 ? phv_data_30 : _GEN_842; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_844 = 8'h1f == _match_key_bytes_18_T_1 ? phv_data_31 : _GEN_843; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_845 = 8'h20 == _match_key_bytes_18_T_1 ? phv_data_32 : _GEN_844; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_846 = 8'h21 == _match_key_bytes_18_T_1 ? phv_data_33 : _GEN_845; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_847 = 8'h22 == _match_key_bytes_18_T_1 ? phv_data_34 : _GEN_846; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_848 = 8'h23 == _match_key_bytes_18_T_1 ? phv_data_35 : _GEN_847; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_849 = 8'h24 == _match_key_bytes_18_T_1 ? phv_data_36 : _GEN_848; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_850 = 8'h25 == _match_key_bytes_18_T_1 ? phv_data_37 : _GEN_849; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_851 = 8'h26 == _match_key_bytes_18_T_1 ? phv_data_38 : _GEN_850; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_852 = 8'h27 == _match_key_bytes_18_T_1 ? phv_data_39 : _GEN_851; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_853 = 8'h28 == _match_key_bytes_18_T_1 ? phv_data_40 : _GEN_852; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_854 = 8'h29 == _match_key_bytes_18_T_1 ? phv_data_41 : _GEN_853; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_855 = 8'h2a == _match_key_bytes_18_T_1 ? phv_data_42 : _GEN_854; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_856 = 8'h2b == _match_key_bytes_18_T_1 ? phv_data_43 : _GEN_855; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_857 = 8'h2c == _match_key_bytes_18_T_1 ? phv_data_44 : _GEN_856; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_858 = 8'h2d == _match_key_bytes_18_T_1 ? phv_data_45 : _GEN_857; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_859 = 8'h2e == _match_key_bytes_18_T_1 ? phv_data_46 : _GEN_858; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_860 = 8'h2f == _match_key_bytes_18_T_1 ? phv_data_47 : _GEN_859; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_861 = 8'h30 == _match_key_bytes_18_T_1 ? phv_data_48 : _GEN_860; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_862 = 8'h31 == _match_key_bytes_18_T_1 ? phv_data_49 : _GEN_861; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_863 = 8'h32 == _match_key_bytes_18_T_1 ? phv_data_50 : _GEN_862; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_864 = 8'h33 == _match_key_bytes_18_T_1 ? phv_data_51 : _GEN_863; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_865 = 8'h34 == _match_key_bytes_18_T_1 ? phv_data_52 : _GEN_864; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_866 = 8'h35 == _match_key_bytes_18_T_1 ? phv_data_53 : _GEN_865; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_867 = 8'h36 == _match_key_bytes_18_T_1 ? phv_data_54 : _GEN_866; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_868 = 8'h37 == _match_key_bytes_18_T_1 ? phv_data_55 : _GEN_867; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_869 = 8'h38 == _match_key_bytes_18_T_1 ? phv_data_56 : _GEN_868; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_870 = 8'h39 == _match_key_bytes_18_T_1 ? phv_data_57 : _GEN_869; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_871 = 8'h3a == _match_key_bytes_18_T_1 ? phv_data_58 : _GEN_870; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_872 = 8'h3b == _match_key_bytes_18_T_1 ? phv_data_59 : _GEN_871; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_873 = 8'h3c == _match_key_bytes_18_T_1 ? phv_data_60 : _GEN_872; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_874 = 8'h3d == _match_key_bytes_18_T_1 ? phv_data_61 : _GEN_873; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_875 = 8'h3e == _match_key_bytes_18_T_1 ? phv_data_62 : _GEN_874; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_876 = 8'h3f == _match_key_bytes_18_T_1 ? phv_data_63 : _GEN_875; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_877 = 8'h40 == _match_key_bytes_18_T_1 ? phv_data_64 : _GEN_876; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_878 = 8'h41 == _match_key_bytes_18_T_1 ? phv_data_65 : _GEN_877; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_879 = 8'h42 == _match_key_bytes_18_T_1 ? phv_data_66 : _GEN_878; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_880 = 8'h43 == _match_key_bytes_18_T_1 ? phv_data_67 : _GEN_879; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_881 = 8'h44 == _match_key_bytes_18_T_1 ? phv_data_68 : _GEN_880; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_882 = 8'h45 == _match_key_bytes_18_T_1 ? phv_data_69 : _GEN_881; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_883 = 8'h46 == _match_key_bytes_18_T_1 ? phv_data_70 : _GEN_882; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_884 = 8'h47 == _match_key_bytes_18_T_1 ? phv_data_71 : _GEN_883; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_885 = 8'h48 == _match_key_bytes_18_T_1 ? phv_data_72 : _GEN_884; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_886 = 8'h49 == _match_key_bytes_18_T_1 ? phv_data_73 : _GEN_885; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_887 = 8'h4a == _match_key_bytes_18_T_1 ? phv_data_74 : _GEN_886; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_888 = 8'h4b == _match_key_bytes_18_T_1 ? phv_data_75 : _GEN_887; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_889 = 8'h4c == _match_key_bytes_18_T_1 ? phv_data_76 : _GEN_888; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_890 = 8'h4d == _match_key_bytes_18_T_1 ? phv_data_77 : _GEN_889; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_891 = 8'h4e == _match_key_bytes_18_T_1 ? phv_data_78 : _GEN_890; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_892 = 8'h4f == _match_key_bytes_18_T_1 ? phv_data_79 : _GEN_891; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_893 = 8'h50 == _match_key_bytes_18_T_1 ? phv_data_80 : _GEN_892; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_894 = 8'h51 == _match_key_bytes_18_T_1 ? phv_data_81 : _GEN_893; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_895 = 8'h52 == _match_key_bytes_18_T_1 ? phv_data_82 : _GEN_894; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_896 = 8'h53 == _match_key_bytes_18_T_1 ? phv_data_83 : _GEN_895; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_897 = 8'h54 == _match_key_bytes_18_T_1 ? phv_data_84 : _GEN_896; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_898 = 8'h55 == _match_key_bytes_18_T_1 ? phv_data_85 : _GEN_897; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_899 = 8'h56 == _match_key_bytes_18_T_1 ? phv_data_86 : _GEN_898; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_900 = 8'h57 == _match_key_bytes_18_T_1 ? phv_data_87 : _GEN_899; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_901 = 8'h58 == _match_key_bytes_18_T_1 ? phv_data_88 : _GEN_900; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_902 = 8'h59 == _match_key_bytes_18_T_1 ? phv_data_89 : _GEN_901; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_903 = 8'h5a == _match_key_bytes_18_T_1 ? phv_data_90 : _GEN_902; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_904 = 8'h5b == _match_key_bytes_18_T_1 ? phv_data_91 : _GEN_903; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_905 = 8'h5c == _match_key_bytes_18_T_1 ? phv_data_92 : _GEN_904; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_906 = 8'h5d == _match_key_bytes_18_T_1 ? phv_data_93 : _GEN_905; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_907 = 8'h5e == _match_key_bytes_18_T_1 ? phv_data_94 : _GEN_906; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_908 = 8'h5f == _match_key_bytes_18_T_1 ? phv_data_95 : _GEN_907; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_909 = 8'h60 == _match_key_bytes_18_T_1 ? phv_data_96 : _GEN_908; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_910 = 8'h61 == _match_key_bytes_18_T_1 ? phv_data_97 : _GEN_909; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_911 = 8'h62 == _match_key_bytes_18_T_1 ? phv_data_98 : _GEN_910; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_912 = 8'h63 == _match_key_bytes_18_T_1 ? phv_data_99 : _GEN_911; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_913 = 8'h64 == _match_key_bytes_18_T_1 ? phv_data_100 : _GEN_912; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_914 = 8'h65 == _match_key_bytes_18_T_1 ? phv_data_101 : _GEN_913; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_915 = 8'h66 == _match_key_bytes_18_T_1 ? phv_data_102 : _GEN_914; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_916 = 8'h67 == _match_key_bytes_18_T_1 ? phv_data_103 : _GEN_915; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_917 = 8'h68 == _match_key_bytes_18_T_1 ? phv_data_104 : _GEN_916; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_918 = 8'h69 == _match_key_bytes_18_T_1 ? phv_data_105 : _GEN_917; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_919 = 8'h6a == _match_key_bytes_18_T_1 ? phv_data_106 : _GEN_918; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_920 = 8'h6b == _match_key_bytes_18_T_1 ? phv_data_107 : _GEN_919; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_921 = 8'h6c == _match_key_bytes_18_T_1 ? phv_data_108 : _GEN_920; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_922 = 8'h6d == _match_key_bytes_18_T_1 ? phv_data_109 : _GEN_921; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_923 = 8'h6e == _match_key_bytes_18_T_1 ? phv_data_110 : _GEN_922; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_924 = 8'h6f == _match_key_bytes_18_T_1 ? phv_data_111 : _GEN_923; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_925 = 8'h70 == _match_key_bytes_18_T_1 ? phv_data_112 : _GEN_924; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_926 = 8'h71 == _match_key_bytes_18_T_1 ? phv_data_113 : _GEN_925; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_927 = 8'h72 == _match_key_bytes_18_T_1 ? phv_data_114 : _GEN_926; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_928 = 8'h73 == _match_key_bytes_18_T_1 ? phv_data_115 : _GEN_927; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_929 = 8'h74 == _match_key_bytes_18_T_1 ? phv_data_116 : _GEN_928; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_930 = 8'h75 == _match_key_bytes_18_T_1 ? phv_data_117 : _GEN_929; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_931 = 8'h76 == _match_key_bytes_18_T_1 ? phv_data_118 : _GEN_930; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_932 = 8'h77 == _match_key_bytes_18_T_1 ? phv_data_119 : _GEN_931; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_933 = 8'h78 == _match_key_bytes_18_T_1 ? phv_data_120 : _GEN_932; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_934 = 8'h79 == _match_key_bytes_18_T_1 ? phv_data_121 : _GEN_933; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_935 = 8'h7a == _match_key_bytes_18_T_1 ? phv_data_122 : _GEN_934; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_936 = 8'h7b == _match_key_bytes_18_T_1 ? phv_data_123 : _GEN_935; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_937 = 8'h7c == _match_key_bytes_18_T_1 ? phv_data_124 : _GEN_936; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_938 = 8'h7d == _match_key_bytes_18_T_1 ? phv_data_125 : _GEN_937; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_939 = 8'h7e == _match_key_bytes_18_T_1 ? phv_data_126 : _GEN_938; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_940 = 8'h7f == _match_key_bytes_18_T_1 ? phv_data_127 : _GEN_939; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_941 = 8'h80 == _match_key_bytes_18_T_1 ? phv_data_128 : _GEN_940; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_942 = 8'h81 == _match_key_bytes_18_T_1 ? phv_data_129 : _GEN_941; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_943 = 8'h82 == _match_key_bytes_18_T_1 ? phv_data_130 : _GEN_942; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_944 = 8'h83 == _match_key_bytes_18_T_1 ? phv_data_131 : _GEN_943; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_945 = 8'h84 == _match_key_bytes_18_T_1 ? phv_data_132 : _GEN_944; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_946 = 8'h85 == _match_key_bytes_18_T_1 ? phv_data_133 : _GEN_945; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_947 = 8'h86 == _match_key_bytes_18_T_1 ? phv_data_134 : _GEN_946; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_948 = 8'h87 == _match_key_bytes_18_T_1 ? phv_data_135 : _GEN_947; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_949 = 8'h88 == _match_key_bytes_18_T_1 ? phv_data_136 : _GEN_948; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_950 = 8'h89 == _match_key_bytes_18_T_1 ? phv_data_137 : _GEN_949; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_951 = 8'h8a == _match_key_bytes_18_T_1 ? phv_data_138 : _GEN_950; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_952 = 8'h8b == _match_key_bytes_18_T_1 ? phv_data_139 : _GEN_951; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_953 = 8'h8c == _match_key_bytes_18_T_1 ? phv_data_140 : _GEN_952; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_954 = 8'h8d == _match_key_bytes_18_T_1 ? phv_data_141 : _GEN_953; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_955 = 8'h8e == _match_key_bytes_18_T_1 ? phv_data_142 : _GEN_954; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_956 = 8'h8f == _match_key_bytes_18_T_1 ? phv_data_143 : _GEN_955; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_957 = 8'h90 == _match_key_bytes_18_T_1 ? phv_data_144 : _GEN_956; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_958 = 8'h91 == _match_key_bytes_18_T_1 ? phv_data_145 : _GEN_957; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_959 = 8'h92 == _match_key_bytes_18_T_1 ? phv_data_146 : _GEN_958; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_960 = 8'h93 == _match_key_bytes_18_T_1 ? phv_data_147 : _GEN_959; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_961 = 8'h94 == _match_key_bytes_18_T_1 ? phv_data_148 : _GEN_960; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_962 = 8'h95 == _match_key_bytes_18_T_1 ? phv_data_149 : _GEN_961; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_963 = 8'h96 == _match_key_bytes_18_T_1 ? phv_data_150 : _GEN_962; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_964 = 8'h97 == _match_key_bytes_18_T_1 ? phv_data_151 : _GEN_963; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_965 = 8'h98 == _match_key_bytes_18_T_1 ? phv_data_152 : _GEN_964; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_966 = 8'h99 == _match_key_bytes_18_T_1 ? phv_data_153 : _GEN_965; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_967 = 8'h9a == _match_key_bytes_18_T_1 ? phv_data_154 : _GEN_966; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_968 = 8'h9b == _match_key_bytes_18_T_1 ? phv_data_155 : _GEN_967; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_969 = 8'h9c == _match_key_bytes_18_T_1 ? phv_data_156 : _GEN_968; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_970 = 8'h9d == _match_key_bytes_18_T_1 ? phv_data_157 : _GEN_969; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_971 = 8'h9e == _match_key_bytes_18_T_1 ? phv_data_158 : _GEN_970; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_972 = 8'h9f == _match_key_bytes_18_T_1 ? phv_data_159 : _GEN_971; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_18 = 8'h5 < _GEN_6 ? _GEN_972 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_17_T_1 = key_offset + 8'h6; // @[matcher.scala 72:98]
  wire [7:0] _GEN_975 = 8'h1 == _match_key_bytes_17_T_1 ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_976 = 8'h2 == _match_key_bytes_17_T_1 ? phv_data_2 : _GEN_975; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_977 = 8'h3 == _match_key_bytes_17_T_1 ? phv_data_3 : _GEN_976; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_978 = 8'h4 == _match_key_bytes_17_T_1 ? phv_data_4 : _GEN_977; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_979 = 8'h5 == _match_key_bytes_17_T_1 ? phv_data_5 : _GEN_978; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_980 = 8'h6 == _match_key_bytes_17_T_1 ? phv_data_6 : _GEN_979; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_981 = 8'h7 == _match_key_bytes_17_T_1 ? phv_data_7 : _GEN_980; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_982 = 8'h8 == _match_key_bytes_17_T_1 ? phv_data_8 : _GEN_981; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_983 = 8'h9 == _match_key_bytes_17_T_1 ? phv_data_9 : _GEN_982; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_984 = 8'ha == _match_key_bytes_17_T_1 ? phv_data_10 : _GEN_983; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_985 = 8'hb == _match_key_bytes_17_T_1 ? phv_data_11 : _GEN_984; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_986 = 8'hc == _match_key_bytes_17_T_1 ? phv_data_12 : _GEN_985; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_987 = 8'hd == _match_key_bytes_17_T_1 ? phv_data_13 : _GEN_986; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_988 = 8'he == _match_key_bytes_17_T_1 ? phv_data_14 : _GEN_987; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_989 = 8'hf == _match_key_bytes_17_T_1 ? phv_data_15 : _GEN_988; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_990 = 8'h10 == _match_key_bytes_17_T_1 ? phv_data_16 : _GEN_989; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_991 = 8'h11 == _match_key_bytes_17_T_1 ? phv_data_17 : _GEN_990; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_992 = 8'h12 == _match_key_bytes_17_T_1 ? phv_data_18 : _GEN_991; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_993 = 8'h13 == _match_key_bytes_17_T_1 ? phv_data_19 : _GEN_992; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_994 = 8'h14 == _match_key_bytes_17_T_1 ? phv_data_20 : _GEN_993; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_995 = 8'h15 == _match_key_bytes_17_T_1 ? phv_data_21 : _GEN_994; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_996 = 8'h16 == _match_key_bytes_17_T_1 ? phv_data_22 : _GEN_995; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_997 = 8'h17 == _match_key_bytes_17_T_1 ? phv_data_23 : _GEN_996; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_998 = 8'h18 == _match_key_bytes_17_T_1 ? phv_data_24 : _GEN_997; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_999 = 8'h19 == _match_key_bytes_17_T_1 ? phv_data_25 : _GEN_998; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1000 = 8'h1a == _match_key_bytes_17_T_1 ? phv_data_26 : _GEN_999; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1001 = 8'h1b == _match_key_bytes_17_T_1 ? phv_data_27 : _GEN_1000; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1002 = 8'h1c == _match_key_bytes_17_T_1 ? phv_data_28 : _GEN_1001; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1003 = 8'h1d == _match_key_bytes_17_T_1 ? phv_data_29 : _GEN_1002; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1004 = 8'h1e == _match_key_bytes_17_T_1 ? phv_data_30 : _GEN_1003; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1005 = 8'h1f == _match_key_bytes_17_T_1 ? phv_data_31 : _GEN_1004; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1006 = 8'h20 == _match_key_bytes_17_T_1 ? phv_data_32 : _GEN_1005; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1007 = 8'h21 == _match_key_bytes_17_T_1 ? phv_data_33 : _GEN_1006; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1008 = 8'h22 == _match_key_bytes_17_T_1 ? phv_data_34 : _GEN_1007; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1009 = 8'h23 == _match_key_bytes_17_T_1 ? phv_data_35 : _GEN_1008; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1010 = 8'h24 == _match_key_bytes_17_T_1 ? phv_data_36 : _GEN_1009; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1011 = 8'h25 == _match_key_bytes_17_T_1 ? phv_data_37 : _GEN_1010; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1012 = 8'h26 == _match_key_bytes_17_T_1 ? phv_data_38 : _GEN_1011; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1013 = 8'h27 == _match_key_bytes_17_T_1 ? phv_data_39 : _GEN_1012; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1014 = 8'h28 == _match_key_bytes_17_T_1 ? phv_data_40 : _GEN_1013; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1015 = 8'h29 == _match_key_bytes_17_T_1 ? phv_data_41 : _GEN_1014; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1016 = 8'h2a == _match_key_bytes_17_T_1 ? phv_data_42 : _GEN_1015; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1017 = 8'h2b == _match_key_bytes_17_T_1 ? phv_data_43 : _GEN_1016; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1018 = 8'h2c == _match_key_bytes_17_T_1 ? phv_data_44 : _GEN_1017; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1019 = 8'h2d == _match_key_bytes_17_T_1 ? phv_data_45 : _GEN_1018; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1020 = 8'h2e == _match_key_bytes_17_T_1 ? phv_data_46 : _GEN_1019; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1021 = 8'h2f == _match_key_bytes_17_T_1 ? phv_data_47 : _GEN_1020; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1022 = 8'h30 == _match_key_bytes_17_T_1 ? phv_data_48 : _GEN_1021; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1023 = 8'h31 == _match_key_bytes_17_T_1 ? phv_data_49 : _GEN_1022; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1024 = 8'h32 == _match_key_bytes_17_T_1 ? phv_data_50 : _GEN_1023; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1025 = 8'h33 == _match_key_bytes_17_T_1 ? phv_data_51 : _GEN_1024; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1026 = 8'h34 == _match_key_bytes_17_T_1 ? phv_data_52 : _GEN_1025; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1027 = 8'h35 == _match_key_bytes_17_T_1 ? phv_data_53 : _GEN_1026; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1028 = 8'h36 == _match_key_bytes_17_T_1 ? phv_data_54 : _GEN_1027; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1029 = 8'h37 == _match_key_bytes_17_T_1 ? phv_data_55 : _GEN_1028; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1030 = 8'h38 == _match_key_bytes_17_T_1 ? phv_data_56 : _GEN_1029; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1031 = 8'h39 == _match_key_bytes_17_T_1 ? phv_data_57 : _GEN_1030; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1032 = 8'h3a == _match_key_bytes_17_T_1 ? phv_data_58 : _GEN_1031; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1033 = 8'h3b == _match_key_bytes_17_T_1 ? phv_data_59 : _GEN_1032; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1034 = 8'h3c == _match_key_bytes_17_T_1 ? phv_data_60 : _GEN_1033; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1035 = 8'h3d == _match_key_bytes_17_T_1 ? phv_data_61 : _GEN_1034; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1036 = 8'h3e == _match_key_bytes_17_T_1 ? phv_data_62 : _GEN_1035; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1037 = 8'h3f == _match_key_bytes_17_T_1 ? phv_data_63 : _GEN_1036; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1038 = 8'h40 == _match_key_bytes_17_T_1 ? phv_data_64 : _GEN_1037; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1039 = 8'h41 == _match_key_bytes_17_T_1 ? phv_data_65 : _GEN_1038; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1040 = 8'h42 == _match_key_bytes_17_T_1 ? phv_data_66 : _GEN_1039; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1041 = 8'h43 == _match_key_bytes_17_T_1 ? phv_data_67 : _GEN_1040; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1042 = 8'h44 == _match_key_bytes_17_T_1 ? phv_data_68 : _GEN_1041; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1043 = 8'h45 == _match_key_bytes_17_T_1 ? phv_data_69 : _GEN_1042; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1044 = 8'h46 == _match_key_bytes_17_T_1 ? phv_data_70 : _GEN_1043; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1045 = 8'h47 == _match_key_bytes_17_T_1 ? phv_data_71 : _GEN_1044; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1046 = 8'h48 == _match_key_bytes_17_T_1 ? phv_data_72 : _GEN_1045; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1047 = 8'h49 == _match_key_bytes_17_T_1 ? phv_data_73 : _GEN_1046; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1048 = 8'h4a == _match_key_bytes_17_T_1 ? phv_data_74 : _GEN_1047; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1049 = 8'h4b == _match_key_bytes_17_T_1 ? phv_data_75 : _GEN_1048; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1050 = 8'h4c == _match_key_bytes_17_T_1 ? phv_data_76 : _GEN_1049; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1051 = 8'h4d == _match_key_bytes_17_T_1 ? phv_data_77 : _GEN_1050; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1052 = 8'h4e == _match_key_bytes_17_T_1 ? phv_data_78 : _GEN_1051; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1053 = 8'h4f == _match_key_bytes_17_T_1 ? phv_data_79 : _GEN_1052; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1054 = 8'h50 == _match_key_bytes_17_T_1 ? phv_data_80 : _GEN_1053; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1055 = 8'h51 == _match_key_bytes_17_T_1 ? phv_data_81 : _GEN_1054; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1056 = 8'h52 == _match_key_bytes_17_T_1 ? phv_data_82 : _GEN_1055; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1057 = 8'h53 == _match_key_bytes_17_T_1 ? phv_data_83 : _GEN_1056; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1058 = 8'h54 == _match_key_bytes_17_T_1 ? phv_data_84 : _GEN_1057; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1059 = 8'h55 == _match_key_bytes_17_T_1 ? phv_data_85 : _GEN_1058; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1060 = 8'h56 == _match_key_bytes_17_T_1 ? phv_data_86 : _GEN_1059; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1061 = 8'h57 == _match_key_bytes_17_T_1 ? phv_data_87 : _GEN_1060; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1062 = 8'h58 == _match_key_bytes_17_T_1 ? phv_data_88 : _GEN_1061; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1063 = 8'h59 == _match_key_bytes_17_T_1 ? phv_data_89 : _GEN_1062; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1064 = 8'h5a == _match_key_bytes_17_T_1 ? phv_data_90 : _GEN_1063; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1065 = 8'h5b == _match_key_bytes_17_T_1 ? phv_data_91 : _GEN_1064; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1066 = 8'h5c == _match_key_bytes_17_T_1 ? phv_data_92 : _GEN_1065; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1067 = 8'h5d == _match_key_bytes_17_T_1 ? phv_data_93 : _GEN_1066; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1068 = 8'h5e == _match_key_bytes_17_T_1 ? phv_data_94 : _GEN_1067; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1069 = 8'h5f == _match_key_bytes_17_T_1 ? phv_data_95 : _GEN_1068; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1070 = 8'h60 == _match_key_bytes_17_T_1 ? phv_data_96 : _GEN_1069; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1071 = 8'h61 == _match_key_bytes_17_T_1 ? phv_data_97 : _GEN_1070; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1072 = 8'h62 == _match_key_bytes_17_T_1 ? phv_data_98 : _GEN_1071; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1073 = 8'h63 == _match_key_bytes_17_T_1 ? phv_data_99 : _GEN_1072; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1074 = 8'h64 == _match_key_bytes_17_T_1 ? phv_data_100 : _GEN_1073; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1075 = 8'h65 == _match_key_bytes_17_T_1 ? phv_data_101 : _GEN_1074; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1076 = 8'h66 == _match_key_bytes_17_T_1 ? phv_data_102 : _GEN_1075; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1077 = 8'h67 == _match_key_bytes_17_T_1 ? phv_data_103 : _GEN_1076; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1078 = 8'h68 == _match_key_bytes_17_T_1 ? phv_data_104 : _GEN_1077; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1079 = 8'h69 == _match_key_bytes_17_T_1 ? phv_data_105 : _GEN_1078; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1080 = 8'h6a == _match_key_bytes_17_T_1 ? phv_data_106 : _GEN_1079; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1081 = 8'h6b == _match_key_bytes_17_T_1 ? phv_data_107 : _GEN_1080; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1082 = 8'h6c == _match_key_bytes_17_T_1 ? phv_data_108 : _GEN_1081; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1083 = 8'h6d == _match_key_bytes_17_T_1 ? phv_data_109 : _GEN_1082; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1084 = 8'h6e == _match_key_bytes_17_T_1 ? phv_data_110 : _GEN_1083; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1085 = 8'h6f == _match_key_bytes_17_T_1 ? phv_data_111 : _GEN_1084; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1086 = 8'h70 == _match_key_bytes_17_T_1 ? phv_data_112 : _GEN_1085; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1087 = 8'h71 == _match_key_bytes_17_T_1 ? phv_data_113 : _GEN_1086; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1088 = 8'h72 == _match_key_bytes_17_T_1 ? phv_data_114 : _GEN_1087; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1089 = 8'h73 == _match_key_bytes_17_T_1 ? phv_data_115 : _GEN_1088; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1090 = 8'h74 == _match_key_bytes_17_T_1 ? phv_data_116 : _GEN_1089; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1091 = 8'h75 == _match_key_bytes_17_T_1 ? phv_data_117 : _GEN_1090; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1092 = 8'h76 == _match_key_bytes_17_T_1 ? phv_data_118 : _GEN_1091; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1093 = 8'h77 == _match_key_bytes_17_T_1 ? phv_data_119 : _GEN_1092; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1094 = 8'h78 == _match_key_bytes_17_T_1 ? phv_data_120 : _GEN_1093; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1095 = 8'h79 == _match_key_bytes_17_T_1 ? phv_data_121 : _GEN_1094; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1096 = 8'h7a == _match_key_bytes_17_T_1 ? phv_data_122 : _GEN_1095; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1097 = 8'h7b == _match_key_bytes_17_T_1 ? phv_data_123 : _GEN_1096; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1098 = 8'h7c == _match_key_bytes_17_T_1 ? phv_data_124 : _GEN_1097; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1099 = 8'h7d == _match_key_bytes_17_T_1 ? phv_data_125 : _GEN_1098; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1100 = 8'h7e == _match_key_bytes_17_T_1 ? phv_data_126 : _GEN_1099; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1101 = 8'h7f == _match_key_bytes_17_T_1 ? phv_data_127 : _GEN_1100; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1102 = 8'h80 == _match_key_bytes_17_T_1 ? phv_data_128 : _GEN_1101; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1103 = 8'h81 == _match_key_bytes_17_T_1 ? phv_data_129 : _GEN_1102; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1104 = 8'h82 == _match_key_bytes_17_T_1 ? phv_data_130 : _GEN_1103; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1105 = 8'h83 == _match_key_bytes_17_T_1 ? phv_data_131 : _GEN_1104; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1106 = 8'h84 == _match_key_bytes_17_T_1 ? phv_data_132 : _GEN_1105; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1107 = 8'h85 == _match_key_bytes_17_T_1 ? phv_data_133 : _GEN_1106; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1108 = 8'h86 == _match_key_bytes_17_T_1 ? phv_data_134 : _GEN_1107; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1109 = 8'h87 == _match_key_bytes_17_T_1 ? phv_data_135 : _GEN_1108; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1110 = 8'h88 == _match_key_bytes_17_T_1 ? phv_data_136 : _GEN_1109; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1111 = 8'h89 == _match_key_bytes_17_T_1 ? phv_data_137 : _GEN_1110; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1112 = 8'h8a == _match_key_bytes_17_T_1 ? phv_data_138 : _GEN_1111; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1113 = 8'h8b == _match_key_bytes_17_T_1 ? phv_data_139 : _GEN_1112; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1114 = 8'h8c == _match_key_bytes_17_T_1 ? phv_data_140 : _GEN_1113; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1115 = 8'h8d == _match_key_bytes_17_T_1 ? phv_data_141 : _GEN_1114; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1116 = 8'h8e == _match_key_bytes_17_T_1 ? phv_data_142 : _GEN_1115; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1117 = 8'h8f == _match_key_bytes_17_T_1 ? phv_data_143 : _GEN_1116; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1118 = 8'h90 == _match_key_bytes_17_T_1 ? phv_data_144 : _GEN_1117; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1119 = 8'h91 == _match_key_bytes_17_T_1 ? phv_data_145 : _GEN_1118; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1120 = 8'h92 == _match_key_bytes_17_T_1 ? phv_data_146 : _GEN_1119; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1121 = 8'h93 == _match_key_bytes_17_T_1 ? phv_data_147 : _GEN_1120; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1122 = 8'h94 == _match_key_bytes_17_T_1 ? phv_data_148 : _GEN_1121; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1123 = 8'h95 == _match_key_bytes_17_T_1 ? phv_data_149 : _GEN_1122; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1124 = 8'h96 == _match_key_bytes_17_T_1 ? phv_data_150 : _GEN_1123; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1125 = 8'h97 == _match_key_bytes_17_T_1 ? phv_data_151 : _GEN_1124; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1126 = 8'h98 == _match_key_bytes_17_T_1 ? phv_data_152 : _GEN_1125; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1127 = 8'h99 == _match_key_bytes_17_T_1 ? phv_data_153 : _GEN_1126; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1128 = 8'h9a == _match_key_bytes_17_T_1 ? phv_data_154 : _GEN_1127; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1129 = 8'h9b == _match_key_bytes_17_T_1 ? phv_data_155 : _GEN_1128; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1130 = 8'h9c == _match_key_bytes_17_T_1 ? phv_data_156 : _GEN_1129; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1131 = 8'h9d == _match_key_bytes_17_T_1 ? phv_data_157 : _GEN_1130; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1132 = 8'h9e == _match_key_bytes_17_T_1 ? phv_data_158 : _GEN_1131; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1133 = 8'h9f == _match_key_bytes_17_T_1 ? phv_data_159 : _GEN_1132; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_17 = 8'h6 < _GEN_6 ? _GEN_1133 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_16_T_1 = key_offset + 8'h7; // @[matcher.scala 72:98]
  wire [7:0] _GEN_1136 = 8'h1 == _match_key_bytes_16_T_1 ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1137 = 8'h2 == _match_key_bytes_16_T_1 ? phv_data_2 : _GEN_1136; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1138 = 8'h3 == _match_key_bytes_16_T_1 ? phv_data_3 : _GEN_1137; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1139 = 8'h4 == _match_key_bytes_16_T_1 ? phv_data_4 : _GEN_1138; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1140 = 8'h5 == _match_key_bytes_16_T_1 ? phv_data_5 : _GEN_1139; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1141 = 8'h6 == _match_key_bytes_16_T_1 ? phv_data_6 : _GEN_1140; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1142 = 8'h7 == _match_key_bytes_16_T_1 ? phv_data_7 : _GEN_1141; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1143 = 8'h8 == _match_key_bytes_16_T_1 ? phv_data_8 : _GEN_1142; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1144 = 8'h9 == _match_key_bytes_16_T_1 ? phv_data_9 : _GEN_1143; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1145 = 8'ha == _match_key_bytes_16_T_1 ? phv_data_10 : _GEN_1144; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1146 = 8'hb == _match_key_bytes_16_T_1 ? phv_data_11 : _GEN_1145; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1147 = 8'hc == _match_key_bytes_16_T_1 ? phv_data_12 : _GEN_1146; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1148 = 8'hd == _match_key_bytes_16_T_1 ? phv_data_13 : _GEN_1147; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1149 = 8'he == _match_key_bytes_16_T_1 ? phv_data_14 : _GEN_1148; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1150 = 8'hf == _match_key_bytes_16_T_1 ? phv_data_15 : _GEN_1149; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1151 = 8'h10 == _match_key_bytes_16_T_1 ? phv_data_16 : _GEN_1150; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1152 = 8'h11 == _match_key_bytes_16_T_1 ? phv_data_17 : _GEN_1151; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1153 = 8'h12 == _match_key_bytes_16_T_1 ? phv_data_18 : _GEN_1152; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1154 = 8'h13 == _match_key_bytes_16_T_1 ? phv_data_19 : _GEN_1153; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1155 = 8'h14 == _match_key_bytes_16_T_1 ? phv_data_20 : _GEN_1154; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1156 = 8'h15 == _match_key_bytes_16_T_1 ? phv_data_21 : _GEN_1155; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1157 = 8'h16 == _match_key_bytes_16_T_1 ? phv_data_22 : _GEN_1156; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1158 = 8'h17 == _match_key_bytes_16_T_1 ? phv_data_23 : _GEN_1157; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1159 = 8'h18 == _match_key_bytes_16_T_1 ? phv_data_24 : _GEN_1158; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1160 = 8'h19 == _match_key_bytes_16_T_1 ? phv_data_25 : _GEN_1159; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1161 = 8'h1a == _match_key_bytes_16_T_1 ? phv_data_26 : _GEN_1160; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1162 = 8'h1b == _match_key_bytes_16_T_1 ? phv_data_27 : _GEN_1161; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1163 = 8'h1c == _match_key_bytes_16_T_1 ? phv_data_28 : _GEN_1162; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1164 = 8'h1d == _match_key_bytes_16_T_1 ? phv_data_29 : _GEN_1163; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1165 = 8'h1e == _match_key_bytes_16_T_1 ? phv_data_30 : _GEN_1164; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1166 = 8'h1f == _match_key_bytes_16_T_1 ? phv_data_31 : _GEN_1165; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1167 = 8'h20 == _match_key_bytes_16_T_1 ? phv_data_32 : _GEN_1166; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1168 = 8'h21 == _match_key_bytes_16_T_1 ? phv_data_33 : _GEN_1167; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1169 = 8'h22 == _match_key_bytes_16_T_1 ? phv_data_34 : _GEN_1168; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1170 = 8'h23 == _match_key_bytes_16_T_1 ? phv_data_35 : _GEN_1169; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1171 = 8'h24 == _match_key_bytes_16_T_1 ? phv_data_36 : _GEN_1170; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1172 = 8'h25 == _match_key_bytes_16_T_1 ? phv_data_37 : _GEN_1171; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1173 = 8'h26 == _match_key_bytes_16_T_1 ? phv_data_38 : _GEN_1172; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1174 = 8'h27 == _match_key_bytes_16_T_1 ? phv_data_39 : _GEN_1173; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1175 = 8'h28 == _match_key_bytes_16_T_1 ? phv_data_40 : _GEN_1174; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1176 = 8'h29 == _match_key_bytes_16_T_1 ? phv_data_41 : _GEN_1175; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1177 = 8'h2a == _match_key_bytes_16_T_1 ? phv_data_42 : _GEN_1176; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1178 = 8'h2b == _match_key_bytes_16_T_1 ? phv_data_43 : _GEN_1177; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1179 = 8'h2c == _match_key_bytes_16_T_1 ? phv_data_44 : _GEN_1178; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1180 = 8'h2d == _match_key_bytes_16_T_1 ? phv_data_45 : _GEN_1179; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1181 = 8'h2e == _match_key_bytes_16_T_1 ? phv_data_46 : _GEN_1180; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1182 = 8'h2f == _match_key_bytes_16_T_1 ? phv_data_47 : _GEN_1181; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1183 = 8'h30 == _match_key_bytes_16_T_1 ? phv_data_48 : _GEN_1182; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1184 = 8'h31 == _match_key_bytes_16_T_1 ? phv_data_49 : _GEN_1183; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1185 = 8'h32 == _match_key_bytes_16_T_1 ? phv_data_50 : _GEN_1184; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1186 = 8'h33 == _match_key_bytes_16_T_1 ? phv_data_51 : _GEN_1185; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1187 = 8'h34 == _match_key_bytes_16_T_1 ? phv_data_52 : _GEN_1186; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1188 = 8'h35 == _match_key_bytes_16_T_1 ? phv_data_53 : _GEN_1187; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1189 = 8'h36 == _match_key_bytes_16_T_1 ? phv_data_54 : _GEN_1188; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1190 = 8'h37 == _match_key_bytes_16_T_1 ? phv_data_55 : _GEN_1189; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1191 = 8'h38 == _match_key_bytes_16_T_1 ? phv_data_56 : _GEN_1190; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1192 = 8'h39 == _match_key_bytes_16_T_1 ? phv_data_57 : _GEN_1191; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1193 = 8'h3a == _match_key_bytes_16_T_1 ? phv_data_58 : _GEN_1192; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1194 = 8'h3b == _match_key_bytes_16_T_1 ? phv_data_59 : _GEN_1193; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1195 = 8'h3c == _match_key_bytes_16_T_1 ? phv_data_60 : _GEN_1194; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1196 = 8'h3d == _match_key_bytes_16_T_1 ? phv_data_61 : _GEN_1195; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1197 = 8'h3e == _match_key_bytes_16_T_1 ? phv_data_62 : _GEN_1196; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1198 = 8'h3f == _match_key_bytes_16_T_1 ? phv_data_63 : _GEN_1197; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1199 = 8'h40 == _match_key_bytes_16_T_1 ? phv_data_64 : _GEN_1198; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1200 = 8'h41 == _match_key_bytes_16_T_1 ? phv_data_65 : _GEN_1199; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1201 = 8'h42 == _match_key_bytes_16_T_1 ? phv_data_66 : _GEN_1200; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1202 = 8'h43 == _match_key_bytes_16_T_1 ? phv_data_67 : _GEN_1201; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1203 = 8'h44 == _match_key_bytes_16_T_1 ? phv_data_68 : _GEN_1202; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1204 = 8'h45 == _match_key_bytes_16_T_1 ? phv_data_69 : _GEN_1203; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1205 = 8'h46 == _match_key_bytes_16_T_1 ? phv_data_70 : _GEN_1204; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1206 = 8'h47 == _match_key_bytes_16_T_1 ? phv_data_71 : _GEN_1205; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1207 = 8'h48 == _match_key_bytes_16_T_1 ? phv_data_72 : _GEN_1206; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1208 = 8'h49 == _match_key_bytes_16_T_1 ? phv_data_73 : _GEN_1207; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1209 = 8'h4a == _match_key_bytes_16_T_1 ? phv_data_74 : _GEN_1208; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1210 = 8'h4b == _match_key_bytes_16_T_1 ? phv_data_75 : _GEN_1209; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1211 = 8'h4c == _match_key_bytes_16_T_1 ? phv_data_76 : _GEN_1210; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1212 = 8'h4d == _match_key_bytes_16_T_1 ? phv_data_77 : _GEN_1211; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1213 = 8'h4e == _match_key_bytes_16_T_1 ? phv_data_78 : _GEN_1212; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1214 = 8'h4f == _match_key_bytes_16_T_1 ? phv_data_79 : _GEN_1213; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1215 = 8'h50 == _match_key_bytes_16_T_1 ? phv_data_80 : _GEN_1214; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1216 = 8'h51 == _match_key_bytes_16_T_1 ? phv_data_81 : _GEN_1215; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1217 = 8'h52 == _match_key_bytes_16_T_1 ? phv_data_82 : _GEN_1216; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1218 = 8'h53 == _match_key_bytes_16_T_1 ? phv_data_83 : _GEN_1217; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1219 = 8'h54 == _match_key_bytes_16_T_1 ? phv_data_84 : _GEN_1218; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1220 = 8'h55 == _match_key_bytes_16_T_1 ? phv_data_85 : _GEN_1219; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1221 = 8'h56 == _match_key_bytes_16_T_1 ? phv_data_86 : _GEN_1220; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1222 = 8'h57 == _match_key_bytes_16_T_1 ? phv_data_87 : _GEN_1221; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1223 = 8'h58 == _match_key_bytes_16_T_1 ? phv_data_88 : _GEN_1222; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1224 = 8'h59 == _match_key_bytes_16_T_1 ? phv_data_89 : _GEN_1223; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1225 = 8'h5a == _match_key_bytes_16_T_1 ? phv_data_90 : _GEN_1224; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1226 = 8'h5b == _match_key_bytes_16_T_1 ? phv_data_91 : _GEN_1225; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1227 = 8'h5c == _match_key_bytes_16_T_1 ? phv_data_92 : _GEN_1226; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1228 = 8'h5d == _match_key_bytes_16_T_1 ? phv_data_93 : _GEN_1227; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1229 = 8'h5e == _match_key_bytes_16_T_1 ? phv_data_94 : _GEN_1228; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1230 = 8'h5f == _match_key_bytes_16_T_1 ? phv_data_95 : _GEN_1229; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1231 = 8'h60 == _match_key_bytes_16_T_1 ? phv_data_96 : _GEN_1230; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1232 = 8'h61 == _match_key_bytes_16_T_1 ? phv_data_97 : _GEN_1231; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1233 = 8'h62 == _match_key_bytes_16_T_1 ? phv_data_98 : _GEN_1232; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1234 = 8'h63 == _match_key_bytes_16_T_1 ? phv_data_99 : _GEN_1233; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1235 = 8'h64 == _match_key_bytes_16_T_1 ? phv_data_100 : _GEN_1234; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1236 = 8'h65 == _match_key_bytes_16_T_1 ? phv_data_101 : _GEN_1235; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1237 = 8'h66 == _match_key_bytes_16_T_1 ? phv_data_102 : _GEN_1236; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1238 = 8'h67 == _match_key_bytes_16_T_1 ? phv_data_103 : _GEN_1237; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1239 = 8'h68 == _match_key_bytes_16_T_1 ? phv_data_104 : _GEN_1238; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1240 = 8'h69 == _match_key_bytes_16_T_1 ? phv_data_105 : _GEN_1239; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1241 = 8'h6a == _match_key_bytes_16_T_1 ? phv_data_106 : _GEN_1240; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1242 = 8'h6b == _match_key_bytes_16_T_1 ? phv_data_107 : _GEN_1241; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1243 = 8'h6c == _match_key_bytes_16_T_1 ? phv_data_108 : _GEN_1242; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1244 = 8'h6d == _match_key_bytes_16_T_1 ? phv_data_109 : _GEN_1243; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1245 = 8'h6e == _match_key_bytes_16_T_1 ? phv_data_110 : _GEN_1244; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1246 = 8'h6f == _match_key_bytes_16_T_1 ? phv_data_111 : _GEN_1245; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1247 = 8'h70 == _match_key_bytes_16_T_1 ? phv_data_112 : _GEN_1246; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1248 = 8'h71 == _match_key_bytes_16_T_1 ? phv_data_113 : _GEN_1247; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1249 = 8'h72 == _match_key_bytes_16_T_1 ? phv_data_114 : _GEN_1248; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1250 = 8'h73 == _match_key_bytes_16_T_1 ? phv_data_115 : _GEN_1249; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1251 = 8'h74 == _match_key_bytes_16_T_1 ? phv_data_116 : _GEN_1250; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1252 = 8'h75 == _match_key_bytes_16_T_1 ? phv_data_117 : _GEN_1251; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1253 = 8'h76 == _match_key_bytes_16_T_1 ? phv_data_118 : _GEN_1252; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1254 = 8'h77 == _match_key_bytes_16_T_1 ? phv_data_119 : _GEN_1253; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1255 = 8'h78 == _match_key_bytes_16_T_1 ? phv_data_120 : _GEN_1254; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1256 = 8'h79 == _match_key_bytes_16_T_1 ? phv_data_121 : _GEN_1255; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1257 = 8'h7a == _match_key_bytes_16_T_1 ? phv_data_122 : _GEN_1256; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1258 = 8'h7b == _match_key_bytes_16_T_1 ? phv_data_123 : _GEN_1257; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1259 = 8'h7c == _match_key_bytes_16_T_1 ? phv_data_124 : _GEN_1258; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1260 = 8'h7d == _match_key_bytes_16_T_1 ? phv_data_125 : _GEN_1259; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1261 = 8'h7e == _match_key_bytes_16_T_1 ? phv_data_126 : _GEN_1260; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1262 = 8'h7f == _match_key_bytes_16_T_1 ? phv_data_127 : _GEN_1261; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1263 = 8'h80 == _match_key_bytes_16_T_1 ? phv_data_128 : _GEN_1262; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1264 = 8'h81 == _match_key_bytes_16_T_1 ? phv_data_129 : _GEN_1263; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1265 = 8'h82 == _match_key_bytes_16_T_1 ? phv_data_130 : _GEN_1264; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1266 = 8'h83 == _match_key_bytes_16_T_1 ? phv_data_131 : _GEN_1265; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1267 = 8'h84 == _match_key_bytes_16_T_1 ? phv_data_132 : _GEN_1266; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1268 = 8'h85 == _match_key_bytes_16_T_1 ? phv_data_133 : _GEN_1267; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1269 = 8'h86 == _match_key_bytes_16_T_1 ? phv_data_134 : _GEN_1268; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1270 = 8'h87 == _match_key_bytes_16_T_1 ? phv_data_135 : _GEN_1269; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1271 = 8'h88 == _match_key_bytes_16_T_1 ? phv_data_136 : _GEN_1270; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1272 = 8'h89 == _match_key_bytes_16_T_1 ? phv_data_137 : _GEN_1271; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1273 = 8'h8a == _match_key_bytes_16_T_1 ? phv_data_138 : _GEN_1272; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1274 = 8'h8b == _match_key_bytes_16_T_1 ? phv_data_139 : _GEN_1273; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1275 = 8'h8c == _match_key_bytes_16_T_1 ? phv_data_140 : _GEN_1274; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1276 = 8'h8d == _match_key_bytes_16_T_1 ? phv_data_141 : _GEN_1275; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1277 = 8'h8e == _match_key_bytes_16_T_1 ? phv_data_142 : _GEN_1276; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1278 = 8'h8f == _match_key_bytes_16_T_1 ? phv_data_143 : _GEN_1277; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1279 = 8'h90 == _match_key_bytes_16_T_1 ? phv_data_144 : _GEN_1278; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1280 = 8'h91 == _match_key_bytes_16_T_1 ? phv_data_145 : _GEN_1279; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1281 = 8'h92 == _match_key_bytes_16_T_1 ? phv_data_146 : _GEN_1280; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1282 = 8'h93 == _match_key_bytes_16_T_1 ? phv_data_147 : _GEN_1281; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1283 = 8'h94 == _match_key_bytes_16_T_1 ? phv_data_148 : _GEN_1282; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1284 = 8'h95 == _match_key_bytes_16_T_1 ? phv_data_149 : _GEN_1283; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1285 = 8'h96 == _match_key_bytes_16_T_1 ? phv_data_150 : _GEN_1284; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1286 = 8'h97 == _match_key_bytes_16_T_1 ? phv_data_151 : _GEN_1285; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1287 = 8'h98 == _match_key_bytes_16_T_1 ? phv_data_152 : _GEN_1286; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1288 = 8'h99 == _match_key_bytes_16_T_1 ? phv_data_153 : _GEN_1287; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1289 = 8'h9a == _match_key_bytes_16_T_1 ? phv_data_154 : _GEN_1288; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1290 = 8'h9b == _match_key_bytes_16_T_1 ? phv_data_155 : _GEN_1289; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1291 = 8'h9c == _match_key_bytes_16_T_1 ? phv_data_156 : _GEN_1290; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1292 = 8'h9d == _match_key_bytes_16_T_1 ? phv_data_157 : _GEN_1291; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1293 = 8'h9e == _match_key_bytes_16_T_1 ? phv_data_158 : _GEN_1292; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1294 = 8'h9f == _match_key_bytes_16_T_1 ? phv_data_159 : _GEN_1293; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_16 = 8'h7 < _GEN_6 ? _GEN_1294 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_15_T_1 = key_offset + 8'h8; // @[matcher.scala 72:98]
  wire [7:0] _GEN_1297 = 8'h1 == _match_key_bytes_15_T_1 ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1298 = 8'h2 == _match_key_bytes_15_T_1 ? phv_data_2 : _GEN_1297; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1299 = 8'h3 == _match_key_bytes_15_T_1 ? phv_data_3 : _GEN_1298; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1300 = 8'h4 == _match_key_bytes_15_T_1 ? phv_data_4 : _GEN_1299; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1301 = 8'h5 == _match_key_bytes_15_T_1 ? phv_data_5 : _GEN_1300; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1302 = 8'h6 == _match_key_bytes_15_T_1 ? phv_data_6 : _GEN_1301; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1303 = 8'h7 == _match_key_bytes_15_T_1 ? phv_data_7 : _GEN_1302; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1304 = 8'h8 == _match_key_bytes_15_T_1 ? phv_data_8 : _GEN_1303; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1305 = 8'h9 == _match_key_bytes_15_T_1 ? phv_data_9 : _GEN_1304; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1306 = 8'ha == _match_key_bytes_15_T_1 ? phv_data_10 : _GEN_1305; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1307 = 8'hb == _match_key_bytes_15_T_1 ? phv_data_11 : _GEN_1306; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1308 = 8'hc == _match_key_bytes_15_T_1 ? phv_data_12 : _GEN_1307; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1309 = 8'hd == _match_key_bytes_15_T_1 ? phv_data_13 : _GEN_1308; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1310 = 8'he == _match_key_bytes_15_T_1 ? phv_data_14 : _GEN_1309; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1311 = 8'hf == _match_key_bytes_15_T_1 ? phv_data_15 : _GEN_1310; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1312 = 8'h10 == _match_key_bytes_15_T_1 ? phv_data_16 : _GEN_1311; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1313 = 8'h11 == _match_key_bytes_15_T_1 ? phv_data_17 : _GEN_1312; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1314 = 8'h12 == _match_key_bytes_15_T_1 ? phv_data_18 : _GEN_1313; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1315 = 8'h13 == _match_key_bytes_15_T_1 ? phv_data_19 : _GEN_1314; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1316 = 8'h14 == _match_key_bytes_15_T_1 ? phv_data_20 : _GEN_1315; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1317 = 8'h15 == _match_key_bytes_15_T_1 ? phv_data_21 : _GEN_1316; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1318 = 8'h16 == _match_key_bytes_15_T_1 ? phv_data_22 : _GEN_1317; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1319 = 8'h17 == _match_key_bytes_15_T_1 ? phv_data_23 : _GEN_1318; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1320 = 8'h18 == _match_key_bytes_15_T_1 ? phv_data_24 : _GEN_1319; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1321 = 8'h19 == _match_key_bytes_15_T_1 ? phv_data_25 : _GEN_1320; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1322 = 8'h1a == _match_key_bytes_15_T_1 ? phv_data_26 : _GEN_1321; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1323 = 8'h1b == _match_key_bytes_15_T_1 ? phv_data_27 : _GEN_1322; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1324 = 8'h1c == _match_key_bytes_15_T_1 ? phv_data_28 : _GEN_1323; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1325 = 8'h1d == _match_key_bytes_15_T_1 ? phv_data_29 : _GEN_1324; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1326 = 8'h1e == _match_key_bytes_15_T_1 ? phv_data_30 : _GEN_1325; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1327 = 8'h1f == _match_key_bytes_15_T_1 ? phv_data_31 : _GEN_1326; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1328 = 8'h20 == _match_key_bytes_15_T_1 ? phv_data_32 : _GEN_1327; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1329 = 8'h21 == _match_key_bytes_15_T_1 ? phv_data_33 : _GEN_1328; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1330 = 8'h22 == _match_key_bytes_15_T_1 ? phv_data_34 : _GEN_1329; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1331 = 8'h23 == _match_key_bytes_15_T_1 ? phv_data_35 : _GEN_1330; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1332 = 8'h24 == _match_key_bytes_15_T_1 ? phv_data_36 : _GEN_1331; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1333 = 8'h25 == _match_key_bytes_15_T_1 ? phv_data_37 : _GEN_1332; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1334 = 8'h26 == _match_key_bytes_15_T_1 ? phv_data_38 : _GEN_1333; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1335 = 8'h27 == _match_key_bytes_15_T_1 ? phv_data_39 : _GEN_1334; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1336 = 8'h28 == _match_key_bytes_15_T_1 ? phv_data_40 : _GEN_1335; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1337 = 8'h29 == _match_key_bytes_15_T_1 ? phv_data_41 : _GEN_1336; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1338 = 8'h2a == _match_key_bytes_15_T_1 ? phv_data_42 : _GEN_1337; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1339 = 8'h2b == _match_key_bytes_15_T_1 ? phv_data_43 : _GEN_1338; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1340 = 8'h2c == _match_key_bytes_15_T_1 ? phv_data_44 : _GEN_1339; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1341 = 8'h2d == _match_key_bytes_15_T_1 ? phv_data_45 : _GEN_1340; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1342 = 8'h2e == _match_key_bytes_15_T_1 ? phv_data_46 : _GEN_1341; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1343 = 8'h2f == _match_key_bytes_15_T_1 ? phv_data_47 : _GEN_1342; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1344 = 8'h30 == _match_key_bytes_15_T_1 ? phv_data_48 : _GEN_1343; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1345 = 8'h31 == _match_key_bytes_15_T_1 ? phv_data_49 : _GEN_1344; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1346 = 8'h32 == _match_key_bytes_15_T_1 ? phv_data_50 : _GEN_1345; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1347 = 8'h33 == _match_key_bytes_15_T_1 ? phv_data_51 : _GEN_1346; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1348 = 8'h34 == _match_key_bytes_15_T_1 ? phv_data_52 : _GEN_1347; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1349 = 8'h35 == _match_key_bytes_15_T_1 ? phv_data_53 : _GEN_1348; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1350 = 8'h36 == _match_key_bytes_15_T_1 ? phv_data_54 : _GEN_1349; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1351 = 8'h37 == _match_key_bytes_15_T_1 ? phv_data_55 : _GEN_1350; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1352 = 8'h38 == _match_key_bytes_15_T_1 ? phv_data_56 : _GEN_1351; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1353 = 8'h39 == _match_key_bytes_15_T_1 ? phv_data_57 : _GEN_1352; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1354 = 8'h3a == _match_key_bytes_15_T_1 ? phv_data_58 : _GEN_1353; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1355 = 8'h3b == _match_key_bytes_15_T_1 ? phv_data_59 : _GEN_1354; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1356 = 8'h3c == _match_key_bytes_15_T_1 ? phv_data_60 : _GEN_1355; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1357 = 8'h3d == _match_key_bytes_15_T_1 ? phv_data_61 : _GEN_1356; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1358 = 8'h3e == _match_key_bytes_15_T_1 ? phv_data_62 : _GEN_1357; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1359 = 8'h3f == _match_key_bytes_15_T_1 ? phv_data_63 : _GEN_1358; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1360 = 8'h40 == _match_key_bytes_15_T_1 ? phv_data_64 : _GEN_1359; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1361 = 8'h41 == _match_key_bytes_15_T_1 ? phv_data_65 : _GEN_1360; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1362 = 8'h42 == _match_key_bytes_15_T_1 ? phv_data_66 : _GEN_1361; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1363 = 8'h43 == _match_key_bytes_15_T_1 ? phv_data_67 : _GEN_1362; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1364 = 8'h44 == _match_key_bytes_15_T_1 ? phv_data_68 : _GEN_1363; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1365 = 8'h45 == _match_key_bytes_15_T_1 ? phv_data_69 : _GEN_1364; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1366 = 8'h46 == _match_key_bytes_15_T_1 ? phv_data_70 : _GEN_1365; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1367 = 8'h47 == _match_key_bytes_15_T_1 ? phv_data_71 : _GEN_1366; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1368 = 8'h48 == _match_key_bytes_15_T_1 ? phv_data_72 : _GEN_1367; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1369 = 8'h49 == _match_key_bytes_15_T_1 ? phv_data_73 : _GEN_1368; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1370 = 8'h4a == _match_key_bytes_15_T_1 ? phv_data_74 : _GEN_1369; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1371 = 8'h4b == _match_key_bytes_15_T_1 ? phv_data_75 : _GEN_1370; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1372 = 8'h4c == _match_key_bytes_15_T_1 ? phv_data_76 : _GEN_1371; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1373 = 8'h4d == _match_key_bytes_15_T_1 ? phv_data_77 : _GEN_1372; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1374 = 8'h4e == _match_key_bytes_15_T_1 ? phv_data_78 : _GEN_1373; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1375 = 8'h4f == _match_key_bytes_15_T_1 ? phv_data_79 : _GEN_1374; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1376 = 8'h50 == _match_key_bytes_15_T_1 ? phv_data_80 : _GEN_1375; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1377 = 8'h51 == _match_key_bytes_15_T_1 ? phv_data_81 : _GEN_1376; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1378 = 8'h52 == _match_key_bytes_15_T_1 ? phv_data_82 : _GEN_1377; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1379 = 8'h53 == _match_key_bytes_15_T_1 ? phv_data_83 : _GEN_1378; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1380 = 8'h54 == _match_key_bytes_15_T_1 ? phv_data_84 : _GEN_1379; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1381 = 8'h55 == _match_key_bytes_15_T_1 ? phv_data_85 : _GEN_1380; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1382 = 8'h56 == _match_key_bytes_15_T_1 ? phv_data_86 : _GEN_1381; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1383 = 8'h57 == _match_key_bytes_15_T_1 ? phv_data_87 : _GEN_1382; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1384 = 8'h58 == _match_key_bytes_15_T_1 ? phv_data_88 : _GEN_1383; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1385 = 8'h59 == _match_key_bytes_15_T_1 ? phv_data_89 : _GEN_1384; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1386 = 8'h5a == _match_key_bytes_15_T_1 ? phv_data_90 : _GEN_1385; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1387 = 8'h5b == _match_key_bytes_15_T_1 ? phv_data_91 : _GEN_1386; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1388 = 8'h5c == _match_key_bytes_15_T_1 ? phv_data_92 : _GEN_1387; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1389 = 8'h5d == _match_key_bytes_15_T_1 ? phv_data_93 : _GEN_1388; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1390 = 8'h5e == _match_key_bytes_15_T_1 ? phv_data_94 : _GEN_1389; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1391 = 8'h5f == _match_key_bytes_15_T_1 ? phv_data_95 : _GEN_1390; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1392 = 8'h60 == _match_key_bytes_15_T_1 ? phv_data_96 : _GEN_1391; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1393 = 8'h61 == _match_key_bytes_15_T_1 ? phv_data_97 : _GEN_1392; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1394 = 8'h62 == _match_key_bytes_15_T_1 ? phv_data_98 : _GEN_1393; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1395 = 8'h63 == _match_key_bytes_15_T_1 ? phv_data_99 : _GEN_1394; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1396 = 8'h64 == _match_key_bytes_15_T_1 ? phv_data_100 : _GEN_1395; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1397 = 8'h65 == _match_key_bytes_15_T_1 ? phv_data_101 : _GEN_1396; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1398 = 8'h66 == _match_key_bytes_15_T_1 ? phv_data_102 : _GEN_1397; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1399 = 8'h67 == _match_key_bytes_15_T_1 ? phv_data_103 : _GEN_1398; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1400 = 8'h68 == _match_key_bytes_15_T_1 ? phv_data_104 : _GEN_1399; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1401 = 8'h69 == _match_key_bytes_15_T_1 ? phv_data_105 : _GEN_1400; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1402 = 8'h6a == _match_key_bytes_15_T_1 ? phv_data_106 : _GEN_1401; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1403 = 8'h6b == _match_key_bytes_15_T_1 ? phv_data_107 : _GEN_1402; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1404 = 8'h6c == _match_key_bytes_15_T_1 ? phv_data_108 : _GEN_1403; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1405 = 8'h6d == _match_key_bytes_15_T_1 ? phv_data_109 : _GEN_1404; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1406 = 8'h6e == _match_key_bytes_15_T_1 ? phv_data_110 : _GEN_1405; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1407 = 8'h6f == _match_key_bytes_15_T_1 ? phv_data_111 : _GEN_1406; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1408 = 8'h70 == _match_key_bytes_15_T_1 ? phv_data_112 : _GEN_1407; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1409 = 8'h71 == _match_key_bytes_15_T_1 ? phv_data_113 : _GEN_1408; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1410 = 8'h72 == _match_key_bytes_15_T_1 ? phv_data_114 : _GEN_1409; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1411 = 8'h73 == _match_key_bytes_15_T_1 ? phv_data_115 : _GEN_1410; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1412 = 8'h74 == _match_key_bytes_15_T_1 ? phv_data_116 : _GEN_1411; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1413 = 8'h75 == _match_key_bytes_15_T_1 ? phv_data_117 : _GEN_1412; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1414 = 8'h76 == _match_key_bytes_15_T_1 ? phv_data_118 : _GEN_1413; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1415 = 8'h77 == _match_key_bytes_15_T_1 ? phv_data_119 : _GEN_1414; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1416 = 8'h78 == _match_key_bytes_15_T_1 ? phv_data_120 : _GEN_1415; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1417 = 8'h79 == _match_key_bytes_15_T_1 ? phv_data_121 : _GEN_1416; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1418 = 8'h7a == _match_key_bytes_15_T_1 ? phv_data_122 : _GEN_1417; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1419 = 8'h7b == _match_key_bytes_15_T_1 ? phv_data_123 : _GEN_1418; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1420 = 8'h7c == _match_key_bytes_15_T_1 ? phv_data_124 : _GEN_1419; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1421 = 8'h7d == _match_key_bytes_15_T_1 ? phv_data_125 : _GEN_1420; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1422 = 8'h7e == _match_key_bytes_15_T_1 ? phv_data_126 : _GEN_1421; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1423 = 8'h7f == _match_key_bytes_15_T_1 ? phv_data_127 : _GEN_1422; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1424 = 8'h80 == _match_key_bytes_15_T_1 ? phv_data_128 : _GEN_1423; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1425 = 8'h81 == _match_key_bytes_15_T_1 ? phv_data_129 : _GEN_1424; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1426 = 8'h82 == _match_key_bytes_15_T_1 ? phv_data_130 : _GEN_1425; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1427 = 8'h83 == _match_key_bytes_15_T_1 ? phv_data_131 : _GEN_1426; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1428 = 8'h84 == _match_key_bytes_15_T_1 ? phv_data_132 : _GEN_1427; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1429 = 8'h85 == _match_key_bytes_15_T_1 ? phv_data_133 : _GEN_1428; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1430 = 8'h86 == _match_key_bytes_15_T_1 ? phv_data_134 : _GEN_1429; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1431 = 8'h87 == _match_key_bytes_15_T_1 ? phv_data_135 : _GEN_1430; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1432 = 8'h88 == _match_key_bytes_15_T_1 ? phv_data_136 : _GEN_1431; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1433 = 8'h89 == _match_key_bytes_15_T_1 ? phv_data_137 : _GEN_1432; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1434 = 8'h8a == _match_key_bytes_15_T_1 ? phv_data_138 : _GEN_1433; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1435 = 8'h8b == _match_key_bytes_15_T_1 ? phv_data_139 : _GEN_1434; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1436 = 8'h8c == _match_key_bytes_15_T_1 ? phv_data_140 : _GEN_1435; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1437 = 8'h8d == _match_key_bytes_15_T_1 ? phv_data_141 : _GEN_1436; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1438 = 8'h8e == _match_key_bytes_15_T_1 ? phv_data_142 : _GEN_1437; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1439 = 8'h8f == _match_key_bytes_15_T_1 ? phv_data_143 : _GEN_1438; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1440 = 8'h90 == _match_key_bytes_15_T_1 ? phv_data_144 : _GEN_1439; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1441 = 8'h91 == _match_key_bytes_15_T_1 ? phv_data_145 : _GEN_1440; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1442 = 8'h92 == _match_key_bytes_15_T_1 ? phv_data_146 : _GEN_1441; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1443 = 8'h93 == _match_key_bytes_15_T_1 ? phv_data_147 : _GEN_1442; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1444 = 8'h94 == _match_key_bytes_15_T_1 ? phv_data_148 : _GEN_1443; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1445 = 8'h95 == _match_key_bytes_15_T_1 ? phv_data_149 : _GEN_1444; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1446 = 8'h96 == _match_key_bytes_15_T_1 ? phv_data_150 : _GEN_1445; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1447 = 8'h97 == _match_key_bytes_15_T_1 ? phv_data_151 : _GEN_1446; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1448 = 8'h98 == _match_key_bytes_15_T_1 ? phv_data_152 : _GEN_1447; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1449 = 8'h99 == _match_key_bytes_15_T_1 ? phv_data_153 : _GEN_1448; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1450 = 8'h9a == _match_key_bytes_15_T_1 ? phv_data_154 : _GEN_1449; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1451 = 8'h9b == _match_key_bytes_15_T_1 ? phv_data_155 : _GEN_1450; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1452 = 8'h9c == _match_key_bytes_15_T_1 ? phv_data_156 : _GEN_1451; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1453 = 8'h9d == _match_key_bytes_15_T_1 ? phv_data_157 : _GEN_1452; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1454 = 8'h9e == _match_key_bytes_15_T_1 ? phv_data_158 : _GEN_1453; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1455 = 8'h9f == _match_key_bytes_15_T_1 ? phv_data_159 : _GEN_1454; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_15 = 8'h8 < _GEN_6 ? _GEN_1455 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_14_T_1 = key_offset + 8'h9; // @[matcher.scala 72:98]
  wire [7:0] _GEN_1458 = 8'h1 == _match_key_bytes_14_T_1 ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1459 = 8'h2 == _match_key_bytes_14_T_1 ? phv_data_2 : _GEN_1458; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1460 = 8'h3 == _match_key_bytes_14_T_1 ? phv_data_3 : _GEN_1459; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1461 = 8'h4 == _match_key_bytes_14_T_1 ? phv_data_4 : _GEN_1460; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1462 = 8'h5 == _match_key_bytes_14_T_1 ? phv_data_5 : _GEN_1461; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1463 = 8'h6 == _match_key_bytes_14_T_1 ? phv_data_6 : _GEN_1462; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1464 = 8'h7 == _match_key_bytes_14_T_1 ? phv_data_7 : _GEN_1463; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1465 = 8'h8 == _match_key_bytes_14_T_1 ? phv_data_8 : _GEN_1464; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1466 = 8'h9 == _match_key_bytes_14_T_1 ? phv_data_9 : _GEN_1465; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1467 = 8'ha == _match_key_bytes_14_T_1 ? phv_data_10 : _GEN_1466; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1468 = 8'hb == _match_key_bytes_14_T_1 ? phv_data_11 : _GEN_1467; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1469 = 8'hc == _match_key_bytes_14_T_1 ? phv_data_12 : _GEN_1468; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1470 = 8'hd == _match_key_bytes_14_T_1 ? phv_data_13 : _GEN_1469; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1471 = 8'he == _match_key_bytes_14_T_1 ? phv_data_14 : _GEN_1470; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1472 = 8'hf == _match_key_bytes_14_T_1 ? phv_data_15 : _GEN_1471; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1473 = 8'h10 == _match_key_bytes_14_T_1 ? phv_data_16 : _GEN_1472; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1474 = 8'h11 == _match_key_bytes_14_T_1 ? phv_data_17 : _GEN_1473; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1475 = 8'h12 == _match_key_bytes_14_T_1 ? phv_data_18 : _GEN_1474; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1476 = 8'h13 == _match_key_bytes_14_T_1 ? phv_data_19 : _GEN_1475; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1477 = 8'h14 == _match_key_bytes_14_T_1 ? phv_data_20 : _GEN_1476; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1478 = 8'h15 == _match_key_bytes_14_T_1 ? phv_data_21 : _GEN_1477; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1479 = 8'h16 == _match_key_bytes_14_T_1 ? phv_data_22 : _GEN_1478; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1480 = 8'h17 == _match_key_bytes_14_T_1 ? phv_data_23 : _GEN_1479; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1481 = 8'h18 == _match_key_bytes_14_T_1 ? phv_data_24 : _GEN_1480; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1482 = 8'h19 == _match_key_bytes_14_T_1 ? phv_data_25 : _GEN_1481; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1483 = 8'h1a == _match_key_bytes_14_T_1 ? phv_data_26 : _GEN_1482; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1484 = 8'h1b == _match_key_bytes_14_T_1 ? phv_data_27 : _GEN_1483; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1485 = 8'h1c == _match_key_bytes_14_T_1 ? phv_data_28 : _GEN_1484; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1486 = 8'h1d == _match_key_bytes_14_T_1 ? phv_data_29 : _GEN_1485; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1487 = 8'h1e == _match_key_bytes_14_T_1 ? phv_data_30 : _GEN_1486; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1488 = 8'h1f == _match_key_bytes_14_T_1 ? phv_data_31 : _GEN_1487; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1489 = 8'h20 == _match_key_bytes_14_T_1 ? phv_data_32 : _GEN_1488; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1490 = 8'h21 == _match_key_bytes_14_T_1 ? phv_data_33 : _GEN_1489; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1491 = 8'h22 == _match_key_bytes_14_T_1 ? phv_data_34 : _GEN_1490; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1492 = 8'h23 == _match_key_bytes_14_T_1 ? phv_data_35 : _GEN_1491; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1493 = 8'h24 == _match_key_bytes_14_T_1 ? phv_data_36 : _GEN_1492; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1494 = 8'h25 == _match_key_bytes_14_T_1 ? phv_data_37 : _GEN_1493; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1495 = 8'h26 == _match_key_bytes_14_T_1 ? phv_data_38 : _GEN_1494; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1496 = 8'h27 == _match_key_bytes_14_T_1 ? phv_data_39 : _GEN_1495; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1497 = 8'h28 == _match_key_bytes_14_T_1 ? phv_data_40 : _GEN_1496; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1498 = 8'h29 == _match_key_bytes_14_T_1 ? phv_data_41 : _GEN_1497; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1499 = 8'h2a == _match_key_bytes_14_T_1 ? phv_data_42 : _GEN_1498; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1500 = 8'h2b == _match_key_bytes_14_T_1 ? phv_data_43 : _GEN_1499; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1501 = 8'h2c == _match_key_bytes_14_T_1 ? phv_data_44 : _GEN_1500; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1502 = 8'h2d == _match_key_bytes_14_T_1 ? phv_data_45 : _GEN_1501; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1503 = 8'h2e == _match_key_bytes_14_T_1 ? phv_data_46 : _GEN_1502; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1504 = 8'h2f == _match_key_bytes_14_T_1 ? phv_data_47 : _GEN_1503; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1505 = 8'h30 == _match_key_bytes_14_T_1 ? phv_data_48 : _GEN_1504; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1506 = 8'h31 == _match_key_bytes_14_T_1 ? phv_data_49 : _GEN_1505; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1507 = 8'h32 == _match_key_bytes_14_T_1 ? phv_data_50 : _GEN_1506; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1508 = 8'h33 == _match_key_bytes_14_T_1 ? phv_data_51 : _GEN_1507; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1509 = 8'h34 == _match_key_bytes_14_T_1 ? phv_data_52 : _GEN_1508; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1510 = 8'h35 == _match_key_bytes_14_T_1 ? phv_data_53 : _GEN_1509; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1511 = 8'h36 == _match_key_bytes_14_T_1 ? phv_data_54 : _GEN_1510; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1512 = 8'h37 == _match_key_bytes_14_T_1 ? phv_data_55 : _GEN_1511; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1513 = 8'h38 == _match_key_bytes_14_T_1 ? phv_data_56 : _GEN_1512; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1514 = 8'h39 == _match_key_bytes_14_T_1 ? phv_data_57 : _GEN_1513; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1515 = 8'h3a == _match_key_bytes_14_T_1 ? phv_data_58 : _GEN_1514; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1516 = 8'h3b == _match_key_bytes_14_T_1 ? phv_data_59 : _GEN_1515; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1517 = 8'h3c == _match_key_bytes_14_T_1 ? phv_data_60 : _GEN_1516; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1518 = 8'h3d == _match_key_bytes_14_T_1 ? phv_data_61 : _GEN_1517; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1519 = 8'h3e == _match_key_bytes_14_T_1 ? phv_data_62 : _GEN_1518; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1520 = 8'h3f == _match_key_bytes_14_T_1 ? phv_data_63 : _GEN_1519; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1521 = 8'h40 == _match_key_bytes_14_T_1 ? phv_data_64 : _GEN_1520; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1522 = 8'h41 == _match_key_bytes_14_T_1 ? phv_data_65 : _GEN_1521; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1523 = 8'h42 == _match_key_bytes_14_T_1 ? phv_data_66 : _GEN_1522; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1524 = 8'h43 == _match_key_bytes_14_T_1 ? phv_data_67 : _GEN_1523; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1525 = 8'h44 == _match_key_bytes_14_T_1 ? phv_data_68 : _GEN_1524; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1526 = 8'h45 == _match_key_bytes_14_T_1 ? phv_data_69 : _GEN_1525; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1527 = 8'h46 == _match_key_bytes_14_T_1 ? phv_data_70 : _GEN_1526; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1528 = 8'h47 == _match_key_bytes_14_T_1 ? phv_data_71 : _GEN_1527; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1529 = 8'h48 == _match_key_bytes_14_T_1 ? phv_data_72 : _GEN_1528; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1530 = 8'h49 == _match_key_bytes_14_T_1 ? phv_data_73 : _GEN_1529; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1531 = 8'h4a == _match_key_bytes_14_T_1 ? phv_data_74 : _GEN_1530; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1532 = 8'h4b == _match_key_bytes_14_T_1 ? phv_data_75 : _GEN_1531; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1533 = 8'h4c == _match_key_bytes_14_T_1 ? phv_data_76 : _GEN_1532; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1534 = 8'h4d == _match_key_bytes_14_T_1 ? phv_data_77 : _GEN_1533; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1535 = 8'h4e == _match_key_bytes_14_T_1 ? phv_data_78 : _GEN_1534; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1536 = 8'h4f == _match_key_bytes_14_T_1 ? phv_data_79 : _GEN_1535; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1537 = 8'h50 == _match_key_bytes_14_T_1 ? phv_data_80 : _GEN_1536; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1538 = 8'h51 == _match_key_bytes_14_T_1 ? phv_data_81 : _GEN_1537; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1539 = 8'h52 == _match_key_bytes_14_T_1 ? phv_data_82 : _GEN_1538; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1540 = 8'h53 == _match_key_bytes_14_T_1 ? phv_data_83 : _GEN_1539; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1541 = 8'h54 == _match_key_bytes_14_T_1 ? phv_data_84 : _GEN_1540; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1542 = 8'h55 == _match_key_bytes_14_T_1 ? phv_data_85 : _GEN_1541; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1543 = 8'h56 == _match_key_bytes_14_T_1 ? phv_data_86 : _GEN_1542; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1544 = 8'h57 == _match_key_bytes_14_T_1 ? phv_data_87 : _GEN_1543; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1545 = 8'h58 == _match_key_bytes_14_T_1 ? phv_data_88 : _GEN_1544; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1546 = 8'h59 == _match_key_bytes_14_T_1 ? phv_data_89 : _GEN_1545; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1547 = 8'h5a == _match_key_bytes_14_T_1 ? phv_data_90 : _GEN_1546; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1548 = 8'h5b == _match_key_bytes_14_T_1 ? phv_data_91 : _GEN_1547; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1549 = 8'h5c == _match_key_bytes_14_T_1 ? phv_data_92 : _GEN_1548; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1550 = 8'h5d == _match_key_bytes_14_T_1 ? phv_data_93 : _GEN_1549; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1551 = 8'h5e == _match_key_bytes_14_T_1 ? phv_data_94 : _GEN_1550; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1552 = 8'h5f == _match_key_bytes_14_T_1 ? phv_data_95 : _GEN_1551; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1553 = 8'h60 == _match_key_bytes_14_T_1 ? phv_data_96 : _GEN_1552; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1554 = 8'h61 == _match_key_bytes_14_T_1 ? phv_data_97 : _GEN_1553; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1555 = 8'h62 == _match_key_bytes_14_T_1 ? phv_data_98 : _GEN_1554; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1556 = 8'h63 == _match_key_bytes_14_T_1 ? phv_data_99 : _GEN_1555; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1557 = 8'h64 == _match_key_bytes_14_T_1 ? phv_data_100 : _GEN_1556; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1558 = 8'h65 == _match_key_bytes_14_T_1 ? phv_data_101 : _GEN_1557; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1559 = 8'h66 == _match_key_bytes_14_T_1 ? phv_data_102 : _GEN_1558; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1560 = 8'h67 == _match_key_bytes_14_T_1 ? phv_data_103 : _GEN_1559; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1561 = 8'h68 == _match_key_bytes_14_T_1 ? phv_data_104 : _GEN_1560; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1562 = 8'h69 == _match_key_bytes_14_T_1 ? phv_data_105 : _GEN_1561; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1563 = 8'h6a == _match_key_bytes_14_T_1 ? phv_data_106 : _GEN_1562; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1564 = 8'h6b == _match_key_bytes_14_T_1 ? phv_data_107 : _GEN_1563; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1565 = 8'h6c == _match_key_bytes_14_T_1 ? phv_data_108 : _GEN_1564; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1566 = 8'h6d == _match_key_bytes_14_T_1 ? phv_data_109 : _GEN_1565; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1567 = 8'h6e == _match_key_bytes_14_T_1 ? phv_data_110 : _GEN_1566; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1568 = 8'h6f == _match_key_bytes_14_T_1 ? phv_data_111 : _GEN_1567; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1569 = 8'h70 == _match_key_bytes_14_T_1 ? phv_data_112 : _GEN_1568; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1570 = 8'h71 == _match_key_bytes_14_T_1 ? phv_data_113 : _GEN_1569; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1571 = 8'h72 == _match_key_bytes_14_T_1 ? phv_data_114 : _GEN_1570; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1572 = 8'h73 == _match_key_bytes_14_T_1 ? phv_data_115 : _GEN_1571; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1573 = 8'h74 == _match_key_bytes_14_T_1 ? phv_data_116 : _GEN_1572; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1574 = 8'h75 == _match_key_bytes_14_T_1 ? phv_data_117 : _GEN_1573; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1575 = 8'h76 == _match_key_bytes_14_T_1 ? phv_data_118 : _GEN_1574; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1576 = 8'h77 == _match_key_bytes_14_T_1 ? phv_data_119 : _GEN_1575; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1577 = 8'h78 == _match_key_bytes_14_T_1 ? phv_data_120 : _GEN_1576; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1578 = 8'h79 == _match_key_bytes_14_T_1 ? phv_data_121 : _GEN_1577; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1579 = 8'h7a == _match_key_bytes_14_T_1 ? phv_data_122 : _GEN_1578; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1580 = 8'h7b == _match_key_bytes_14_T_1 ? phv_data_123 : _GEN_1579; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1581 = 8'h7c == _match_key_bytes_14_T_1 ? phv_data_124 : _GEN_1580; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1582 = 8'h7d == _match_key_bytes_14_T_1 ? phv_data_125 : _GEN_1581; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1583 = 8'h7e == _match_key_bytes_14_T_1 ? phv_data_126 : _GEN_1582; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1584 = 8'h7f == _match_key_bytes_14_T_1 ? phv_data_127 : _GEN_1583; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1585 = 8'h80 == _match_key_bytes_14_T_1 ? phv_data_128 : _GEN_1584; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1586 = 8'h81 == _match_key_bytes_14_T_1 ? phv_data_129 : _GEN_1585; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1587 = 8'h82 == _match_key_bytes_14_T_1 ? phv_data_130 : _GEN_1586; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1588 = 8'h83 == _match_key_bytes_14_T_1 ? phv_data_131 : _GEN_1587; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1589 = 8'h84 == _match_key_bytes_14_T_1 ? phv_data_132 : _GEN_1588; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1590 = 8'h85 == _match_key_bytes_14_T_1 ? phv_data_133 : _GEN_1589; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1591 = 8'h86 == _match_key_bytes_14_T_1 ? phv_data_134 : _GEN_1590; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1592 = 8'h87 == _match_key_bytes_14_T_1 ? phv_data_135 : _GEN_1591; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1593 = 8'h88 == _match_key_bytes_14_T_1 ? phv_data_136 : _GEN_1592; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1594 = 8'h89 == _match_key_bytes_14_T_1 ? phv_data_137 : _GEN_1593; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1595 = 8'h8a == _match_key_bytes_14_T_1 ? phv_data_138 : _GEN_1594; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1596 = 8'h8b == _match_key_bytes_14_T_1 ? phv_data_139 : _GEN_1595; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1597 = 8'h8c == _match_key_bytes_14_T_1 ? phv_data_140 : _GEN_1596; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1598 = 8'h8d == _match_key_bytes_14_T_1 ? phv_data_141 : _GEN_1597; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1599 = 8'h8e == _match_key_bytes_14_T_1 ? phv_data_142 : _GEN_1598; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1600 = 8'h8f == _match_key_bytes_14_T_1 ? phv_data_143 : _GEN_1599; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1601 = 8'h90 == _match_key_bytes_14_T_1 ? phv_data_144 : _GEN_1600; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1602 = 8'h91 == _match_key_bytes_14_T_1 ? phv_data_145 : _GEN_1601; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1603 = 8'h92 == _match_key_bytes_14_T_1 ? phv_data_146 : _GEN_1602; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1604 = 8'h93 == _match_key_bytes_14_T_1 ? phv_data_147 : _GEN_1603; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1605 = 8'h94 == _match_key_bytes_14_T_1 ? phv_data_148 : _GEN_1604; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1606 = 8'h95 == _match_key_bytes_14_T_1 ? phv_data_149 : _GEN_1605; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1607 = 8'h96 == _match_key_bytes_14_T_1 ? phv_data_150 : _GEN_1606; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1608 = 8'h97 == _match_key_bytes_14_T_1 ? phv_data_151 : _GEN_1607; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1609 = 8'h98 == _match_key_bytes_14_T_1 ? phv_data_152 : _GEN_1608; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1610 = 8'h99 == _match_key_bytes_14_T_1 ? phv_data_153 : _GEN_1609; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1611 = 8'h9a == _match_key_bytes_14_T_1 ? phv_data_154 : _GEN_1610; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1612 = 8'h9b == _match_key_bytes_14_T_1 ? phv_data_155 : _GEN_1611; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1613 = 8'h9c == _match_key_bytes_14_T_1 ? phv_data_156 : _GEN_1612; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1614 = 8'h9d == _match_key_bytes_14_T_1 ? phv_data_157 : _GEN_1613; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1615 = 8'h9e == _match_key_bytes_14_T_1 ? phv_data_158 : _GEN_1614; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1616 = 8'h9f == _match_key_bytes_14_T_1 ? phv_data_159 : _GEN_1615; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_14 = 8'h9 < _GEN_6 ? _GEN_1616 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_13_T_1 = key_offset + 8'ha; // @[matcher.scala 72:98]
  wire [7:0] _GEN_1619 = 8'h1 == _match_key_bytes_13_T_1 ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1620 = 8'h2 == _match_key_bytes_13_T_1 ? phv_data_2 : _GEN_1619; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1621 = 8'h3 == _match_key_bytes_13_T_1 ? phv_data_3 : _GEN_1620; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1622 = 8'h4 == _match_key_bytes_13_T_1 ? phv_data_4 : _GEN_1621; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1623 = 8'h5 == _match_key_bytes_13_T_1 ? phv_data_5 : _GEN_1622; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1624 = 8'h6 == _match_key_bytes_13_T_1 ? phv_data_6 : _GEN_1623; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1625 = 8'h7 == _match_key_bytes_13_T_1 ? phv_data_7 : _GEN_1624; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1626 = 8'h8 == _match_key_bytes_13_T_1 ? phv_data_8 : _GEN_1625; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1627 = 8'h9 == _match_key_bytes_13_T_1 ? phv_data_9 : _GEN_1626; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1628 = 8'ha == _match_key_bytes_13_T_1 ? phv_data_10 : _GEN_1627; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1629 = 8'hb == _match_key_bytes_13_T_1 ? phv_data_11 : _GEN_1628; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1630 = 8'hc == _match_key_bytes_13_T_1 ? phv_data_12 : _GEN_1629; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1631 = 8'hd == _match_key_bytes_13_T_1 ? phv_data_13 : _GEN_1630; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1632 = 8'he == _match_key_bytes_13_T_1 ? phv_data_14 : _GEN_1631; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1633 = 8'hf == _match_key_bytes_13_T_1 ? phv_data_15 : _GEN_1632; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1634 = 8'h10 == _match_key_bytes_13_T_1 ? phv_data_16 : _GEN_1633; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1635 = 8'h11 == _match_key_bytes_13_T_1 ? phv_data_17 : _GEN_1634; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1636 = 8'h12 == _match_key_bytes_13_T_1 ? phv_data_18 : _GEN_1635; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1637 = 8'h13 == _match_key_bytes_13_T_1 ? phv_data_19 : _GEN_1636; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1638 = 8'h14 == _match_key_bytes_13_T_1 ? phv_data_20 : _GEN_1637; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1639 = 8'h15 == _match_key_bytes_13_T_1 ? phv_data_21 : _GEN_1638; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1640 = 8'h16 == _match_key_bytes_13_T_1 ? phv_data_22 : _GEN_1639; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1641 = 8'h17 == _match_key_bytes_13_T_1 ? phv_data_23 : _GEN_1640; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1642 = 8'h18 == _match_key_bytes_13_T_1 ? phv_data_24 : _GEN_1641; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1643 = 8'h19 == _match_key_bytes_13_T_1 ? phv_data_25 : _GEN_1642; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1644 = 8'h1a == _match_key_bytes_13_T_1 ? phv_data_26 : _GEN_1643; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1645 = 8'h1b == _match_key_bytes_13_T_1 ? phv_data_27 : _GEN_1644; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1646 = 8'h1c == _match_key_bytes_13_T_1 ? phv_data_28 : _GEN_1645; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1647 = 8'h1d == _match_key_bytes_13_T_1 ? phv_data_29 : _GEN_1646; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1648 = 8'h1e == _match_key_bytes_13_T_1 ? phv_data_30 : _GEN_1647; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1649 = 8'h1f == _match_key_bytes_13_T_1 ? phv_data_31 : _GEN_1648; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1650 = 8'h20 == _match_key_bytes_13_T_1 ? phv_data_32 : _GEN_1649; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1651 = 8'h21 == _match_key_bytes_13_T_1 ? phv_data_33 : _GEN_1650; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1652 = 8'h22 == _match_key_bytes_13_T_1 ? phv_data_34 : _GEN_1651; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1653 = 8'h23 == _match_key_bytes_13_T_1 ? phv_data_35 : _GEN_1652; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1654 = 8'h24 == _match_key_bytes_13_T_1 ? phv_data_36 : _GEN_1653; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1655 = 8'h25 == _match_key_bytes_13_T_1 ? phv_data_37 : _GEN_1654; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1656 = 8'h26 == _match_key_bytes_13_T_1 ? phv_data_38 : _GEN_1655; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1657 = 8'h27 == _match_key_bytes_13_T_1 ? phv_data_39 : _GEN_1656; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1658 = 8'h28 == _match_key_bytes_13_T_1 ? phv_data_40 : _GEN_1657; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1659 = 8'h29 == _match_key_bytes_13_T_1 ? phv_data_41 : _GEN_1658; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1660 = 8'h2a == _match_key_bytes_13_T_1 ? phv_data_42 : _GEN_1659; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1661 = 8'h2b == _match_key_bytes_13_T_1 ? phv_data_43 : _GEN_1660; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1662 = 8'h2c == _match_key_bytes_13_T_1 ? phv_data_44 : _GEN_1661; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1663 = 8'h2d == _match_key_bytes_13_T_1 ? phv_data_45 : _GEN_1662; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1664 = 8'h2e == _match_key_bytes_13_T_1 ? phv_data_46 : _GEN_1663; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1665 = 8'h2f == _match_key_bytes_13_T_1 ? phv_data_47 : _GEN_1664; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1666 = 8'h30 == _match_key_bytes_13_T_1 ? phv_data_48 : _GEN_1665; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1667 = 8'h31 == _match_key_bytes_13_T_1 ? phv_data_49 : _GEN_1666; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1668 = 8'h32 == _match_key_bytes_13_T_1 ? phv_data_50 : _GEN_1667; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1669 = 8'h33 == _match_key_bytes_13_T_1 ? phv_data_51 : _GEN_1668; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1670 = 8'h34 == _match_key_bytes_13_T_1 ? phv_data_52 : _GEN_1669; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1671 = 8'h35 == _match_key_bytes_13_T_1 ? phv_data_53 : _GEN_1670; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1672 = 8'h36 == _match_key_bytes_13_T_1 ? phv_data_54 : _GEN_1671; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1673 = 8'h37 == _match_key_bytes_13_T_1 ? phv_data_55 : _GEN_1672; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1674 = 8'h38 == _match_key_bytes_13_T_1 ? phv_data_56 : _GEN_1673; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1675 = 8'h39 == _match_key_bytes_13_T_1 ? phv_data_57 : _GEN_1674; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1676 = 8'h3a == _match_key_bytes_13_T_1 ? phv_data_58 : _GEN_1675; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1677 = 8'h3b == _match_key_bytes_13_T_1 ? phv_data_59 : _GEN_1676; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1678 = 8'h3c == _match_key_bytes_13_T_1 ? phv_data_60 : _GEN_1677; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1679 = 8'h3d == _match_key_bytes_13_T_1 ? phv_data_61 : _GEN_1678; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1680 = 8'h3e == _match_key_bytes_13_T_1 ? phv_data_62 : _GEN_1679; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1681 = 8'h3f == _match_key_bytes_13_T_1 ? phv_data_63 : _GEN_1680; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1682 = 8'h40 == _match_key_bytes_13_T_1 ? phv_data_64 : _GEN_1681; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1683 = 8'h41 == _match_key_bytes_13_T_1 ? phv_data_65 : _GEN_1682; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1684 = 8'h42 == _match_key_bytes_13_T_1 ? phv_data_66 : _GEN_1683; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1685 = 8'h43 == _match_key_bytes_13_T_1 ? phv_data_67 : _GEN_1684; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1686 = 8'h44 == _match_key_bytes_13_T_1 ? phv_data_68 : _GEN_1685; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1687 = 8'h45 == _match_key_bytes_13_T_1 ? phv_data_69 : _GEN_1686; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1688 = 8'h46 == _match_key_bytes_13_T_1 ? phv_data_70 : _GEN_1687; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1689 = 8'h47 == _match_key_bytes_13_T_1 ? phv_data_71 : _GEN_1688; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1690 = 8'h48 == _match_key_bytes_13_T_1 ? phv_data_72 : _GEN_1689; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1691 = 8'h49 == _match_key_bytes_13_T_1 ? phv_data_73 : _GEN_1690; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1692 = 8'h4a == _match_key_bytes_13_T_1 ? phv_data_74 : _GEN_1691; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1693 = 8'h4b == _match_key_bytes_13_T_1 ? phv_data_75 : _GEN_1692; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1694 = 8'h4c == _match_key_bytes_13_T_1 ? phv_data_76 : _GEN_1693; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1695 = 8'h4d == _match_key_bytes_13_T_1 ? phv_data_77 : _GEN_1694; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1696 = 8'h4e == _match_key_bytes_13_T_1 ? phv_data_78 : _GEN_1695; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1697 = 8'h4f == _match_key_bytes_13_T_1 ? phv_data_79 : _GEN_1696; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1698 = 8'h50 == _match_key_bytes_13_T_1 ? phv_data_80 : _GEN_1697; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1699 = 8'h51 == _match_key_bytes_13_T_1 ? phv_data_81 : _GEN_1698; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1700 = 8'h52 == _match_key_bytes_13_T_1 ? phv_data_82 : _GEN_1699; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1701 = 8'h53 == _match_key_bytes_13_T_1 ? phv_data_83 : _GEN_1700; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1702 = 8'h54 == _match_key_bytes_13_T_1 ? phv_data_84 : _GEN_1701; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1703 = 8'h55 == _match_key_bytes_13_T_1 ? phv_data_85 : _GEN_1702; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1704 = 8'h56 == _match_key_bytes_13_T_1 ? phv_data_86 : _GEN_1703; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1705 = 8'h57 == _match_key_bytes_13_T_1 ? phv_data_87 : _GEN_1704; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1706 = 8'h58 == _match_key_bytes_13_T_1 ? phv_data_88 : _GEN_1705; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1707 = 8'h59 == _match_key_bytes_13_T_1 ? phv_data_89 : _GEN_1706; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1708 = 8'h5a == _match_key_bytes_13_T_1 ? phv_data_90 : _GEN_1707; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1709 = 8'h5b == _match_key_bytes_13_T_1 ? phv_data_91 : _GEN_1708; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1710 = 8'h5c == _match_key_bytes_13_T_1 ? phv_data_92 : _GEN_1709; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1711 = 8'h5d == _match_key_bytes_13_T_1 ? phv_data_93 : _GEN_1710; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1712 = 8'h5e == _match_key_bytes_13_T_1 ? phv_data_94 : _GEN_1711; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1713 = 8'h5f == _match_key_bytes_13_T_1 ? phv_data_95 : _GEN_1712; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1714 = 8'h60 == _match_key_bytes_13_T_1 ? phv_data_96 : _GEN_1713; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1715 = 8'h61 == _match_key_bytes_13_T_1 ? phv_data_97 : _GEN_1714; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1716 = 8'h62 == _match_key_bytes_13_T_1 ? phv_data_98 : _GEN_1715; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1717 = 8'h63 == _match_key_bytes_13_T_1 ? phv_data_99 : _GEN_1716; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1718 = 8'h64 == _match_key_bytes_13_T_1 ? phv_data_100 : _GEN_1717; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1719 = 8'h65 == _match_key_bytes_13_T_1 ? phv_data_101 : _GEN_1718; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1720 = 8'h66 == _match_key_bytes_13_T_1 ? phv_data_102 : _GEN_1719; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1721 = 8'h67 == _match_key_bytes_13_T_1 ? phv_data_103 : _GEN_1720; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1722 = 8'h68 == _match_key_bytes_13_T_1 ? phv_data_104 : _GEN_1721; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1723 = 8'h69 == _match_key_bytes_13_T_1 ? phv_data_105 : _GEN_1722; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1724 = 8'h6a == _match_key_bytes_13_T_1 ? phv_data_106 : _GEN_1723; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1725 = 8'h6b == _match_key_bytes_13_T_1 ? phv_data_107 : _GEN_1724; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1726 = 8'h6c == _match_key_bytes_13_T_1 ? phv_data_108 : _GEN_1725; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1727 = 8'h6d == _match_key_bytes_13_T_1 ? phv_data_109 : _GEN_1726; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1728 = 8'h6e == _match_key_bytes_13_T_1 ? phv_data_110 : _GEN_1727; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1729 = 8'h6f == _match_key_bytes_13_T_1 ? phv_data_111 : _GEN_1728; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1730 = 8'h70 == _match_key_bytes_13_T_1 ? phv_data_112 : _GEN_1729; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1731 = 8'h71 == _match_key_bytes_13_T_1 ? phv_data_113 : _GEN_1730; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1732 = 8'h72 == _match_key_bytes_13_T_1 ? phv_data_114 : _GEN_1731; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1733 = 8'h73 == _match_key_bytes_13_T_1 ? phv_data_115 : _GEN_1732; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1734 = 8'h74 == _match_key_bytes_13_T_1 ? phv_data_116 : _GEN_1733; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1735 = 8'h75 == _match_key_bytes_13_T_1 ? phv_data_117 : _GEN_1734; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1736 = 8'h76 == _match_key_bytes_13_T_1 ? phv_data_118 : _GEN_1735; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1737 = 8'h77 == _match_key_bytes_13_T_1 ? phv_data_119 : _GEN_1736; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1738 = 8'h78 == _match_key_bytes_13_T_1 ? phv_data_120 : _GEN_1737; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1739 = 8'h79 == _match_key_bytes_13_T_1 ? phv_data_121 : _GEN_1738; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1740 = 8'h7a == _match_key_bytes_13_T_1 ? phv_data_122 : _GEN_1739; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1741 = 8'h7b == _match_key_bytes_13_T_1 ? phv_data_123 : _GEN_1740; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1742 = 8'h7c == _match_key_bytes_13_T_1 ? phv_data_124 : _GEN_1741; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1743 = 8'h7d == _match_key_bytes_13_T_1 ? phv_data_125 : _GEN_1742; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1744 = 8'h7e == _match_key_bytes_13_T_1 ? phv_data_126 : _GEN_1743; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1745 = 8'h7f == _match_key_bytes_13_T_1 ? phv_data_127 : _GEN_1744; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1746 = 8'h80 == _match_key_bytes_13_T_1 ? phv_data_128 : _GEN_1745; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1747 = 8'h81 == _match_key_bytes_13_T_1 ? phv_data_129 : _GEN_1746; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1748 = 8'h82 == _match_key_bytes_13_T_1 ? phv_data_130 : _GEN_1747; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1749 = 8'h83 == _match_key_bytes_13_T_1 ? phv_data_131 : _GEN_1748; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1750 = 8'h84 == _match_key_bytes_13_T_1 ? phv_data_132 : _GEN_1749; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1751 = 8'h85 == _match_key_bytes_13_T_1 ? phv_data_133 : _GEN_1750; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1752 = 8'h86 == _match_key_bytes_13_T_1 ? phv_data_134 : _GEN_1751; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1753 = 8'h87 == _match_key_bytes_13_T_1 ? phv_data_135 : _GEN_1752; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1754 = 8'h88 == _match_key_bytes_13_T_1 ? phv_data_136 : _GEN_1753; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1755 = 8'h89 == _match_key_bytes_13_T_1 ? phv_data_137 : _GEN_1754; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1756 = 8'h8a == _match_key_bytes_13_T_1 ? phv_data_138 : _GEN_1755; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1757 = 8'h8b == _match_key_bytes_13_T_1 ? phv_data_139 : _GEN_1756; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1758 = 8'h8c == _match_key_bytes_13_T_1 ? phv_data_140 : _GEN_1757; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1759 = 8'h8d == _match_key_bytes_13_T_1 ? phv_data_141 : _GEN_1758; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1760 = 8'h8e == _match_key_bytes_13_T_1 ? phv_data_142 : _GEN_1759; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1761 = 8'h8f == _match_key_bytes_13_T_1 ? phv_data_143 : _GEN_1760; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1762 = 8'h90 == _match_key_bytes_13_T_1 ? phv_data_144 : _GEN_1761; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1763 = 8'h91 == _match_key_bytes_13_T_1 ? phv_data_145 : _GEN_1762; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1764 = 8'h92 == _match_key_bytes_13_T_1 ? phv_data_146 : _GEN_1763; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1765 = 8'h93 == _match_key_bytes_13_T_1 ? phv_data_147 : _GEN_1764; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1766 = 8'h94 == _match_key_bytes_13_T_1 ? phv_data_148 : _GEN_1765; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1767 = 8'h95 == _match_key_bytes_13_T_1 ? phv_data_149 : _GEN_1766; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1768 = 8'h96 == _match_key_bytes_13_T_1 ? phv_data_150 : _GEN_1767; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1769 = 8'h97 == _match_key_bytes_13_T_1 ? phv_data_151 : _GEN_1768; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1770 = 8'h98 == _match_key_bytes_13_T_1 ? phv_data_152 : _GEN_1769; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1771 = 8'h99 == _match_key_bytes_13_T_1 ? phv_data_153 : _GEN_1770; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1772 = 8'h9a == _match_key_bytes_13_T_1 ? phv_data_154 : _GEN_1771; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1773 = 8'h9b == _match_key_bytes_13_T_1 ? phv_data_155 : _GEN_1772; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1774 = 8'h9c == _match_key_bytes_13_T_1 ? phv_data_156 : _GEN_1773; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1775 = 8'h9d == _match_key_bytes_13_T_1 ? phv_data_157 : _GEN_1774; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1776 = 8'h9e == _match_key_bytes_13_T_1 ? phv_data_158 : _GEN_1775; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1777 = 8'h9f == _match_key_bytes_13_T_1 ? phv_data_159 : _GEN_1776; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_13 = 8'ha < _GEN_6 ? _GEN_1777 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_12_T_1 = key_offset + 8'hb; // @[matcher.scala 72:98]
  wire [7:0] _GEN_1780 = 8'h1 == _match_key_bytes_12_T_1 ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1781 = 8'h2 == _match_key_bytes_12_T_1 ? phv_data_2 : _GEN_1780; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1782 = 8'h3 == _match_key_bytes_12_T_1 ? phv_data_3 : _GEN_1781; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1783 = 8'h4 == _match_key_bytes_12_T_1 ? phv_data_4 : _GEN_1782; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1784 = 8'h5 == _match_key_bytes_12_T_1 ? phv_data_5 : _GEN_1783; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1785 = 8'h6 == _match_key_bytes_12_T_1 ? phv_data_6 : _GEN_1784; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1786 = 8'h7 == _match_key_bytes_12_T_1 ? phv_data_7 : _GEN_1785; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1787 = 8'h8 == _match_key_bytes_12_T_1 ? phv_data_8 : _GEN_1786; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1788 = 8'h9 == _match_key_bytes_12_T_1 ? phv_data_9 : _GEN_1787; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1789 = 8'ha == _match_key_bytes_12_T_1 ? phv_data_10 : _GEN_1788; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1790 = 8'hb == _match_key_bytes_12_T_1 ? phv_data_11 : _GEN_1789; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1791 = 8'hc == _match_key_bytes_12_T_1 ? phv_data_12 : _GEN_1790; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1792 = 8'hd == _match_key_bytes_12_T_1 ? phv_data_13 : _GEN_1791; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1793 = 8'he == _match_key_bytes_12_T_1 ? phv_data_14 : _GEN_1792; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1794 = 8'hf == _match_key_bytes_12_T_1 ? phv_data_15 : _GEN_1793; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1795 = 8'h10 == _match_key_bytes_12_T_1 ? phv_data_16 : _GEN_1794; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1796 = 8'h11 == _match_key_bytes_12_T_1 ? phv_data_17 : _GEN_1795; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1797 = 8'h12 == _match_key_bytes_12_T_1 ? phv_data_18 : _GEN_1796; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1798 = 8'h13 == _match_key_bytes_12_T_1 ? phv_data_19 : _GEN_1797; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1799 = 8'h14 == _match_key_bytes_12_T_1 ? phv_data_20 : _GEN_1798; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1800 = 8'h15 == _match_key_bytes_12_T_1 ? phv_data_21 : _GEN_1799; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1801 = 8'h16 == _match_key_bytes_12_T_1 ? phv_data_22 : _GEN_1800; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1802 = 8'h17 == _match_key_bytes_12_T_1 ? phv_data_23 : _GEN_1801; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1803 = 8'h18 == _match_key_bytes_12_T_1 ? phv_data_24 : _GEN_1802; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1804 = 8'h19 == _match_key_bytes_12_T_1 ? phv_data_25 : _GEN_1803; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1805 = 8'h1a == _match_key_bytes_12_T_1 ? phv_data_26 : _GEN_1804; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1806 = 8'h1b == _match_key_bytes_12_T_1 ? phv_data_27 : _GEN_1805; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1807 = 8'h1c == _match_key_bytes_12_T_1 ? phv_data_28 : _GEN_1806; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1808 = 8'h1d == _match_key_bytes_12_T_1 ? phv_data_29 : _GEN_1807; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1809 = 8'h1e == _match_key_bytes_12_T_1 ? phv_data_30 : _GEN_1808; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1810 = 8'h1f == _match_key_bytes_12_T_1 ? phv_data_31 : _GEN_1809; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1811 = 8'h20 == _match_key_bytes_12_T_1 ? phv_data_32 : _GEN_1810; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1812 = 8'h21 == _match_key_bytes_12_T_1 ? phv_data_33 : _GEN_1811; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1813 = 8'h22 == _match_key_bytes_12_T_1 ? phv_data_34 : _GEN_1812; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1814 = 8'h23 == _match_key_bytes_12_T_1 ? phv_data_35 : _GEN_1813; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1815 = 8'h24 == _match_key_bytes_12_T_1 ? phv_data_36 : _GEN_1814; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1816 = 8'h25 == _match_key_bytes_12_T_1 ? phv_data_37 : _GEN_1815; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1817 = 8'h26 == _match_key_bytes_12_T_1 ? phv_data_38 : _GEN_1816; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1818 = 8'h27 == _match_key_bytes_12_T_1 ? phv_data_39 : _GEN_1817; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1819 = 8'h28 == _match_key_bytes_12_T_1 ? phv_data_40 : _GEN_1818; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1820 = 8'h29 == _match_key_bytes_12_T_1 ? phv_data_41 : _GEN_1819; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1821 = 8'h2a == _match_key_bytes_12_T_1 ? phv_data_42 : _GEN_1820; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1822 = 8'h2b == _match_key_bytes_12_T_1 ? phv_data_43 : _GEN_1821; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1823 = 8'h2c == _match_key_bytes_12_T_1 ? phv_data_44 : _GEN_1822; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1824 = 8'h2d == _match_key_bytes_12_T_1 ? phv_data_45 : _GEN_1823; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1825 = 8'h2e == _match_key_bytes_12_T_1 ? phv_data_46 : _GEN_1824; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1826 = 8'h2f == _match_key_bytes_12_T_1 ? phv_data_47 : _GEN_1825; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1827 = 8'h30 == _match_key_bytes_12_T_1 ? phv_data_48 : _GEN_1826; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1828 = 8'h31 == _match_key_bytes_12_T_1 ? phv_data_49 : _GEN_1827; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1829 = 8'h32 == _match_key_bytes_12_T_1 ? phv_data_50 : _GEN_1828; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1830 = 8'h33 == _match_key_bytes_12_T_1 ? phv_data_51 : _GEN_1829; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1831 = 8'h34 == _match_key_bytes_12_T_1 ? phv_data_52 : _GEN_1830; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1832 = 8'h35 == _match_key_bytes_12_T_1 ? phv_data_53 : _GEN_1831; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1833 = 8'h36 == _match_key_bytes_12_T_1 ? phv_data_54 : _GEN_1832; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1834 = 8'h37 == _match_key_bytes_12_T_1 ? phv_data_55 : _GEN_1833; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1835 = 8'h38 == _match_key_bytes_12_T_1 ? phv_data_56 : _GEN_1834; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1836 = 8'h39 == _match_key_bytes_12_T_1 ? phv_data_57 : _GEN_1835; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1837 = 8'h3a == _match_key_bytes_12_T_1 ? phv_data_58 : _GEN_1836; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1838 = 8'h3b == _match_key_bytes_12_T_1 ? phv_data_59 : _GEN_1837; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1839 = 8'h3c == _match_key_bytes_12_T_1 ? phv_data_60 : _GEN_1838; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1840 = 8'h3d == _match_key_bytes_12_T_1 ? phv_data_61 : _GEN_1839; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1841 = 8'h3e == _match_key_bytes_12_T_1 ? phv_data_62 : _GEN_1840; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1842 = 8'h3f == _match_key_bytes_12_T_1 ? phv_data_63 : _GEN_1841; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1843 = 8'h40 == _match_key_bytes_12_T_1 ? phv_data_64 : _GEN_1842; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1844 = 8'h41 == _match_key_bytes_12_T_1 ? phv_data_65 : _GEN_1843; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1845 = 8'h42 == _match_key_bytes_12_T_1 ? phv_data_66 : _GEN_1844; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1846 = 8'h43 == _match_key_bytes_12_T_1 ? phv_data_67 : _GEN_1845; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1847 = 8'h44 == _match_key_bytes_12_T_1 ? phv_data_68 : _GEN_1846; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1848 = 8'h45 == _match_key_bytes_12_T_1 ? phv_data_69 : _GEN_1847; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1849 = 8'h46 == _match_key_bytes_12_T_1 ? phv_data_70 : _GEN_1848; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1850 = 8'h47 == _match_key_bytes_12_T_1 ? phv_data_71 : _GEN_1849; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1851 = 8'h48 == _match_key_bytes_12_T_1 ? phv_data_72 : _GEN_1850; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1852 = 8'h49 == _match_key_bytes_12_T_1 ? phv_data_73 : _GEN_1851; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1853 = 8'h4a == _match_key_bytes_12_T_1 ? phv_data_74 : _GEN_1852; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1854 = 8'h4b == _match_key_bytes_12_T_1 ? phv_data_75 : _GEN_1853; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1855 = 8'h4c == _match_key_bytes_12_T_1 ? phv_data_76 : _GEN_1854; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1856 = 8'h4d == _match_key_bytes_12_T_1 ? phv_data_77 : _GEN_1855; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1857 = 8'h4e == _match_key_bytes_12_T_1 ? phv_data_78 : _GEN_1856; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1858 = 8'h4f == _match_key_bytes_12_T_1 ? phv_data_79 : _GEN_1857; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1859 = 8'h50 == _match_key_bytes_12_T_1 ? phv_data_80 : _GEN_1858; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1860 = 8'h51 == _match_key_bytes_12_T_1 ? phv_data_81 : _GEN_1859; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1861 = 8'h52 == _match_key_bytes_12_T_1 ? phv_data_82 : _GEN_1860; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1862 = 8'h53 == _match_key_bytes_12_T_1 ? phv_data_83 : _GEN_1861; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1863 = 8'h54 == _match_key_bytes_12_T_1 ? phv_data_84 : _GEN_1862; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1864 = 8'h55 == _match_key_bytes_12_T_1 ? phv_data_85 : _GEN_1863; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1865 = 8'h56 == _match_key_bytes_12_T_1 ? phv_data_86 : _GEN_1864; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1866 = 8'h57 == _match_key_bytes_12_T_1 ? phv_data_87 : _GEN_1865; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1867 = 8'h58 == _match_key_bytes_12_T_1 ? phv_data_88 : _GEN_1866; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1868 = 8'h59 == _match_key_bytes_12_T_1 ? phv_data_89 : _GEN_1867; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1869 = 8'h5a == _match_key_bytes_12_T_1 ? phv_data_90 : _GEN_1868; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1870 = 8'h5b == _match_key_bytes_12_T_1 ? phv_data_91 : _GEN_1869; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1871 = 8'h5c == _match_key_bytes_12_T_1 ? phv_data_92 : _GEN_1870; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1872 = 8'h5d == _match_key_bytes_12_T_1 ? phv_data_93 : _GEN_1871; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1873 = 8'h5e == _match_key_bytes_12_T_1 ? phv_data_94 : _GEN_1872; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1874 = 8'h5f == _match_key_bytes_12_T_1 ? phv_data_95 : _GEN_1873; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1875 = 8'h60 == _match_key_bytes_12_T_1 ? phv_data_96 : _GEN_1874; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1876 = 8'h61 == _match_key_bytes_12_T_1 ? phv_data_97 : _GEN_1875; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1877 = 8'h62 == _match_key_bytes_12_T_1 ? phv_data_98 : _GEN_1876; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1878 = 8'h63 == _match_key_bytes_12_T_1 ? phv_data_99 : _GEN_1877; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1879 = 8'h64 == _match_key_bytes_12_T_1 ? phv_data_100 : _GEN_1878; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1880 = 8'h65 == _match_key_bytes_12_T_1 ? phv_data_101 : _GEN_1879; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1881 = 8'h66 == _match_key_bytes_12_T_1 ? phv_data_102 : _GEN_1880; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1882 = 8'h67 == _match_key_bytes_12_T_1 ? phv_data_103 : _GEN_1881; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1883 = 8'h68 == _match_key_bytes_12_T_1 ? phv_data_104 : _GEN_1882; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1884 = 8'h69 == _match_key_bytes_12_T_1 ? phv_data_105 : _GEN_1883; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1885 = 8'h6a == _match_key_bytes_12_T_1 ? phv_data_106 : _GEN_1884; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1886 = 8'h6b == _match_key_bytes_12_T_1 ? phv_data_107 : _GEN_1885; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1887 = 8'h6c == _match_key_bytes_12_T_1 ? phv_data_108 : _GEN_1886; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1888 = 8'h6d == _match_key_bytes_12_T_1 ? phv_data_109 : _GEN_1887; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1889 = 8'h6e == _match_key_bytes_12_T_1 ? phv_data_110 : _GEN_1888; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1890 = 8'h6f == _match_key_bytes_12_T_1 ? phv_data_111 : _GEN_1889; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1891 = 8'h70 == _match_key_bytes_12_T_1 ? phv_data_112 : _GEN_1890; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1892 = 8'h71 == _match_key_bytes_12_T_1 ? phv_data_113 : _GEN_1891; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1893 = 8'h72 == _match_key_bytes_12_T_1 ? phv_data_114 : _GEN_1892; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1894 = 8'h73 == _match_key_bytes_12_T_1 ? phv_data_115 : _GEN_1893; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1895 = 8'h74 == _match_key_bytes_12_T_1 ? phv_data_116 : _GEN_1894; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1896 = 8'h75 == _match_key_bytes_12_T_1 ? phv_data_117 : _GEN_1895; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1897 = 8'h76 == _match_key_bytes_12_T_1 ? phv_data_118 : _GEN_1896; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1898 = 8'h77 == _match_key_bytes_12_T_1 ? phv_data_119 : _GEN_1897; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1899 = 8'h78 == _match_key_bytes_12_T_1 ? phv_data_120 : _GEN_1898; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1900 = 8'h79 == _match_key_bytes_12_T_1 ? phv_data_121 : _GEN_1899; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1901 = 8'h7a == _match_key_bytes_12_T_1 ? phv_data_122 : _GEN_1900; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1902 = 8'h7b == _match_key_bytes_12_T_1 ? phv_data_123 : _GEN_1901; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1903 = 8'h7c == _match_key_bytes_12_T_1 ? phv_data_124 : _GEN_1902; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1904 = 8'h7d == _match_key_bytes_12_T_1 ? phv_data_125 : _GEN_1903; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1905 = 8'h7e == _match_key_bytes_12_T_1 ? phv_data_126 : _GEN_1904; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1906 = 8'h7f == _match_key_bytes_12_T_1 ? phv_data_127 : _GEN_1905; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1907 = 8'h80 == _match_key_bytes_12_T_1 ? phv_data_128 : _GEN_1906; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1908 = 8'h81 == _match_key_bytes_12_T_1 ? phv_data_129 : _GEN_1907; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1909 = 8'h82 == _match_key_bytes_12_T_1 ? phv_data_130 : _GEN_1908; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1910 = 8'h83 == _match_key_bytes_12_T_1 ? phv_data_131 : _GEN_1909; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1911 = 8'h84 == _match_key_bytes_12_T_1 ? phv_data_132 : _GEN_1910; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1912 = 8'h85 == _match_key_bytes_12_T_1 ? phv_data_133 : _GEN_1911; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1913 = 8'h86 == _match_key_bytes_12_T_1 ? phv_data_134 : _GEN_1912; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1914 = 8'h87 == _match_key_bytes_12_T_1 ? phv_data_135 : _GEN_1913; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1915 = 8'h88 == _match_key_bytes_12_T_1 ? phv_data_136 : _GEN_1914; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1916 = 8'h89 == _match_key_bytes_12_T_1 ? phv_data_137 : _GEN_1915; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1917 = 8'h8a == _match_key_bytes_12_T_1 ? phv_data_138 : _GEN_1916; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1918 = 8'h8b == _match_key_bytes_12_T_1 ? phv_data_139 : _GEN_1917; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1919 = 8'h8c == _match_key_bytes_12_T_1 ? phv_data_140 : _GEN_1918; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1920 = 8'h8d == _match_key_bytes_12_T_1 ? phv_data_141 : _GEN_1919; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1921 = 8'h8e == _match_key_bytes_12_T_1 ? phv_data_142 : _GEN_1920; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1922 = 8'h8f == _match_key_bytes_12_T_1 ? phv_data_143 : _GEN_1921; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1923 = 8'h90 == _match_key_bytes_12_T_1 ? phv_data_144 : _GEN_1922; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1924 = 8'h91 == _match_key_bytes_12_T_1 ? phv_data_145 : _GEN_1923; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1925 = 8'h92 == _match_key_bytes_12_T_1 ? phv_data_146 : _GEN_1924; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1926 = 8'h93 == _match_key_bytes_12_T_1 ? phv_data_147 : _GEN_1925; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1927 = 8'h94 == _match_key_bytes_12_T_1 ? phv_data_148 : _GEN_1926; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1928 = 8'h95 == _match_key_bytes_12_T_1 ? phv_data_149 : _GEN_1927; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1929 = 8'h96 == _match_key_bytes_12_T_1 ? phv_data_150 : _GEN_1928; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1930 = 8'h97 == _match_key_bytes_12_T_1 ? phv_data_151 : _GEN_1929; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1931 = 8'h98 == _match_key_bytes_12_T_1 ? phv_data_152 : _GEN_1930; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1932 = 8'h99 == _match_key_bytes_12_T_1 ? phv_data_153 : _GEN_1931; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1933 = 8'h9a == _match_key_bytes_12_T_1 ? phv_data_154 : _GEN_1932; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1934 = 8'h9b == _match_key_bytes_12_T_1 ? phv_data_155 : _GEN_1933; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1935 = 8'h9c == _match_key_bytes_12_T_1 ? phv_data_156 : _GEN_1934; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1936 = 8'h9d == _match_key_bytes_12_T_1 ? phv_data_157 : _GEN_1935; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1937 = 8'h9e == _match_key_bytes_12_T_1 ? phv_data_158 : _GEN_1936; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1938 = 8'h9f == _match_key_bytes_12_T_1 ? phv_data_159 : _GEN_1937; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_12 = 8'hb < _GEN_6 ? _GEN_1938 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_11_T_1 = key_offset + 8'hc; // @[matcher.scala 72:98]
  wire [7:0] _GEN_1941 = 8'h1 == _match_key_bytes_11_T_1 ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1942 = 8'h2 == _match_key_bytes_11_T_1 ? phv_data_2 : _GEN_1941; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1943 = 8'h3 == _match_key_bytes_11_T_1 ? phv_data_3 : _GEN_1942; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1944 = 8'h4 == _match_key_bytes_11_T_1 ? phv_data_4 : _GEN_1943; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1945 = 8'h5 == _match_key_bytes_11_T_1 ? phv_data_5 : _GEN_1944; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1946 = 8'h6 == _match_key_bytes_11_T_1 ? phv_data_6 : _GEN_1945; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1947 = 8'h7 == _match_key_bytes_11_T_1 ? phv_data_7 : _GEN_1946; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1948 = 8'h8 == _match_key_bytes_11_T_1 ? phv_data_8 : _GEN_1947; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1949 = 8'h9 == _match_key_bytes_11_T_1 ? phv_data_9 : _GEN_1948; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1950 = 8'ha == _match_key_bytes_11_T_1 ? phv_data_10 : _GEN_1949; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1951 = 8'hb == _match_key_bytes_11_T_1 ? phv_data_11 : _GEN_1950; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1952 = 8'hc == _match_key_bytes_11_T_1 ? phv_data_12 : _GEN_1951; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1953 = 8'hd == _match_key_bytes_11_T_1 ? phv_data_13 : _GEN_1952; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1954 = 8'he == _match_key_bytes_11_T_1 ? phv_data_14 : _GEN_1953; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1955 = 8'hf == _match_key_bytes_11_T_1 ? phv_data_15 : _GEN_1954; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1956 = 8'h10 == _match_key_bytes_11_T_1 ? phv_data_16 : _GEN_1955; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1957 = 8'h11 == _match_key_bytes_11_T_1 ? phv_data_17 : _GEN_1956; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1958 = 8'h12 == _match_key_bytes_11_T_1 ? phv_data_18 : _GEN_1957; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1959 = 8'h13 == _match_key_bytes_11_T_1 ? phv_data_19 : _GEN_1958; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1960 = 8'h14 == _match_key_bytes_11_T_1 ? phv_data_20 : _GEN_1959; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1961 = 8'h15 == _match_key_bytes_11_T_1 ? phv_data_21 : _GEN_1960; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1962 = 8'h16 == _match_key_bytes_11_T_1 ? phv_data_22 : _GEN_1961; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1963 = 8'h17 == _match_key_bytes_11_T_1 ? phv_data_23 : _GEN_1962; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1964 = 8'h18 == _match_key_bytes_11_T_1 ? phv_data_24 : _GEN_1963; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1965 = 8'h19 == _match_key_bytes_11_T_1 ? phv_data_25 : _GEN_1964; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1966 = 8'h1a == _match_key_bytes_11_T_1 ? phv_data_26 : _GEN_1965; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1967 = 8'h1b == _match_key_bytes_11_T_1 ? phv_data_27 : _GEN_1966; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1968 = 8'h1c == _match_key_bytes_11_T_1 ? phv_data_28 : _GEN_1967; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1969 = 8'h1d == _match_key_bytes_11_T_1 ? phv_data_29 : _GEN_1968; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1970 = 8'h1e == _match_key_bytes_11_T_1 ? phv_data_30 : _GEN_1969; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1971 = 8'h1f == _match_key_bytes_11_T_1 ? phv_data_31 : _GEN_1970; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1972 = 8'h20 == _match_key_bytes_11_T_1 ? phv_data_32 : _GEN_1971; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1973 = 8'h21 == _match_key_bytes_11_T_1 ? phv_data_33 : _GEN_1972; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1974 = 8'h22 == _match_key_bytes_11_T_1 ? phv_data_34 : _GEN_1973; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1975 = 8'h23 == _match_key_bytes_11_T_1 ? phv_data_35 : _GEN_1974; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1976 = 8'h24 == _match_key_bytes_11_T_1 ? phv_data_36 : _GEN_1975; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1977 = 8'h25 == _match_key_bytes_11_T_1 ? phv_data_37 : _GEN_1976; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1978 = 8'h26 == _match_key_bytes_11_T_1 ? phv_data_38 : _GEN_1977; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1979 = 8'h27 == _match_key_bytes_11_T_1 ? phv_data_39 : _GEN_1978; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1980 = 8'h28 == _match_key_bytes_11_T_1 ? phv_data_40 : _GEN_1979; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1981 = 8'h29 == _match_key_bytes_11_T_1 ? phv_data_41 : _GEN_1980; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1982 = 8'h2a == _match_key_bytes_11_T_1 ? phv_data_42 : _GEN_1981; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1983 = 8'h2b == _match_key_bytes_11_T_1 ? phv_data_43 : _GEN_1982; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1984 = 8'h2c == _match_key_bytes_11_T_1 ? phv_data_44 : _GEN_1983; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1985 = 8'h2d == _match_key_bytes_11_T_1 ? phv_data_45 : _GEN_1984; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1986 = 8'h2e == _match_key_bytes_11_T_1 ? phv_data_46 : _GEN_1985; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1987 = 8'h2f == _match_key_bytes_11_T_1 ? phv_data_47 : _GEN_1986; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1988 = 8'h30 == _match_key_bytes_11_T_1 ? phv_data_48 : _GEN_1987; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1989 = 8'h31 == _match_key_bytes_11_T_1 ? phv_data_49 : _GEN_1988; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1990 = 8'h32 == _match_key_bytes_11_T_1 ? phv_data_50 : _GEN_1989; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1991 = 8'h33 == _match_key_bytes_11_T_1 ? phv_data_51 : _GEN_1990; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1992 = 8'h34 == _match_key_bytes_11_T_1 ? phv_data_52 : _GEN_1991; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1993 = 8'h35 == _match_key_bytes_11_T_1 ? phv_data_53 : _GEN_1992; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1994 = 8'h36 == _match_key_bytes_11_T_1 ? phv_data_54 : _GEN_1993; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1995 = 8'h37 == _match_key_bytes_11_T_1 ? phv_data_55 : _GEN_1994; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1996 = 8'h38 == _match_key_bytes_11_T_1 ? phv_data_56 : _GEN_1995; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1997 = 8'h39 == _match_key_bytes_11_T_1 ? phv_data_57 : _GEN_1996; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1998 = 8'h3a == _match_key_bytes_11_T_1 ? phv_data_58 : _GEN_1997; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_1999 = 8'h3b == _match_key_bytes_11_T_1 ? phv_data_59 : _GEN_1998; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2000 = 8'h3c == _match_key_bytes_11_T_1 ? phv_data_60 : _GEN_1999; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2001 = 8'h3d == _match_key_bytes_11_T_1 ? phv_data_61 : _GEN_2000; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2002 = 8'h3e == _match_key_bytes_11_T_1 ? phv_data_62 : _GEN_2001; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2003 = 8'h3f == _match_key_bytes_11_T_1 ? phv_data_63 : _GEN_2002; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2004 = 8'h40 == _match_key_bytes_11_T_1 ? phv_data_64 : _GEN_2003; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2005 = 8'h41 == _match_key_bytes_11_T_1 ? phv_data_65 : _GEN_2004; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2006 = 8'h42 == _match_key_bytes_11_T_1 ? phv_data_66 : _GEN_2005; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2007 = 8'h43 == _match_key_bytes_11_T_1 ? phv_data_67 : _GEN_2006; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2008 = 8'h44 == _match_key_bytes_11_T_1 ? phv_data_68 : _GEN_2007; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2009 = 8'h45 == _match_key_bytes_11_T_1 ? phv_data_69 : _GEN_2008; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2010 = 8'h46 == _match_key_bytes_11_T_1 ? phv_data_70 : _GEN_2009; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2011 = 8'h47 == _match_key_bytes_11_T_1 ? phv_data_71 : _GEN_2010; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2012 = 8'h48 == _match_key_bytes_11_T_1 ? phv_data_72 : _GEN_2011; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2013 = 8'h49 == _match_key_bytes_11_T_1 ? phv_data_73 : _GEN_2012; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2014 = 8'h4a == _match_key_bytes_11_T_1 ? phv_data_74 : _GEN_2013; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2015 = 8'h4b == _match_key_bytes_11_T_1 ? phv_data_75 : _GEN_2014; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2016 = 8'h4c == _match_key_bytes_11_T_1 ? phv_data_76 : _GEN_2015; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2017 = 8'h4d == _match_key_bytes_11_T_1 ? phv_data_77 : _GEN_2016; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2018 = 8'h4e == _match_key_bytes_11_T_1 ? phv_data_78 : _GEN_2017; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2019 = 8'h4f == _match_key_bytes_11_T_1 ? phv_data_79 : _GEN_2018; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2020 = 8'h50 == _match_key_bytes_11_T_1 ? phv_data_80 : _GEN_2019; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2021 = 8'h51 == _match_key_bytes_11_T_1 ? phv_data_81 : _GEN_2020; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2022 = 8'h52 == _match_key_bytes_11_T_1 ? phv_data_82 : _GEN_2021; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2023 = 8'h53 == _match_key_bytes_11_T_1 ? phv_data_83 : _GEN_2022; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2024 = 8'h54 == _match_key_bytes_11_T_1 ? phv_data_84 : _GEN_2023; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2025 = 8'h55 == _match_key_bytes_11_T_1 ? phv_data_85 : _GEN_2024; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2026 = 8'h56 == _match_key_bytes_11_T_1 ? phv_data_86 : _GEN_2025; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2027 = 8'h57 == _match_key_bytes_11_T_1 ? phv_data_87 : _GEN_2026; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2028 = 8'h58 == _match_key_bytes_11_T_1 ? phv_data_88 : _GEN_2027; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2029 = 8'h59 == _match_key_bytes_11_T_1 ? phv_data_89 : _GEN_2028; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2030 = 8'h5a == _match_key_bytes_11_T_1 ? phv_data_90 : _GEN_2029; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2031 = 8'h5b == _match_key_bytes_11_T_1 ? phv_data_91 : _GEN_2030; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2032 = 8'h5c == _match_key_bytes_11_T_1 ? phv_data_92 : _GEN_2031; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2033 = 8'h5d == _match_key_bytes_11_T_1 ? phv_data_93 : _GEN_2032; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2034 = 8'h5e == _match_key_bytes_11_T_1 ? phv_data_94 : _GEN_2033; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2035 = 8'h5f == _match_key_bytes_11_T_1 ? phv_data_95 : _GEN_2034; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2036 = 8'h60 == _match_key_bytes_11_T_1 ? phv_data_96 : _GEN_2035; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2037 = 8'h61 == _match_key_bytes_11_T_1 ? phv_data_97 : _GEN_2036; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2038 = 8'h62 == _match_key_bytes_11_T_1 ? phv_data_98 : _GEN_2037; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2039 = 8'h63 == _match_key_bytes_11_T_1 ? phv_data_99 : _GEN_2038; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2040 = 8'h64 == _match_key_bytes_11_T_1 ? phv_data_100 : _GEN_2039; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2041 = 8'h65 == _match_key_bytes_11_T_1 ? phv_data_101 : _GEN_2040; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2042 = 8'h66 == _match_key_bytes_11_T_1 ? phv_data_102 : _GEN_2041; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2043 = 8'h67 == _match_key_bytes_11_T_1 ? phv_data_103 : _GEN_2042; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2044 = 8'h68 == _match_key_bytes_11_T_1 ? phv_data_104 : _GEN_2043; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2045 = 8'h69 == _match_key_bytes_11_T_1 ? phv_data_105 : _GEN_2044; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2046 = 8'h6a == _match_key_bytes_11_T_1 ? phv_data_106 : _GEN_2045; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2047 = 8'h6b == _match_key_bytes_11_T_1 ? phv_data_107 : _GEN_2046; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2048 = 8'h6c == _match_key_bytes_11_T_1 ? phv_data_108 : _GEN_2047; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2049 = 8'h6d == _match_key_bytes_11_T_1 ? phv_data_109 : _GEN_2048; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2050 = 8'h6e == _match_key_bytes_11_T_1 ? phv_data_110 : _GEN_2049; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2051 = 8'h6f == _match_key_bytes_11_T_1 ? phv_data_111 : _GEN_2050; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2052 = 8'h70 == _match_key_bytes_11_T_1 ? phv_data_112 : _GEN_2051; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2053 = 8'h71 == _match_key_bytes_11_T_1 ? phv_data_113 : _GEN_2052; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2054 = 8'h72 == _match_key_bytes_11_T_1 ? phv_data_114 : _GEN_2053; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2055 = 8'h73 == _match_key_bytes_11_T_1 ? phv_data_115 : _GEN_2054; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2056 = 8'h74 == _match_key_bytes_11_T_1 ? phv_data_116 : _GEN_2055; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2057 = 8'h75 == _match_key_bytes_11_T_1 ? phv_data_117 : _GEN_2056; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2058 = 8'h76 == _match_key_bytes_11_T_1 ? phv_data_118 : _GEN_2057; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2059 = 8'h77 == _match_key_bytes_11_T_1 ? phv_data_119 : _GEN_2058; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2060 = 8'h78 == _match_key_bytes_11_T_1 ? phv_data_120 : _GEN_2059; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2061 = 8'h79 == _match_key_bytes_11_T_1 ? phv_data_121 : _GEN_2060; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2062 = 8'h7a == _match_key_bytes_11_T_1 ? phv_data_122 : _GEN_2061; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2063 = 8'h7b == _match_key_bytes_11_T_1 ? phv_data_123 : _GEN_2062; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2064 = 8'h7c == _match_key_bytes_11_T_1 ? phv_data_124 : _GEN_2063; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2065 = 8'h7d == _match_key_bytes_11_T_1 ? phv_data_125 : _GEN_2064; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2066 = 8'h7e == _match_key_bytes_11_T_1 ? phv_data_126 : _GEN_2065; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2067 = 8'h7f == _match_key_bytes_11_T_1 ? phv_data_127 : _GEN_2066; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2068 = 8'h80 == _match_key_bytes_11_T_1 ? phv_data_128 : _GEN_2067; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2069 = 8'h81 == _match_key_bytes_11_T_1 ? phv_data_129 : _GEN_2068; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2070 = 8'h82 == _match_key_bytes_11_T_1 ? phv_data_130 : _GEN_2069; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2071 = 8'h83 == _match_key_bytes_11_T_1 ? phv_data_131 : _GEN_2070; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2072 = 8'h84 == _match_key_bytes_11_T_1 ? phv_data_132 : _GEN_2071; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2073 = 8'h85 == _match_key_bytes_11_T_1 ? phv_data_133 : _GEN_2072; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2074 = 8'h86 == _match_key_bytes_11_T_1 ? phv_data_134 : _GEN_2073; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2075 = 8'h87 == _match_key_bytes_11_T_1 ? phv_data_135 : _GEN_2074; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2076 = 8'h88 == _match_key_bytes_11_T_1 ? phv_data_136 : _GEN_2075; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2077 = 8'h89 == _match_key_bytes_11_T_1 ? phv_data_137 : _GEN_2076; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2078 = 8'h8a == _match_key_bytes_11_T_1 ? phv_data_138 : _GEN_2077; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2079 = 8'h8b == _match_key_bytes_11_T_1 ? phv_data_139 : _GEN_2078; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2080 = 8'h8c == _match_key_bytes_11_T_1 ? phv_data_140 : _GEN_2079; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2081 = 8'h8d == _match_key_bytes_11_T_1 ? phv_data_141 : _GEN_2080; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2082 = 8'h8e == _match_key_bytes_11_T_1 ? phv_data_142 : _GEN_2081; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2083 = 8'h8f == _match_key_bytes_11_T_1 ? phv_data_143 : _GEN_2082; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2084 = 8'h90 == _match_key_bytes_11_T_1 ? phv_data_144 : _GEN_2083; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2085 = 8'h91 == _match_key_bytes_11_T_1 ? phv_data_145 : _GEN_2084; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2086 = 8'h92 == _match_key_bytes_11_T_1 ? phv_data_146 : _GEN_2085; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2087 = 8'h93 == _match_key_bytes_11_T_1 ? phv_data_147 : _GEN_2086; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2088 = 8'h94 == _match_key_bytes_11_T_1 ? phv_data_148 : _GEN_2087; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2089 = 8'h95 == _match_key_bytes_11_T_1 ? phv_data_149 : _GEN_2088; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2090 = 8'h96 == _match_key_bytes_11_T_1 ? phv_data_150 : _GEN_2089; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2091 = 8'h97 == _match_key_bytes_11_T_1 ? phv_data_151 : _GEN_2090; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2092 = 8'h98 == _match_key_bytes_11_T_1 ? phv_data_152 : _GEN_2091; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2093 = 8'h99 == _match_key_bytes_11_T_1 ? phv_data_153 : _GEN_2092; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2094 = 8'h9a == _match_key_bytes_11_T_1 ? phv_data_154 : _GEN_2093; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2095 = 8'h9b == _match_key_bytes_11_T_1 ? phv_data_155 : _GEN_2094; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2096 = 8'h9c == _match_key_bytes_11_T_1 ? phv_data_156 : _GEN_2095; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2097 = 8'h9d == _match_key_bytes_11_T_1 ? phv_data_157 : _GEN_2096; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2098 = 8'h9e == _match_key_bytes_11_T_1 ? phv_data_158 : _GEN_2097; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2099 = 8'h9f == _match_key_bytes_11_T_1 ? phv_data_159 : _GEN_2098; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_11 = 8'hc < _GEN_6 ? _GEN_2099 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_10_T_1 = key_offset + 8'hd; // @[matcher.scala 72:98]
  wire [7:0] _GEN_2102 = 8'h1 == _match_key_bytes_10_T_1 ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2103 = 8'h2 == _match_key_bytes_10_T_1 ? phv_data_2 : _GEN_2102; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2104 = 8'h3 == _match_key_bytes_10_T_1 ? phv_data_3 : _GEN_2103; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2105 = 8'h4 == _match_key_bytes_10_T_1 ? phv_data_4 : _GEN_2104; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2106 = 8'h5 == _match_key_bytes_10_T_1 ? phv_data_5 : _GEN_2105; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2107 = 8'h6 == _match_key_bytes_10_T_1 ? phv_data_6 : _GEN_2106; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2108 = 8'h7 == _match_key_bytes_10_T_1 ? phv_data_7 : _GEN_2107; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2109 = 8'h8 == _match_key_bytes_10_T_1 ? phv_data_8 : _GEN_2108; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2110 = 8'h9 == _match_key_bytes_10_T_1 ? phv_data_9 : _GEN_2109; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2111 = 8'ha == _match_key_bytes_10_T_1 ? phv_data_10 : _GEN_2110; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2112 = 8'hb == _match_key_bytes_10_T_1 ? phv_data_11 : _GEN_2111; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2113 = 8'hc == _match_key_bytes_10_T_1 ? phv_data_12 : _GEN_2112; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2114 = 8'hd == _match_key_bytes_10_T_1 ? phv_data_13 : _GEN_2113; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2115 = 8'he == _match_key_bytes_10_T_1 ? phv_data_14 : _GEN_2114; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2116 = 8'hf == _match_key_bytes_10_T_1 ? phv_data_15 : _GEN_2115; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2117 = 8'h10 == _match_key_bytes_10_T_1 ? phv_data_16 : _GEN_2116; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2118 = 8'h11 == _match_key_bytes_10_T_1 ? phv_data_17 : _GEN_2117; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2119 = 8'h12 == _match_key_bytes_10_T_1 ? phv_data_18 : _GEN_2118; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2120 = 8'h13 == _match_key_bytes_10_T_1 ? phv_data_19 : _GEN_2119; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2121 = 8'h14 == _match_key_bytes_10_T_1 ? phv_data_20 : _GEN_2120; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2122 = 8'h15 == _match_key_bytes_10_T_1 ? phv_data_21 : _GEN_2121; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2123 = 8'h16 == _match_key_bytes_10_T_1 ? phv_data_22 : _GEN_2122; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2124 = 8'h17 == _match_key_bytes_10_T_1 ? phv_data_23 : _GEN_2123; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2125 = 8'h18 == _match_key_bytes_10_T_1 ? phv_data_24 : _GEN_2124; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2126 = 8'h19 == _match_key_bytes_10_T_1 ? phv_data_25 : _GEN_2125; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2127 = 8'h1a == _match_key_bytes_10_T_1 ? phv_data_26 : _GEN_2126; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2128 = 8'h1b == _match_key_bytes_10_T_1 ? phv_data_27 : _GEN_2127; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2129 = 8'h1c == _match_key_bytes_10_T_1 ? phv_data_28 : _GEN_2128; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2130 = 8'h1d == _match_key_bytes_10_T_1 ? phv_data_29 : _GEN_2129; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2131 = 8'h1e == _match_key_bytes_10_T_1 ? phv_data_30 : _GEN_2130; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2132 = 8'h1f == _match_key_bytes_10_T_1 ? phv_data_31 : _GEN_2131; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2133 = 8'h20 == _match_key_bytes_10_T_1 ? phv_data_32 : _GEN_2132; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2134 = 8'h21 == _match_key_bytes_10_T_1 ? phv_data_33 : _GEN_2133; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2135 = 8'h22 == _match_key_bytes_10_T_1 ? phv_data_34 : _GEN_2134; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2136 = 8'h23 == _match_key_bytes_10_T_1 ? phv_data_35 : _GEN_2135; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2137 = 8'h24 == _match_key_bytes_10_T_1 ? phv_data_36 : _GEN_2136; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2138 = 8'h25 == _match_key_bytes_10_T_1 ? phv_data_37 : _GEN_2137; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2139 = 8'h26 == _match_key_bytes_10_T_1 ? phv_data_38 : _GEN_2138; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2140 = 8'h27 == _match_key_bytes_10_T_1 ? phv_data_39 : _GEN_2139; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2141 = 8'h28 == _match_key_bytes_10_T_1 ? phv_data_40 : _GEN_2140; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2142 = 8'h29 == _match_key_bytes_10_T_1 ? phv_data_41 : _GEN_2141; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2143 = 8'h2a == _match_key_bytes_10_T_1 ? phv_data_42 : _GEN_2142; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2144 = 8'h2b == _match_key_bytes_10_T_1 ? phv_data_43 : _GEN_2143; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2145 = 8'h2c == _match_key_bytes_10_T_1 ? phv_data_44 : _GEN_2144; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2146 = 8'h2d == _match_key_bytes_10_T_1 ? phv_data_45 : _GEN_2145; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2147 = 8'h2e == _match_key_bytes_10_T_1 ? phv_data_46 : _GEN_2146; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2148 = 8'h2f == _match_key_bytes_10_T_1 ? phv_data_47 : _GEN_2147; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2149 = 8'h30 == _match_key_bytes_10_T_1 ? phv_data_48 : _GEN_2148; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2150 = 8'h31 == _match_key_bytes_10_T_1 ? phv_data_49 : _GEN_2149; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2151 = 8'h32 == _match_key_bytes_10_T_1 ? phv_data_50 : _GEN_2150; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2152 = 8'h33 == _match_key_bytes_10_T_1 ? phv_data_51 : _GEN_2151; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2153 = 8'h34 == _match_key_bytes_10_T_1 ? phv_data_52 : _GEN_2152; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2154 = 8'h35 == _match_key_bytes_10_T_1 ? phv_data_53 : _GEN_2153; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2155 = 8'h36 == _match_key_bytes_10_T_1 ? phv_data_54 : _GEN_2154; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2156 = 8'h37 == _match_key_bytes_10_T_1 ? phv_data_55 : _GEN_2155; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2157 = 8'h38 == _match_key_bytes_10_T_1 ? phv_data_56 : _GEN_2156; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2158 = 8'h39 == _match_key_bytes_10_T_1 ? phv_data_57 : _GEN_2157; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2159 = 8'h3a == _match_key_bytes_10_T_1 ? phv_data_58 : _GEN_2158; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2160 = 8'h3b == _match_key_bytes_10_T_1 ? phv_data_59 : _GEN_2159; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2161 = 8'h3c == _match_key_bytes_10_T_1 ? phv_data_60 : _GEN_2160; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2162 = 8'h3d == _match_key_bytes_10_T_1 ? phv_data_61 : _GEN_2161; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2163 = 8'h3e == _match_key_bytes_10_T_1 ? phv_data_62 : _GEN_2162; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2164 = 8'h3f == _match_key_bytes_10_T_1 ? phv_data_63 : _GEN_2163; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2165 = 8'h40 == _match_key_bytes_10_T_1 ? phv_data_64 : _GEN_2164; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2166 = 8'h41 == _match_key_bytes_10_T_1 ? phv_data_65 : _GEN_2165; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2167 = 8'h42 == _match_key_bytes_10_T_1 ? phv_data_66 : _GEN_2166; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2168 = 8'h43 == _match_key_bytes_10_T_1 ? phv_data_67 : _GEN_2167; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2169 = 8'h44 == _match_key_bytes_10_T_1 ? phv_data_68 : _GEN_2168; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2170 = 8'h45 == _match_key_bytes_10_T_1 ? phv_data_69 : _GEN_2169; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2171 = 8'h46 == _match_key_bytes_10_T_1 ? phv_data_70 : _GEN_2170; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2172 = 8'h47 == _match_key_bytes_10_T_1 ? phv_data_71 : _GEN_2171; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2173 = 8'h48 == _match_key_bytes_10_T_1 ? phv_data_72 : _GEN_2172; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2174 = 8'h49 == _match_key_bytes_10_T_1 ? phv_data_73 : _GEN_2173; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2175 = 8'h4a == _match_key_bytes_10_T_1 ? phv_data_74 : _GEN_2174; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2176 = 8'h4b == _match_key_bytes_10_T_1 ? phv_data_75 : _GEN_2175; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2177 = 8'h4c == _match_key_bytes_10_T_1 ? phv_data_76 : _GEN_2176; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2178 = 8'h4d == _match_key_bytes_10_T_1 ? phv_data_77 : _GEN_2177; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2179 = 8'h4e == _match_key_bytes_10_T_1 ? phv_data_78 : _GEN_2178; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2180 = 8'h4f == _match_key_bytes_10_T_1 ? phv_data_79 : _GEN_2179; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2181 = 8'h50 == _match_key_bytes_10_T_1 ? phv_data_80 : _GEN_2180; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2182 = 8'h51 == _match_key_bytes_10_T_1 ? phv_data_81 : _GEN_2181; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2183 = 8'h52 == _match_key_bytes_10_T_1 ? phv_data_82 : _GEN_2182; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2184 = 8'h53 == _match_key_bytes_10_T_1 ? phv_data_83 : _GEN_2183; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2185 = 8'h54 == _match_key_bytes_10_T_1 ? phv_data_84 : _GEN_2184; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2186 = 8'h55 == _match_key_bytes_10_T_1 ? phv_data_85 : _GEN_2185; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2187 = 8'h56 == _match_key_bytes_10_T_1 ? phv_data_86 : _GEN_2186; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2188 = 8'h57 == _match_key_bytes_10_T_1 ? phv_data_87 : _GEN_2187; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2189 = 8'h58 == _match_key_bytes_10_T_1 ? phv_data_88 : _GEN_2188; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2190 = 8'h59 == _match_key_bytes_10_T_1 ? phv_data_89 : _GEN_2189; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2191 = 8'h5a == _match_key_bytes_10_T_1 ? phv_data_90 : _GEN_2190; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2192 = 8'h5b == _match_key_bytes_10_T_1 ? phv_data_91 : _GEN_2191; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2193 = 8'h5c == _match_key_bytes_10_T_1 ? phv_data_92 : _GEN_2192; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2194 = 8'h5d == _match_key_bytes_10_T_1 ? phv_data_93 : _GEN_2193; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2195 = 8'h5e == _match_key_bytes_10_T_1 ? phv_data_94 : _GEN_2194; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2196 = 8'h5f == _match_key_bytes_10_T_1 ? phv_data_95 : _GEN_2195; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2197 = 8'h60 == _match_key_bytes_10_T_1 ? phv_data_96 : _GEN_2196; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2198 = 8'h61 == _match_key_bytes_10_T_1 ? phv_data_97 : _GEN_2197; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2199 = 8'h62 == _match_key_bytes_10_T_1 ? phv_data_98 : _GEN_2198; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2200 = 8'h63 == _match_key_bytes_10_T_1 ? phv_data_99 : _GEN_2199; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2201 = 8'h64 == _match_key_bytes_10_T_1 ? phv_data_100 : _GEN_2200; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2202 = 8'h65 == _match_key_bytes_10_T_1 ? phv_data_101 : _GEN_2201; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2203 = 8'h66 == _match_key_bytes_10_T_1 ? phv_data_102 : _GEN_2202; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2204 = 8'h67 == _match_key_bytes_10_T_1 ? phv_data_103 : _GEN_2203; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2205 = 8'h68 == _match_key_bytes_10_T_1 ? phv_data_104 : _GEN_2204; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2206 = 8'h69 == _match_key_bytes_10_T_1 ? phv_data_105 : _GEN_2205; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2207 = 8'h6a == _match_key_bytes_10_T_1 ? phv_data_106 : _GEN_2206; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2208 = 8'h6b == _match_key_bytes_10_T_1 ? phv_data_107 : _GEN_2207; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2209 = 8'h6c == _match_key_bytes_10_T_1 ? phv_data_108 : _GEN_2208; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2210 = 8'h6d == _match_key_bytes_10_T_1 ? phv_data_109 : _GEN_2209; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2211 = 8'h6e == _match_key_bytes_10_T_1 ? phv_data_110 : _GEN_2210; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2212 = 8'h6f == _match_key_bytes_10_T_1 ? phv_data_111 : _GEN_2211; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2213 = 8'h70 == _match_key_bytes_10_T_1 ? phv_data_112 : _GEN_2212; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2214 = 8'h71 == _match_key_bytes_10_T_1 ? phv_data_113 : _GEN_2213; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2215 = 8'h72 == _match_key_bytes_10_T_1 ? phv_data_114 : _GEN_2214; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2216 = 8'h73 == _match_key_bytes_10_T_1 ? phv_data_115 : _GEN_2215; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2217 = 8'h74 == _match_key_bytes_10_T_1 ? phv_data_116 : _GEN_2216; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2218 = 8'h75 == _match_key_bytes_10_T_1 ? phv_data_117 : _GEN_2217; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2219 = 8'h76 == _match_key_bytes_10_T_1 ? phv_data_118 : _GEN_2218; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2220 = 8'h77 == _match_key_bytes_10_T_1 ? phv_data_119 : _GEN_2219; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2221 = 8'h78 == _match_key_bytes_10_T_1 ? phv_data_120 : _GEN_2220; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2222 = 8'h79 == _match_key_bytes_10_T_1 ? phv_data_121 : _GEN_2221; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2223 = 8'h7a == _match_key_bytes_10_T_1 ? phv_data_122 : _GEN_2222; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2224 = 8'h7b == _match_key_bytes_10_T_1 ? phv_data_123 : _GEN_2223; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2225 = 8'h7c == _match_key_bytes_10_T_1 ? phv_data_124 : _GEN_2224; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2226 = 8'h7d == _match_key_bytes_10_T_1 ? phv_data_125 : _GEN_2225; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2227 = 8'h7e == _match_key_bytes_10_T_1 ? phv_data_126 : _GEN_2226; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2228 = 8'h7f == _match_key_bytes_10_T_1 ? phv_data_127 : _GEN_2227; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2229 = 8'h80 == _match_key_bytes_10_T_1 ? phv_data_128 : _GEN_2228; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2230 = 8'h81 == _match_key_bytes_10_T_1 ? phv_data_129 : _GEN_2229; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2231 = 8'h82 == _match_key_bytes_10_T_1 ? phv_data_130 : _GEN_2230; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2232 = 8'h83 == _match_key_bytes_10_T_1 ? phv_data_131 : _GEN_2231; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2233 = 8'h84 == _match_key_bytes_10_T_1 ? phv_data_132 : _GEN_2232; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2234 = 8'h85 == _match_key_bytes_10_T_1 ? phv_data_133 : _GEN_2233; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2235 = 8'h86 == _match_key_bytes_10_T_1 ? phv_data_134 : _GEN_2234; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2236 = 8'h87 == _match_key_bytes_10_T_1 ? phv_data_135 : _GEN_2235; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2237 = 8'h88 == _match_key_bytes_10_T_1 ? phv_data_136 : _GEN_2236; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2238 = 8'h89 == _match_key_bytes_10_T_1 ? phv_data_137 : _GEN_2237; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2239 = 8'h8a == _match_key_bytes_10_T_1 ? phv_data_138 : _GEN_2238; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2240 = 8'h8b == _match_key_bytes_10_T_1 ? phv_data_139 : _GEN_2239; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2241 = 8'h8c == _match_key_bytes_10_T_1 ? phv_data_140 : _GEN_2240; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2242 = 8'h8d == _match_key_bytes_10_T_1 ? phv_data_141 : _GEN_2241; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2243 = 8'h8e == _match_key_bytes_10_T_1 ? phv_data_142 : _GEN_2242; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2244 = 8'h8f == _match_key_bytes_10_T_1 ? phv_data_143 : _GEN_2243; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2245 = 8'h90 == _match_key_bytes_10_T_1 ? phv_data_144 : _GEN_2244; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2246 = 8'h91 == _match_key_bytes_10_T_1 ? phv_data_145 : _GEN_2245; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2247 = 8'h92 == _match_key_bytes_10_T_1 ? phv_data_146 : _GEN_2246; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2248 = 8'h93 == _match_key_bytes_10_T_1 ? phv_data_147 : _GEN_2247; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2249 = 8'h94 == _match_key_bytes_10_T_1 ? phv_data_148 : _GEN_2248; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2250 = 8'h95 == _match_key_bytes_10_T_1 ? phv_data_149 : _GEN_2249; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2251 = 8'h96 == _match_key_bytes_10_T_1 ? phv_data_150 : _GEN_2250; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2252 = 8'h97 == _match_key_bytes_10_T_1 ? phv_data_151 : _GEN_2251; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2253 = 8'h98 == _match_key_bytes_10_T_1 ? phv_data_152 : _GEN_2252; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2254 = 8'h99 == _match_key_bytes_10_T_1 ? phv_data_153 : _GEN_2253; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2255 = 8'h9a == _match_key_bytes_10_T_1 ? phv_data_154 : _GEN_2254; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2256 = 8'h9b == _match_key_bytes_10_T_1 ? phv_data_155 : _GEN_2255; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2257 = 8'h9c == _match_key_bytes_10_T_1 ? phv_data_156 : _GEN_2256; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2258 = 8'h9d == _match_key_bytes_10_T_1 ? phv_data_157 : _GEN_2257; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2259 = 8'h9e == _match_key_bytes_10_T_1 ? phv_data_158 : _GEN_2258; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2260 = 8'h9f == _match_key_bytes_10_T_1 ? phv_data_159 : _GEN_2259; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_10 = 8'hd < _GEN_6 ? _GEN_2260 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_9_T_1 = key_offset + 8'he; // @[matcher.scala 72:98]
  wire [7:0] _GEN_2263 = 8'h1 == _match_key_bytes_9_T_1 ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2264 = 8'h2 == _match_key_bytes_9_T_1 ? phv_data_2 : _GEN_2263; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2265 = 8'h3 == _match_key_bytes_9_T_1 ? phv_data_3 : _GEN_2264; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2266 = 8'h4 == _match_key_bytes_9_T_1 ? phv_data_4 : _GEN_2265; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2267 = 8'h5 == _match_key_bytes_9_T_1 ? phv_data_5 : _GEN_2266; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2268 = 8'h6 == _match_key_bytes_9_T_1 ? phv_data_6 : _GEN_2267; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2269 = 8'h7 == _match_key_bytes_9_T_1 ? phv_data_7 : _GEN_2268; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2270 = 8'h8 == _match_key_bytes_9_T_1 ? phv_data_8 : _GEN_2269; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2271 = 8'h9 == _match_key_bytes_9_T_1 ? phv_data_9 : _GEN_2270; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2272 = 8'ha == _match_key_bytes_9_T_1 ? phv_data_10 : _GEN_2271; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2273 = 8'hb == _match_key_bytes_9_T_1 ? phv_data_11 : _GEN_2272; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2274 = 8'hc == _match_key_bytes_9_T_1 ? phv_data_12 : _GEN_2273; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2275 = 8'hd == _match_key_bytes_9_T_1 ? phv_data_13 : _GEN_2274; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2276 = 8'he == _match_key_bytes_9_T_1 ? phv_data_14 : _GEN_2275; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2277 = 8'hf == _match_key_bytes_9_T_1 ? phv_data_15 : _GEN_2276; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2278 = 8'h10 == _match_key_bytes_9_T_1 ? phv_data_16 : _GEN_2277; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2279 = 8'h11 == _match_key_bytes_9_T_1 ? phv_data_17 : _GEN_2278; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2280 = 8'h12 == _match_key_bytes_9_T_1 ? phv_data_18 : _GEN_2279; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2281 = 8'h13 == _match_key_bytes_9_T_1 ? phv_data_19 : _GEN_2280; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2282 = 8'h14 == _match_key_bytes_9_T_1 ? phv_data_20 : _GEN_2281; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2283 = 8'h15 == _match_key_bytes_9_T_1 ? phv_data_21 : _GEN_2282; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2284 = 8'h16 == _match_key_bytes_9_T_1 ? phv_data_22 : _GEN_2283; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2285 = 8'h17 == _match_key_bytes_9_T_1 ? phv_data_23 : _GEN_2284; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2286 = 8'h18 == _match_key_bytes_9_T_1 ? phv_data_24 : _GEN_2285; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2287 = 8'h19 == _match_key_bytes_9_T_1 ? phv_data_25 : _GEN_2286; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2288 = 8'h1a == _match_key_bytes_9_T_1 ? phv_data_26 : _GEN_2287; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2289 = 8'h1b == _match_key_bytes_9_T_1 ? phv_data_27 : _GEN_2288; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2290 = 8'h1c == _match_key_bytes_9_T_1 ? phv_data_28 : _GEN_2289; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2291 = 8'h1d == _match_key_bytes_9_T_1 ? phv_data_29 : _GEN_2290; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2292 = 8'h1e == _match_key_bytes_9_T_1 ? phv_data_30 : _GEN_2291; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2293 = 8'h1f == _match_key_bytes_9_T_1 ? phv_data_31 : _GEN_2292; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2294 = 8'h20 == _match_key_bytes_9_T_1 ? phv_data_32 : _GEN_2293; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2295 = 8'h21 == _match_key_bytes_9_T_1 ? phv_data_33 : _GEN_2294; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2296 = 8'h22 == _match_key_bytes_9_T_1 ? phv_data_34 : _GEN_2295; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2297 = 8'h23 == _match_key_bytes_9_T_1 ? phv_data_35 : _GEN_2296; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2298 = 8'h24 == _match_key_bytes_9_T_1 ? phv_data_36 : _GEN_2297; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2299 = 8'h25 == _match_key_bytes_9_T_1 ? phv_data_37 : _GEN_2298; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2300 = 8'h26 == _match_key_bytes_9_T_1 ? phv_data_38 : _GEN_2299; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2301 = 8'h27 == _match_key_bytes_9_T_1 ? phv_data_39 : _GEN_2300; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2302 = 8'h28 == _match_key_bytes_9_T_1 ? phv_data_40 : _GEN_2301; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2303 = 8'h29 == _match_key_bytes_9_T_1 ? phv_data_41 : _GEN_2302; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2304 = 8'h2a == _match_key_bytes_9_T_1 ? phv_data_42 : _GEN_2303; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2305 = 8'h2b == _match_key_bytes_9_T_1 ? phv_data_43 : _GEN_2304; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2306 = 8'h2c == _match_key_bytes_9_T_1 ? phv_data_44 : _GEN_2305; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2307 = 8'h2d == _match_key_bytes_9_T_1 ? phv_data_45 : _GEN_2306; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2308 = 8'h2e == _match_key_bytes_9_T_1 ? phv_data_46 : _GEN_2307; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2309 = 8'h2f == _match_key_bytes_9_T_1 ? phv_data_47 : _GEN_2308; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2310 = 8'h30 == _match_key_bytes_9_T_1 ? phv_data_48 : _GEN_2309; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2311 = 8'h31 == _match_key_bytes_9_T_1 ? phv_data_49 : _GEN_2310; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2312 = 8'h32 == _match_key_bytes_9_T_1 ? phv_data_50 : _GEN_2311; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2313 = 8'h33 == _match_key_bytes_9_T_1 ? phv_data_51 : _GEN_2312; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2314 = 8'h34 == _match_key_bytes_9_T_1 ? phv_data_52 : _GEN_2313; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2315 = 8'h35 == _match_key_bytes_9_T_1 ? phv_data_53 : _GEN_2314; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2316 = 8'h36 == _match_key_bytes_9_T_1 ? phv_data_54 : _GEN_2315; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2317 = 8'h37 == _match_key_bytes_9_T_1 ? phv_data_55 : _GEN_2316; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2318 = 8'h38 == _match_key_bytes_9_T_1 ? phv_data_56 : _GEN_2317; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2319 = 8'h39 == _match_key_bytes_9_T_1 ? phv_data_57 : _GEN_2318; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2320 = 8'h3a == _match_key_bytes_9_T_1 ? phv_data_58 : _GEN_2319; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2321 = 8'h3b == _match_key_bytes_9_T_1 ? phv_data_59 : _GEN_2320; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2322 = 8'h3c == _match_key_bytes_9_T_1 ? phv_data_60 : _GEN_2321; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2323 = 8'h3d == _match_key_bytes_9_T_1 ? phv_data_61 : _GEN_2322; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2324 = 8'h3e == _match_key_bytes_9_T_1 ? phv_data_62 : _GEN_2323; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2325 = 8'h3f == _match_key_bytes_9_T_1 ? phv_data_63 : _GEN_2324; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2326 = 8'h40 == _match_key_bytes_9_T_1 ? phv_data_64 : _GEN_2325; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2327 = 8'h41 == _match_key_bytes_9_T_1 ? phv_data_65 : _GEN_2326; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2328 = 8'h42 == _match_key_bytes_9_T_1 ? phv_data_66 : _GEN_2327; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2329 = 8'h43 == _match_key_bytes_9_T_1 ? phv_data_67 : _GEN_2328; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2330 = 8'h44 == _match_key_bytes_9_T_1 ? phv_data_68 : _GEN_2329; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2331 = 8'h45 == _match_key_bytes_9_T_1 ? phv_data_69 : _GEN_2330; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2332 = 8'h46 == _match_key_bytes_9_T_1 ? phv_data_70 : _GEN_2331; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2333 = 8'h47 == _match_key_bytes_9_T_1 ? phv_data_71 : _GEN_2332; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2334 = 8'h48 == _match_key_bytes_9_T_1 ? phv_data_72 : _GEN_2333; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2335 = 8'h49 == _match_key_bytes_9_T_1 ? phv_data_73 : _GEN_2334; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2336 = 8'h4a == _match_key_bytes_9_T_1 ? phv_data_74 : _GEN_2335; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2337 = 8'h4b == _match_key_bytes_9_T_1 ? phv_data_75 : _GEN_2336; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2338 = 8'h4c == _match_key_bytes_9_T_1 ? phv_data_76 : _GEN_2337; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2339 = 8'h4d == _match_key_bytes_9_T_1 ? phv_data_77 : _GEN_2338; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2340 = 8'h4e == _match_key_bytes_9_T_1 ? phv_data_78 : _GEN_2339; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2341 = 8'h4f == _match_key_bytes_9_T_1 ? phv_data_79 : _GEN_2340; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2342 = 8'h50 == _match_key_bytes_9_T_1 ? phv_data_80 : _GEN_2341; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2343 = 8'h51 == _match_key_bytes_9_T_1 ? phv_data_81 : _GEN_2342; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2344 = 8'h52 == _match_key_bytes_9_T_1 ? phv_data_82 : _GEN_2343; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2345 = 8'h53 == _match_key_bytes_9_T_1 ? phv_data_83 : _GEN_2344; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2346 = 8'h54 == _match_key_bytes_9_T_1 ? phv_data_84 : _GEN_2345; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2347 = 8'h55 == _match_key_bytes_9_T_1 ? phv_data_85 : _GEN_2346; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2348 = 8'h56 == _match_key_bytes_9_T_1 ? phv_data_86 : _GEN_2347; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2349 = 8'h57 == _match_key_bytes_9_T_1 ? phv_data_87 : _GEN_2348; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2350 = 8'h58 == _match_key_bytes_9_T_1 ? phv_data_88 : _GEN_2349; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2351 = 8'h59 == _match_key_bytes_9_T_1 ? phv_data_89 : _GEN_2350; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2352 = 8'h5a == _match_key_bytes_9_T_1 ? phv_data_90 : _GEN_2351; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2353 = 8'h5b == _match_key_bytes_9_T_1 ? phv_data_91 : _GEN_2352; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2354 = 8'h5c == _match_key_bytes_9_T_1 ? phv_data_92 : _GEN_2353; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2355 = 8'h5d == _match_key_bytes_9_T_1 ? phv_data_93 : _GEN_2354; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2356 = 8'h5e == _match_key_bytes_9_T_1 ? phv_data_94 : _GEN_2355; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2357 = 8'h5f == _match_key_bytes_9_T_1 ? phv_data_95 : _GEN_2356; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2358 = 8'h60 == _match_key_bytes_9_T_1 ? phv_data_96 : _GEN_2357; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2359 = 8'h61 == _match_key_bytes_9_T_1 ? phv_data_97 : _GEN_2358; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2360 = 8'h62 == _match_key_bytes_9_T_1 ? phv_data_98 : _GEN_2359; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2361 = 8'h63 == _match_key_bytes_9_T_1 ? phv_data_99 : _GEN_2360; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2362 = 8'h64 == _match_key_bytes_9_T_1 ? phv_data_100 : _GEN_2361; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2363 = 8'h65 == _match_key_bytes_9_T_1 ? phv_data_101 : _GEN_2362; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2364 = 8'h66 == _match_key_bytes_9_T_1 ? phv_data_102 : _GEN_2363; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2365 = 8'h67 == _match_key_bytes_9_T_1 ? phv_data_103 : _GEN_2364; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2366 = 8'h68 == _match_key_bytes_9_T_1 ? phv_data_104 : _GEN_2365; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2367 = 8'h69 == _match_key_bytes_9_T_1 ? phv_data_105 : _GEN_2366; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2368 = 8'h6a == _match_key_bytes_9_T_1 ? phv_data_106 : _GEN_2367; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2369 = 8'h6b == _match_key_bytes_9_T_1 ? phv_data_107 : _GEN_2368; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2370 = 8'h6c == _match_key_bytes_9_T_1 ? phv_data_108 : _GEN_2369; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2371 = 8'h6d == _match_key_bytes_9_T_1 ? phv_data_109 : _GEN_2370; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2372 = 8'h6e == _match_key_bytes_9_T_1 ? phv_data_110 : _GEN_2371; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2373 = 8'h6f == _match_key_bytes_9_T_1 ? phv_data_111 : _GEN_2372; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2374 = 8'h70 == _match_key_bytes_9_T_1 ? phv_data_112 : _GEN_2373; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2375 = 8'h71 == _match_key_bytes_9_T_1 ? phv_data_113 : _GEN_2374; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2376 = 8'h72 == _match_key_bytes_9_T_1 ? phv_data_114 : _GEN_2375; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2377 = 8'h73 == _match_key_bytes_9_T_1 ? phv_data_115 : _GEN_2376; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2378 = 8'h74 == _match_key_bytes_9_T_1 ? phv_data_116 : _GEN_2377; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2379 = 8'h75 == _match_key_bytes_9_T_1 ? phv_data_117 : _GEN_2378; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2380 = 8'h76 == _match_key_bytes_9_T_1 ? phv_data_118 : _GEN_2379; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2381 = 8'h77 == _match_key_bytes_9_T_1 ? phv_data_119 : _GEN_2380; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2382 = 8'h78 == _match_key_bytes_9_T_1 ? phv_data_120 : _GEN_2381; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2383 = 8'h79 == _match_key_bytes_9_T_1 ? phv_data_121 : _GEN_2382; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2384 = 8'h7a == _match_key_bytes_9_T_1 ? phv_data_122 : _GEN_2383; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2385 = 8'h7b == _match_key_bytes_9_T_1 ? phv_data_123 : _GEN_2384; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2386 = 8'h7c == _match_key_bytes_9_T_1 ? phv_data_124 : _GEN_2385; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2387 = 8'h7d == _match_key_bytes_9_T_1 ? phv_data_125 : _GEN_2386; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2388 = 8'h7e == _match_key_bytes_9_T_1 ? phv_data_126 : _GEN_2387; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2389 = 8'h7f == _match_key_bytes_9_T_1 ? phv_data_127 : _GEN_2388; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2390 = 8'h80 == _match_key_bytes_9_T_1 ? phv_data_128 : _GEN_2389; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2391 = 8'h81 == _match_key_bytes_9_T_1 ? phv_data_129 : _GEN_2390; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2392 = 8'h82 == _match_key_bytes_9_T_1 ? phv_data_130 : _GEN_2391; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2393 = 8'h83 == _match_key_bytes_9_T_1 ? phv_data_131 : _GEN_2392; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2394 = 8'h84 == _match_key_bytes_9_T_1 ? phv_data_132 : _GEN_2393; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2395 = 8'h85 == _match_key_bytes_9_T_1 ? phv_data_133 : _GEN_2394; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2396 = 8'h86 == _match_key_bytes_9_T_1 ? phv_data_134 : _GEN_2395; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2397 = 8'h87 == _match_key_bytes_9_T_1 ? phv_data_135 : _GEN_2396; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2398 = 8'h88 == _match_key_bytes_9_T_1 ? phv_data_136 : _GEN_2397; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2399 = 8'h89 == _match_key_bytes_9_T_1 ? phv_data_137 : _GEN_2398; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2400 = 8'h8a == _match_key_bytes_9_T_1 ? phv_data_138 : _GEN_2399; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2401 = 8'h8b == _match_key_bytes_9_T_1 ? phv_data_139 : _GEN_2400; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2402 = 8'h8c == _match_key_bytes_9_T_1 ? phv_data_140 : _GEN_2401; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2403 = 8'h8d == _match_key_bytes_9_T_1 ? phv_data_141 : _GEN_2402; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2404 = 8'h8e == _match_key_bytes_9_T_1 ? phv_data_142 : _GEN_2403; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2405 = 8'h8f == _match_key_bytes_9_T_1 ? phv_data_143 : _GEN_2404; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2406 = 8'h90 == _match_key_bytes_9_T_1 ? phv_data_144 : _GEN_2405; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2407 = 8'h91 == _match_key_bytes_9_T_1 ? phv_data_145 : _GEN_2406; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2408 = 8'h92 == _match_key_bytes_9_T_1 ? phv_data_146 : _GEN_2407; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2409 = 8'h93 == _match_key_bytes_9_T_1 ? phv_data_147 : _GEN_2408; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2410 = 8'h94 == _match_key_bytes_9_T_1 ? phv_data_148 : _GEN_2409; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2411 = 8'h95 == _match_key_bytes_9_T_1 ? phv_data_149 : _GEN_2410; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2412 = 8'h96 == _match_key_bytes_9_T_1 ? phv_data_150 : _GEN_2411; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2413 = 8'h97 == _match_key_bytes_9_T_1 ? phv_data_151 : _GEN_2412; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2414 = 8'h98 == _match_key_bytes_9_T_1 ? phv_data_152 : _GEN_2413; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2415 = 8'h99 == _match_key_bytes_9_T_1 ? phv_data_153 : _GEN_2414; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2416 = 8'h9a == _match_key_bytes_9_T_1 ? phv_data_154 : _GEN_2415; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2417 = 8'h9b == _match_key_bytes_9_T_1 ? phv_data_155 : _GEN_2416; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2418 = 8'h9c == _match_key_bytes_9_T_1 ? phv_data_156 : _GEN_2417; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2419 = 8'h9d == _match_key_bytes_9_T_1 ? phv_data_157 : _GEN_2418; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2420 = 8'h9e == _match_key_bytes_9_T_1 ? phv_data_158 : _GEN_2419; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2421 = 8'h9f == _match_key_bytes_9_T_1 ? phv_data_159 : _GEN_2420; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_9 = 8'he < _GEN_6 ? _GEN_2421 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_8_T_1 = key_offset + 8'hf; // @[matcher.scala 72:98]
  wire [7:0] _GEN_2424 = 8'h1 == _match_key_bytes_8_T_1 ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2425 = 8'h2 == _match_key_bytes_8_T_1 ? phv_data_2 : _GEN_2424; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2426 = 8'h3 == _match_key_bytes_8_T_1 ? phv_data_3 : _GEN_2425; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2427 = 8'h4 == _match_key_bytes_8_T_1 ? phv_data_4 : _GEN_2426; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2428 = 8'h5 == _match_key_bytes_8_T_1 ? phv_data_5 : _GEN_2427; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2429 = 8'h6 == _match_key_bytes_8_T_1 ? phv_data_6 : _GEN_2428; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2430 = 8'h7 == _match_key_bytes_8_T_1 ? phv_data_7 : _GEN_2429; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2431 = 8'h8 == _match_key_bytes_8_T_1 ? phv_data_8 : _GEN_2430; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2432 = 8'h9 == _match_key_bytes_8_T_1 ? phv_data_9 : _GEN_2431; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2433 = 8'ha == _match_key_bytes_8_T_1 ? phv_data_10 : _GEN_2432; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2434 = 8'hb == _match_key_bytes_8_T_1 ? phv_data_11 : _GEN_2433; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2435 = 8'hc == _match_key_bytes_8_T_1 ? phv_data_12 : _GEN_2434; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2436 = 8'hd == _match_key_bytes_8_T_1 ? phv_data_13 : _GEN_2435; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2437 = 8'he == _match_key_bytes_8_T_1 ? phv_data_14 : _GEN_2436; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2438 = 8'hf == _match_key_bytes_8_T_1 ? phv_data_15 : _GEN_2437; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2439 = 8'h10 == _match_key_bytes_8_T_1 ? phv_data_16 : _GEN_2438; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2440 = 8'h11 == _match_key_bytes_8_T_1 ? phv_data_17 : _GEN_2439; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2441 = 8'h12 == _match_key_bytes_8_T_1 ? phv_data_18 : _GEN_2440; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2442 = 8'h13 == _match_key_bytes_8_T_1 ? phv_data_19 : _GEN_2441; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2443 = 8'h14 == _match_key_bytes_8_T_1 ? phv_data_20 : _GEN_2442; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2444 = 8'h15 == _match_key_bytes_8_T_1 ? phv_data_21 : _GEN_2443; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2445 = 8'h16 == _match_key_bytes_8_T_1 ? phv_data_22 : _GEN_2444; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2446 = 8'h17 == _match_key_bytes_8_T_1 ? phv_data_23 : _GEN_2445; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2447 = 8'h18 == _match_key_bytes_8_T_1 ? phv_data_24 : _GEN_2446; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2448 = 8'h19 == _match_key_bytes_8_T_1 ? phv_data_25 : _GEN_2447; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2449 = 8'h1a == _match_key_bytes_8_T_1 ? phv_data_26 : _GEN_2448; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2450 = 8'h1b == _match_key_bytes_8_T_1 ? phv_data_27 : _GEN_2449; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2451 = 8'h1c == _match_key_bytes_8_T_1 ? phv_data_28 : _GEN_2450; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2452 = 8'h1d == _match_key_bytes_8_T_1 ? phv_data_29 : _GEN_2451; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2453 = 8'h1e == _match_key_bytes_8_T_1 ? phv_data_30 : _GEN_2452; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2454 = 8'h1f == _match_key_bytes_8_T_1 ? phv_data_31 : _GEN_2453; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2455 = 8'h20 == _match_key_bytes_8_T_1 ? phv_data_32 : _GEN_2454; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2456 = 8'h21 == _match_key_bytes_8_T_1 ? phv_data_33 : _GEN_2455; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2457 = 8'h22 == _match_key_bytes_8_T_1 ? phv_data_34 : _GEN_2456; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2458 = 8'h23 == _match_key_bytes_8_T_1 ? phv_data_35 : _GEN_2457; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2459 = 8'h24 == _match_key_bytes_8_T_1 ? phv_data_36 : _GEN_2458; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2460 = 8'h25 == _match_key_bytes_8_T_1 ? phv_data_37 : _GEN_2459; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2461 = 8'h26 == _match_key_bytes_8_T_1 ? phv_data_38 : _GEN_2460; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2462 = 8'h27 == _match_key_bytes_8_T_1 ? phv_data_39 : _GEN_2461; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2463 = 8'h28 == _match_key_bytes_8_T_1 ? phv_data_40 : _GEN_2462; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2464 = 8'h29 == _match_key_bytes_8_T_1 ? phv_data_41 : _GEN_2463; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2465 = 8'h2a == _match_key_bytes_8_T_1 ? phv_data_42 : _GEN_2464; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2466 = 8'h2b == _match_key_bytes_8_T_1 ? phv_data_43 : _GEN_2465; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2467 = 8'h2c == _match_key_bytes_8_T_1 ? phv_data_44 : _GEN_2466; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2468 = 8'h2d == _match_key_bytes_8_T_1 ? phv_data_45 : _GEN_2467; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2469 = 8'h2e == _match_key_bytes_8_T_1 ? phv_data_46 : _GEN_2468; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2470 = 8'h2f == _match_key_bytes_8_T_1 ? phv_data_47 : _GEN_2469; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2471 = 8'h30 == _match_key_bytes_8_T_1 ? phv_data_48 : _GEN_2470; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2472 = 8'h31 == _match_key_bytes_8_T_1 ? phv_data_49 : _GEN_2471; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2473 = 8'h32 == _match_key_bytes_8_T_1 ? phv_data_50 : _GEN_2472; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2474 = 8'h33 == _match_key_bytes_8_T_1 ? phv_data_51 : _GEN_2473; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2475 = 8'h34 == _match_key_bytes_8_T_1 ? phv_data_52 : _GEN_2474; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2476 = 8'h35 == _match_key_bytes_8_T_1 ? phv_data_53 : _GEN_2475; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2477 = 8'h36 == _match_key_bytes_8_T_1 ? phv_data_54 : _GEN_2476; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2478 = 8'h37 == _match_key_bytes_8_T_1 ? phv_data_55 : _GEN_2477; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2479 = 8'h38 == _match_key_bytes_8_T_1 ? phv_data_56 : _GEN_2478; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2480 = 8'h39 == _match_key_bytes_8_T_1 ? phv_data_57 : _GEN_2479; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2481 = 8'h3a == _match_key_bytes_8_T_1 ? phv_data_58 : _GEN_2480; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2482 = 8'h3b == _match_key_bytes_8_T_1 ? phv_data_59 : _GEN_2481; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2483 = 8'h3c == _match_key_bytes_8_T_1 ? phv_data_60 : _GEN_2482; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2484 = 8'h3d == _match_key_bytes_8_T_1 ? phv_data_61 : _GEN_2483; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2485 = 8'h3e == _match_key_bytes_8_T_1 ? phv_data_62 : _GEN_2484; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2486 = 8'h3f == _match_key_bytes_8_T_1 ? phv_data_63 : _GEN_2485; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2487 = 8'h40 == _match_key_bytes_8_T_1 ? phv_data_64 : _GEN_2486; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2488 = 8'h41 == _match_key_bytes_8_T_1 ? phv_data_65 : _GEN_2487; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2489 = 8'h42 == _match_key_bytes_8_T_1 ? phv_data_66 : _GEN_2488; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2490 = 8'h43 == _match_key_bytes_8_T_1 ? phv_data_67 : _GEN_2489; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2491 = 8'h44 == _match_key_bytes_8_T_1 ? phv_data_68 : _GEN_2490; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2492 = 8'h45 == _match_key_bytes_8_T_1 ? phv_data_69 : _GEN_2491; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2493 = 8'h46 == _match_key_bytes_8_T_1 ? phv_data_70 : _GEN_2492; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2494 = 8'h47 == _match_key_bytes_8_T_1 ? phv_data_71 : _GEN_2493; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2495 = 8'h48 == _match_key_bytes_8_T_1 ? phv_data_72 : _GEN_2494; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2496 = 8'h49 == _match_key_bytes_8_T_1 ? phv_data_73 : _GEN_2495; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2497 = 8'h4a == _match_key_bytes_8_T_1 ? phv_data_74 : _GEN_2496; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2498 = 8'h4b == _match_key_bytes_8_T_1 ? phv_data_75 : _GEN_2497; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2499 = 8'h4c == _match_key_bytes_8_T_1 ? phv_data_76 : _GEN_2498; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2500 = 8'h4d == _match_key_bytes_8_T_1 ? phv_data_77 : _GEN_2499; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2501 = 8'h4e == _match_key_bytes_8_T_1 ? phv_data_78 : _GEN_2500; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2502 = 8'h4f == _match_key_bytes_8_T_1 ? phv_data_79 : _GEN_2501; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2503 = 8'h50 == _match_key_bytes_8_T_1 ? phv_data_80 : _GEN_2502; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2504 = 8'h51 == _match_key_bytes_8_T_1 ? phv_data_81 : _GEN_2503; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2505 = 8'h52 == _match_key_bytes_8_T_1 ? phv_data_82 : _GEN_2504; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2506 = 8'h53 == _match_key_bytes_8_T_1 ? phv_data_83 : _GEN_2505; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2507 = 8'h54 == _match_key_bytes_8_T_1 ? phv_data_84 : _GEN_2506; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2508 = 8'h55 == _match_key_bytes_8_T_1 ? phv_data_85 : _GEN_2507; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2509 = 8'h56 == _match_key_bytes_8_T_1 ? phv_data_86 : _GEN_2508; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2510 = 8'h57 == _match_key_bytes_8_T_1 ? phv_data_87 : _GEN_2509; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2511 = 8'h58 == _match_key_bytes_8_T_1 ? phv_data_88 : _GEN_2510; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2512 = 8'h59 == _match_key_bytes_8_T_1 ? phv_data_89 : _GEN_2511; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2513 = 8'h5a == _match_key_bytes_8_T_1 ? phv_data_90 : _GEN_2512; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2514 = 8'h5b == _match_key_bytes_8_T_1 ? phv_data_91 : _GEN_2513; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2515 = 8'h5c == _match_key_bytes_8_T_1 ? phv_data_92 : _GEN_2514; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2516 = 8'h5d == _match_key_bytes_8_T_1 ? phv_data_93 : _GEN_2515; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2517 = 8'h5e == _match_key_bytes_8_T_1 ? phv_data_94 : _GEN_2516; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2518 = 8'h5f == _match_key_bytes_8_T_1 ? phv_data_95 : _GEN_2517; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2519 = 8'h60 == _match_key_bytes_8_T_1 ? phv_data_96 : _GEN_2518; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2520 = 8'h61 == _match_key_bytes_8_T_1 ? phv_data_97 : _GEN_2519; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2521 = 8'h62 == _match_key_bytes_8_T_1 ? phv_data_98 : _GEN_2520; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2522 = 8'h63 == _match_key_bytes_8_T_1 ? phv_data_99 : _GEN_2521; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2523 = 8'h64 == _match_key_bytes_8_T_1 ? phv_data_100 : _GEN_2522; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2524 = 8'h65 == _match_key_bytes_8_T_1 ? phv_data_101 : _GEN_2523; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2525 = 8'h66 == _match_key_bytes_8_T_1 ? phv_data_102 : _GEN_2524; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2526 = 8'h67 == _match_key_bytes_8_T_1 ? phv_data_103 : _GEN_2525; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2527 = 8'h68 == _match_key_bytes_8_T_1 ? phv_data_104 : _GEN_2526; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2528 = 8'h69 == _match_key_bytes_8_T_1 ? phv_data_105 : _GEN_2527; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2529 = 8'h6a == _match_key_bytes_8_T_1 ? phv_data_106 : _GEN_2528; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2530 = 8'h6b == _match_key_bytes_8_T_1 ? phv_data_107 : _GEN_2529; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2531 = 8'h6c == _match_key_bytes_8_T_1 ? phv_data_108 : _GEN_2530; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2532 = 8'h6d == _match_key_bytes_8_T_1 ? phv_data_109 : _GEN_2531; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2533 = 8'h6e == _match_key_bytes_8_T_1 ? phv_data_110 : _GEN_2532; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2534 = 8'h6f == _match_key_bytes_8_T_1 ? phv_data_111 : _GEN_2533; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2535 = 8'h70 == _match_key_bytes_8_T_1 ? phv_data_112 : _GEN_2534; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2536 = 8'h71 == _match_key_bytes_8_T_1 ? phv_data_113 : _GEN_2535; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2537 = 8'h72 == _match_key_bytes_8_T_1 ? phv_data_114 : _GEN_2536; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2538 = 8'h73 == _match_key_bytes_8_T_1 ? phv_data_115 : _GEN_2537; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2539 = 8'h74 == _match_key_bytes_8_T_1 ? phv_data_116 : _GEN_2538; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2540 = 8'h75 == _match_key_bytes_8_T_1 ? phv_data_117 : _GEN_2539; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2541 = 8'h76 == _match_key_bytes_8_T_1 ? phv_data_118 : _GEN_2540; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2542 = 8'h77 == _match_key_bytes_8_T_1 ? phv_data_119 : _GEN_2541; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2543 = 8'h78 == _match_key_bytes_8_T_1 ? phv_data_120 : _GEN_2542; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2544 = 8'h79 == _match_key_bytes_8_T_1 ? phv_data_121 : _GEN_2543; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2545 = 8'h7a == _match_key_bytes_8_T_1 ? phv_data_122 : _GEN_2544; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2546 = 8'h7b == _match_key_bytes_8_T_1 ? phv_data_123 : _GEN_2545; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2547 = 8'h7c == _match_key_bytes_8_T_1 ? phv_data_124 : _GEN_2546; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2548 = 8'h7d == _match_key_bytes_8_T_1 ? phv_data_125 : _GEN_2547; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2549 = 8'h7e == _match_key_bytes_8_T_1 ? phv_data_126 : _GEN_2548; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2550 = 8'h7f == _match_key_bytes_8_T_1 ? phv_data_127 : _GEN_2549; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2551 = 8'h80 == _match_key_bytes_8_T_1 ? phv_data_128 : _GEN_2550; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2552 = 8'h81 == _match_key_bytes_8_T_1 ? phv_data_129 : _GEN_2551; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2553 = 8'h82 == _match_key_bytes_8_T_1 ? phv_data_130 : _GEN_2552; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2554 = 8'h83 == _match_key_bytes_8_T_1 ? phv_data_131 : _GEN_2553; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2555 = 8'h84 == _match_key_bytes_8_T_1 ? phv_data_132 : _GEN_2554; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2556 = 8'h85 == _match_key_bytes_8_T_1 ? phv_data_133 : _GEN_2555; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2557 = 8'h86 == _match_key_bytes_8_T_1 ? phv_data_134 : _GEN_2556; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2558 = 8'h87 == _match_key_bytes_8_T_1 ? phv_data_135 : _GEN_2557; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2559 = 8'h88 == _match_key_bytes_8_T_1 ? phv_data_136 : _GEN_2558; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2560 = 8'h89 == _match_key_bytes_8_T_1 ? phv_data_137 : _GEN_2559; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2561 = 8'h8a == _match_key_bytes_8_T_1 ? phv_data_138 : _GEN_2560; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2562 = 8'h8b == _match_key_bytes_8_T_1 ? phv_data_139 : _GEN_2561; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2563 = 8'h8c == _match_key_bytes_8_T_1 ? phv_data_140 : _GEN_2562; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2564 = 8'h8d == _match_key_bytes_8_T_1 ? phv_data_141 : _GEN_2563; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2565 = 8'h8e == _match_key_bytes_8_T_1 ? phv_data_142 : _GEN_2564; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2566 = 8'h8f == _match_key_bytes_8_T_1 ? phv_data_143 : _GEN_2565; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2567 = 8'h90 == _match_key_bytes_8_T_1 ? phv_data_144 : _GEN_2566; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2568 = 8'h91 == _match_key_bytes_8_T_1 ? phv_data_145 : _GEN_2567; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2569 = 8'h92 == _match_key_bytes_8_T_1 ? phv_data_146 : _GEN_2568; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2570 = 8'h93 == _match_key_bytes_8_T_1 ? phv_data_147 : _GEN_2569; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2571 = 8'h94 == _match_key_bytes_8_T_1 ? phv_data_148 : _GEN_2570; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2572 = 8'h95 == _match_key_bytes_8_T_1 ? phv_data_149 : _GEN_2571; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2573 = 8'h96 == _match_key_bytes_8_T_1 ? phv_data_150 : _GEN_2572; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2574 = 8'h97 == _match_key_bytes_8_T_1 ? phv_data_151 : _GEN_2573; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2575 = 8'h98 == _match_key_bytes_8_T_1 ? phv_data_152 : _GEN_2574; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2576 = 8'h99 == _match_key_bytes_8_T_1 ? phv_data_153 : _GEN_2575; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2577 = 8'h9a == _match_key_bytes_8_T_1 ? phv_data_154 : _GEN_2576; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2578 = 8'h9b == _match_key_bytes_8_T_1 ? phv_data_155 : _GEN_2577; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2579 = 8'h9c == _match_key_bytes_8_T_1 ? phv_data_156 : _GEN_2578; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2580 = 8'h9d == _match_key_bytes_8_T_1 ? phv_data_157 : _GEN_2579; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2581 = 8'h9e == _match_key_bytes_8_T_1 ? phv_data_158 : _GEN_2580; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2582 = 8'h9f == _match_key_bytes_8_T_1 ? phv_data_159 : _GEN_2581; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_8 = 8'hf < _GEN_6 ? _GEN_2582 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_7_T_1 = key_offset + 8'h10; // @[matcher.scala 72:98]
  wire [7:0] _GEN_2585 = 8'h1 == _match_key_bytes_7_T_1 ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2586 = 8'h2 == _match_key_bytes_7_T_1 ? phv_data_2 : _GEN_2585; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2587 = 8'h3 == _match_key_bytes_7_T_1 ? phv_data_3 : _GEN_2586; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2588 = 8'h4 == _match_key_bytes_7_T_1 ? phv_data_4 : _GEN_2587; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2589 = 8'h5 == _match_key_bytes_7_T_1 ? phv_data_5 : _GEN_2588; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2590 = 8'h6 == _match_key_bytes_7_T_1 ? phv_data_6 : _GEN_2589; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2591 = 8'h7 == _match_key_bytes_7_T_1 ? phv_data_7 : _GEN_2590; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2592 = 8'h8 == _match_key_bytes_7_T_1 ? phv_data_8 : _GEN_2591; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2593 = 8'h9 == _match_key_bytes_7_T_1 ? phv_data_9 : _GEN_2592; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2594 = 8'ha == _match_key_bytes_7_T_1 ? phv_data_10 : _GEN_2593; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2595 = 8'hb == _match_key_bytes_7_T_1 ? phv_data_11 : _GEN_2594; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2596 = 8'hc == _match_key_bytes_7_T_1 ? phv_data_12 : _GEN_2595; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2597 = 8'hd == _match_key_bytes_7_T_1 ? phv_data_13 : _GEN_2596; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2598 = 8'he == _match_key_bytes_7_T_1 ? phv_data_14 : _GEN_2597; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2599 = 8'hf == _match_key_bytes_7_T_1 ? phv_data_15 : _GEN_2598; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2600 = 8'h10 == _match_key_bytes_7_T_1 ? phv_data_16 : _GEN_2599; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2601 = 8'h11 == _match_key_bytes_7_T_1 ? phv_data_17 : _GEN_2600; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2602 = 8'h12 == _match_key_bytes_7_T_1 ? phv_data_18 : _GEN_2601; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2603 = 8'h13 == _match_key_bytes_7_T_1 ? phv_data_19 : _GEN_2602; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2604 = 8'h14 == _match_key_bytes_7_T_1 ? phv_data_20 : _GEN_2603; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2605 = 8'h15 == _match_key_bytes_7_T_1 ? phv_data_21 : _GEN_2604; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2606 = 8'h16 == _match_key_bytes_7_T_1 ? phv_data_22 : _GEN_2605; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2607 = 8'h17 == _match_key_bytes_7_T_1 ? phv_data_23 : _GEN_2606; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2608 = 8'h18 == _match_key_bytes_7_T_1 ? phv_data_24 : _GEN_2607; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2609 = 8'h19 == _match_key_bytes_7_T_1 ? phv_data_25 : _GEN_2608; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2610 = 8'h1a == _match_key_bytes_7_T_1 ? phv_data_26 : _GEN_2609; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2611 = 8'h1b == _match_key_bytes_7_T_1 ? phv_data_27 : _GEN_2610; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2612 = 8'h1c == _match_key_bytes_7_T_1 ? phv_data_28 : _GEN_2611; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2613 = 8'h1d == _match_key_bytes_7_T_1 ? phv_data_29 : _GEN_2612; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2614 = 8'h1e == _match_key_bytes_7_T_1 ? phv_data_30 : _GEN_2613; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2615 = 8'h1f == _match_key_bytes_7_T_1 ? phv_data_31 : _GEN_2614; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2616 = 8'h20 == _match_key_bytes_7_T_1 ? phv_data_32 : _GEN_2615; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2617 = 8'h21 == _match_key_bytes_7_T_1 ? phv_data_33 : _GEN_2616; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2618 = 8'h22 == _match_key_bytes_7_T_1 ? phv_data_34 : _GEN_2617; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2619 = 8'h23 == _match_key_bytes_7_T_1 ? phv_data_35 : _GEN_2618; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2620 = 8'h24 == _match_key_bytes_7_T_1 ? phv_data_36 : _GEN_2619; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2621 = 8'h25 == _match_key_bytes_7_T_1 ? phv_data_37 : _GEN_2620; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2622 = 8'h26 == _match_key_bytes_7_T_1 ? phv_data_38 : _GEN_2621; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2623 = 8'h27 == _match_key_bytes_7_T_1 ? phv_data_39 : _GEN_2622; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2624 = 8'h28 == _match_key_bytes_7_T_1 ? phv_data_40 : _GEN_2623; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2625 = 8'h29 == _match_key_bytes_7_T_1 ? phv_data_41 : _GEN_2624; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2626 = 8'h2a == _match_key_bytes_7_T_1 ? phv_data_42 : _GEN_2625; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2627 = 8'h2b == _match_key_bytes_7_T_1 ? phv_data_43 : _GEN_2626; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2628 = 8'h2c == _match_key_bytes_7_T_1 ? phv_data_44 : _GEN_2627; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2629 = 8'h2d == _match_key_bytes_7_T_1 ? phv_data_45 : _GEN_2628; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2630 = 8'h2e == _match_key_bytes_7_T_1 ? phv_data_46 : _GEN_2629; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2631 = 8'h2f == _match_key_bytes_7_T_1 ? phv_data_47 : _GEN_2630; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2632 = 8'h30 == _match_key_bytes_7_T_1 ? phv_data_48 : _GEN_2631; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2633 = 8'h31 == _match_key_bytes_7_T_1 ? phv_data_49 : _GEN_2632; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2634 = 8'h32 == _match_key_bytes_7_T_1 ? phv_data_50 : _GEN_2633; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2635 = 8'h33 == _match_key_bytes_7_T_1 ? phv_data_51 : _GEN_2634; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2636 = 8'h34 == _match_key_bytes_7_T_1 ? phv_data_52 : _GEN_2635; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2637 = 8'h35 == _match_key_bytes_7_T_1 ? phv_data_53 : _GEN_2636; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2638 = 8'h36 == _match_key_bytes_7_T_1 ? phv_data_54 : _GEN_2637; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2639 = 8'h37 == _match_key_bytes_7_T_1 ? phv_data_55 : _GEN_2638; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2640 = 8'h38 == _match_key_bytes_7_T_1 ? phv_data_56 : _GEN_2639; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2641 = 8'h39 == _match_key_bytes_7_T_1 ? phv_data_57 : _GEN_2640; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2642 = 8'h3a == _match_key_bytes_7_T_1 ? phv_data_58 : _GEN_2641; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2643 = 8'h3b == _match_key_bytes_7_T_1 ? phv_data_59 : _GEN_2642; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2644 = 8'h3c == _match_key_bytes_7_T_1 ? phv_data_60 : _GEN_2643; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2645 = 8'h3d == _match_key_bytes_7_T_1 ? phv_data_61 : _GEN_2644; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2646 = 8'h3e == _match_key_bytes_7_T_1 ? phv_data_62 : _GEN_2645; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2647 = 8'h3f == _match_key_bytes_7_T_1 ? phv_data_63 : _GEN_2646; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2648 = 8'h40 == _match_key_bytes_7_T_1 ? phv_data_64 : _GEN_2647; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2649 = 8'h41 == _match_key_bytes_7_T_1 ? phv_data_65 : _GEN_2648; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2650 = 8'h42 == _match_key_bytes_7_T_1 ? phv_data_66 : _GEN_2649; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2651 = 8'h43 == _match_key_bytes_7_T_1 ? phv_data_67 : _GEN_2650; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2652 = 8'h44 == _match_key_bytes_7_T_1 ? phv_data_68 : _GEN_2651; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2653 = 8'h45 == _match_key_bytes_7_T_1 ? phv_data_69 : _GEN_2652; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2654 = 8'h46 == _match_key_bytes_7_T_1 ? phv_data_70 : _GEN_2653; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2655 = 8'h47 == _match_key_bytes_7_T_1 ? phv_data_71 : _GEN_2654; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2656 = 8'h48 == _match_key_bytes_7_T_1 ? phv_data_72 : _GEN_2655; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2657 = 8'h49 == _match_key_bytes_7_T_1 ? phv_data_73 : _GEN_2656; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2658 = 8'h4a == _match_key_bytes_7_T_1 ? phv_data_74 : _GEN_2657; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2659 = 8'h4b == _match_key_bytes_7_T_1 ? phv_data_75 : _GEN_2658; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2660 = 8'h4c == _match_key_bytes_7_T_1 ? phv_data_76 : _GEN_2659; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2661 = 8'h4d == _match_key_bytes_7_T_1 ? phv_data_77 : _GEN_2660; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2662 = 8'h4e == _match_key_bytes_7_T_1 ? phv_data_78 : _GEN_2661; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2663 = 8'h4f == _match_key_bytes_7_T_1 ? phv_data_79 : _GEN_2662; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2664 = 8'h50 == _match_key_bytes_7_T_1 ? phv_data_80 : _GEN_2663; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2665 = 8'h51 == _match_key_bytes_7_T_1 ? phv_data_81 : _GEN_2664; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2666 = 8'h52 == _match_key_bytes_7_T_1 ? phv_data_82 : _GEN_2665; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2667 = 8'h53 == _match_key_bytes_7_T_1 ? phv_data_83 : _GEN_2666; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2668 = 8'h54 == _match_key_bytes_7_T_1 ? phv_data_84 : _GEN_2667; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2669 = 8'h55 == _match_key_bytes_7_T_1 ? phv_data_85 : _GEN_2668; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2670 = 8'h56 == _match_key_bytes_7_T_1 ? phv_data_86 : _GEN_2669; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2671 = 8'h57 == _match_key_bytes_7_T_1 ? phv_data_87 : _GEN_2670; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2672 = 8'h58 == _match_key_bytes_7_T_1 ? phv_data_88 : _GEN_2671; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2673 = 8'h59 == _match_key_bytes_7_T_1 ? phv_data_89 : _GEN_2672; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2674 = 8'h5a == _match_key_bytes_7_T_1 ? phv_data_90 : _GEN_2673; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2675 = 8'h5b == _match_key_bytes_7_T_1 ? phv_data_91 : _GEN_2674; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2676 = 8'h5c == _match_key_bytes_7_T_1 ? phv_data_92 : _GEN_2675; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2677 = 8'h5d == _match_key_bytes_7_T_1 ? phv_data_93 : _GEN_2676; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2678 = 8'h5e == _match_key_bytes_7_T_1 ? phv_data_94 : _GEN_2677; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2679 = 8'h5f == _match_key_bytes_7_T_1 ? phv_data_95 : _GEN_2678; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2680 = 8'h60 == _match_key_bytes_7_T_1 ? phv_data_96 : _GEN_2679; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2681 = 8'h61 == _match_key_bytes_7_T_1 ? phv_data_97 : _GEN_2680; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2682 = 8'h62 == _match_key_bytes_7_T_1 ? phv_data_98 : _GEN_2681; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2683 = 8'h63 == _match_key_bytes_7_T_1 ? phv_data_99 : _GEN_2682; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2684 = 8'h64 == _match_key_bytes_7_T_1 ? phv_data_100 : _GEN_2683; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2685 = 8'h65 == _match_key_bytes_7_T_1 ? phv_data_101 : _GEN_2684; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2686 = 8'h66 == _match_key_bytes_7_T_1 ? phv_data_102 : _GEN_2685; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2687 = 8'h67 == _match_key_bytes_7_T_1 ? phv_data_103 : _GEN_2686; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2688 = 8'h68 == _match_key_bytes_7_T_1 ? phv_data_104 : _GEN_2687; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2689 = 8'h69 == _match_key_bytes_7_T_1 ? phv_data_105 : _GEN_2688; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2690 = 8'h6a == _match_key_bytes_7_T_1 ? phv_data_106 : _GEN_2689; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2691 = 8'h6b == _match_key_bytes_7_T_1 ? phv_data_107 : _GEN_2690; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2692 = 8'h6c == _match_key_bytes_7_T_1 ? phv_data_108 : _GEN_2691; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2693 = 8'h6d == _match_key_bytes_7_T_1 ? phv_data_109 : _GEN_2692; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2694 = 8'h6e == _match_key_bytes_7_T_1 ? phv_data_110 : _GEN_2693; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2695 = 8'h6f == _match_key_bytes_7_T_1 ? phv_data_111 : _GEN_2694; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2696 = 8'h70 == _match_key_bytes_7_T_1 ? phv_data_112 : _GEN_2695; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2697 = 8'h71 == _match_key_bytes_7_T_1 ? phv_data_113 : _GEN_2696; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2698 = 8'h72 == _match_key_bytes_7_T_1 ? phv_data_114 : _GEN_2697; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2699 = 8'h73 == _match_key_bytes_7_T_1 ? phv_data_115 : _GEN_2698; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2700 = 8'h74 == _match_key_bytes_7_T_1 ? phv_data_116 : _GEN_2699; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2701 = 8'h75 == _match_key_bytes_7_T_1 ? phv_data_117 : _GEN_2700; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2702 = 8'h76 == _match_key_bytes_7_T_1 ? phv_data_118 : _GEN_2701; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2703 = 8'h77 == _match_key_bytes_7_T_1 ? phv_data_119 : _GEN_2702; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2704 = 8'h78 == _match_key_bytes_7_T_1 ? phv_data_120 : _GEN_2703; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2705 = 8'h79 == _match_key_bytes_7_T_1 ? phv_data_121 : _GEN_2704; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2706 = 8'h7a == _match_key_bytes_7_T_1 ? phv_data_122 : _GEN_2705; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2707 = 8'h7b == _match_key_bytes_7_T_1 ? phv_data_123 : _GEN_2706; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2708 = 8'h7c == _match_key_bytes_7_T_1 ? phv_data_124 : _GEN_2707; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2709 = 8'h7d == _match_key_bytes_7_T_1 ? phv_data_125 : _GEN_2708; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2710 = 8'h7e == _match_key_bytes_7_T_1 ? phv_data_126 : _GEN_2709; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2711 = 8'h7f == _match_key_bytes_7_T_1 ? phv_data_127 : _GEN_2710; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2712 = 8'h80 == _match_key_bytes_7_T_1 ? phv_data_128 : _GEN_2711; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2713 = 8'h81 == _match_key_bytes_7_T_1 ? phv_data_129 : _GEN_2712; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2714 = 8'h82 == _match_key_bytes_7_T_1 ? phv_data_130 : _GEN_2713; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2715 = 8'h83 == _match_key_bytes_7_T_1 ? phv_data_131 : _GEN_2714; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2716 = 8'h84 == _match_key_bytes_7_T_1 ? phv_data_132 : _GEN_2715; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2717 = 8'h85 == _match_key_bytes_7_T_1 ? phv_data_133 : _GEN_2716; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2718 = 8'h86 == _match_key_bytes_7_T_1 ? phv_data_134 : _GEN_2717; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2719 = 8'h87 == _match_key_bytes_7_T_1 ? phv_data_135 : _GEN_2718; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2720 = 8'h88 == _match_key_bytes_7_T_1 ? phv_data_136 : _GEN_2719; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2721 = 8'h89 == _match_key_bytes_7_T_1 ? phv_data_137 : _GEN_2720; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2722 = 8'h8a == _match_key_bytes_7_T_1 ? phv_data_138 : _GEN_2721; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2723 = 8'h8b == _match_key_bytes_7_T_1 ? phv_data_139 : _GEN_2722; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2724 = 8'h8c == _match_key_bytes_7_T_1 ? phv_data_140 : _GEN_2723; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2725 = 8'h8d == _match_key_bytes_7_T_1 ? phv_data_141 : _GEN_2724; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2726 = 8'h8e == _match_key_bytes_7_T_1 ? phv_data_142 : _GEN_2725; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2727 = 8'h8f == _match_key_bytes_7_T_1 ? phv_data_143 : _GEN_2726; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2728 = 8'h90 == _match_key_bytes_7_T_1 ? phv_data_144 : _GEN_2727; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2729 = 8'h91 == _match_key_bytes_7_T_1 ? phv_data_145 : _GEN_2728; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2730 = 8'h92 == _match_key_bytes_7_T_1 ? phv_data_146 : _GEN_2729; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2731 = 8'h93 == _match_key_bytes_7_T_1 ? phv_data_147 : _GEN_2730; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2732 = 8'h94 == _match_key_bytes_7_T_1 ? phv_data_148 : _GEN_2731; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2733 = 8'h95 == _match_key_bytes_7_T_1 ? phv_data_149 : _GEN_2732; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2734 = 8'h96 == _match_key_bytes_7_T_1 ? phv_data_150 : _GEN_2733; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2735 = 8'h97 == _match_key_bytes_7_T_1 ? phv_data_151 : _GEN_2734; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2736 = 8'h98 == _match_key_bytes_7_T_1 ? phv_data_152 : _GEN_2735; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2737 = 8'h99 == _match_key_bytes_7_T_1 ? phv_data_153 : _GEN_2736; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2738 = 8'h9a == _match_key_bytes_7_T_1 ? phv_data_154 : _GEN_2737; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2739 = 8'h9b == _match_key_bytes_7_T_1 ? phv_data_155 : _GEN_2738; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2740 = 8'h9c == _match_key_bytes_7_T_1 ? phv_data_156 : _GEN_2739; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2741 = 8'h9d == _match_key_bytes_7_T_1 ? phv_data_157 : _GEN_2740; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2742 = 8'h9e == _match_key_bytes_7_T_1 ? phv_data_158 : _GEN_2741; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2743 = 8'h9f == _match_key_bytes_7_T_1 ? phv_data_159 : _GEN_2742; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_7 = 8'h10 < _GEN_6 ? _GEN_2743 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_6_T_1 = key_offset + 8'h11; // @[matcher.scala 72:98]
  wire [7:0] _GEN_2746 = 8'h1 == _match_key_bytes_6_T_1 ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2747 = 8'h2 == _match_key_bytes_6_T_1 ? phv_data_2 : _GEN_2746; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2748 = 8'h3 == _match_key_bytes_6_T_1 ? phv_data_3 : _GEN_2747; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2749 = 8'h4 == _match_key_bytes_6_T_1 ? phv_data_4 : _GEN_2748; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2750 = 8'h5 == _match_key_bytes_6_T_1 ? phv_data_5 : _GEN_2749; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2751 = 8'h6 == _match_key_bytes_6_T_1 ? phv_data_6 : _GEN_2750; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2752 = 8'h7 == _match_key_bytes_6_T_1 ? phv_data_7 : _GEN_2751; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2753 = 8'h8 == _match_key_bytes_6_T_1 ? phv_data_8 : _GEN_2752; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2754 = 8'h9 == _match_key_bytes_6_T_1 ? phv_data_9 : _GEN_2753; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2755 = 8'ha == _match_key_bytes_6_T_1 ? phv_data_10 : _GEN_2754; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2756 = 8'hb == _match_key_bytes_6_T_1 ? phv_data_11 : _GEN_2755; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2757 = 8'hc == _match_key_bytes_6_T_1 ? phv_data_12 : _GEN_2756; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2758 = 8'hd == _match_key_bytes_6_T_1 ? phv_data_13 : _GEN_2757; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2759 = 8'he == _match_key_bytes_6_T_1 ? phv_data_14 : _GEN_2758; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2760 = 8'hf == _match_key_bytes_6_T_1 ? phv_data_15 : _GEN_2759; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2761 = 8'h10 == _match_key_bytes_6_T_1 ? phv_data_16 : _GEN_2760; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2762 = 8'h11 == _match_key_bytes_6_T_1 ? phv_data_17 : _GEN_2761; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2763 = 8'h12 == _match_key_bytes_6_T_1 ? phv_data_18 : _GEN_2762; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2764 = 8'h13 == _match_key_bytes_6_T_1 ? phv_data_19 : _GEN_2763; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2765 = 8'h14 == _match_key_bytes_6_T_1 ? phv_data_20 : _GEN_2764; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2766 = 8'h15 == _match_key_bytes_6_T_1 ? phv_data_21 : _GEN_2765; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2767 = 8'h16 == _match_key_bytes_6_T_1 ? phv_data_22 : _GEN_2766; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2768 = 8'h17 == _match_key_bytes_6_T_1 ? phv_data_23 : _GEN_2767; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2769 = 8'h18 == _match_key_bytes_6_T_1 ? phv_data_24 : _GEN_2768; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2770 = 8'h19 == _match_key_bytes_6_T_1 ? phv_data_25 : _GEN_2769; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2771 = 8'h1a == _match_key_bytes_6_T_1 ? phv_data_26 : _GEN_2770; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2772 = 8'h1b == _match_key_bytes_6_T_1 ? phv_data_27 : _GEN_2771; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2773 = 8'h1c == _match_key_bytes_6_T_1 ? phv_data_28 : _GEN_2772; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2774 = 8'h1d == _match_key_bytes_6_T_1 ? phv_data_29 : _GEN_2773; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2775 = 8'h1e == _match_key_bytes_6_T_1 ? phv_data_30 : _GEN_2774; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2776 = 8'h1f == _match_key_bytes_6_T_1 ? phv_data_31 : _GEN_2775; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2777 = 8'h20 == _match_key_bytes_6_T_1 ? phv_data_32 : _GEN_2776; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2778 = 8'h21 == _match_key_bytes_6_T_1 ? phv_data_33 : _GEN_2777; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2779 = 8'h22 == _match_key_bytes_6_T_1 ? phv_data_34 : _GEN_2778; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2780 = 8'h23 == _match_key_bytes_6_T_1 ? phv_data_35 : _GEN_2779; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2781 = 8'h24 == _match_key_bytes_6_T_1 ? phv_data_36 : _GEN_2780; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2782 = 8'h25 == _match_key_bytes_6_T_1 ? phv_data_37 : _GEN_2781; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2783 = 8'h26 == _match_key_bytes_6_T_1 ? phv_data_38 : _GEN_2782; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2784 = 8'h27 == _match_key_bytes_6_T_1 ? phv_data_39 : _GEN_2783; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2785 = 8'h28 == _match_key_bytes_6_T_1 ? phv_data_40 : _GEN_2784; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2786 = 8'h29 == _match_key_bytes_6_T_1 ? phv_data_41 : _GEN_2785; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2787 = 8'h2a == _match_key_bytes_6_T_1 ? phv_data_42 : _GEN_2786; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2788 = 8'h2b == _match_key_bytes_6_T_1 ? phv_data_43 : _GEN_2787; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2789 = 8'h2c == _match_key_bytes_6_T_1 ? phv_data_44 : _GEN_2788; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2790 = 8'h2d == _match_key_bytes_6_T_1 ? phv_data_45 : _GEN_2789; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2791 = 8'h2e == _match_key_bytes_6_T_1 ? phv_data_46 : _GEN_2790; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2792 = 8'h2f == _match_key_bytes_6_T_1 ? phv_data_47 : _GEN_2791; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2793 = 8'h30 == _match_key_bytes_6_T_1 ? phv_data_48 : _GEN_2792; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2794 = 8'h31 == _match_key_bytes_6_T_1 ? phv_data_49 : _GEN_2793; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2795 = 8'h32 == _match_key_bytes_6_T_1 ? phv_data_50 : _GEN_2794; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2796 = 8'h33 == _match_key_bytes_6_T_1 ? phv_data_51 : _GEN_2795; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2797 = 8'h34 == _match_key_bytes_6_T_1 ? phv_data_52 : _GEN_2796; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2798 = 8'h35 == _match_key_bytes_6_T_1 ? phv_data_53 : _GEN_2797; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2799 = 8'h36 == _match_key_bytes_6_T_1 ? phv_data_54 : _GEN_2798; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2800 = 8'h37 == _match_key_bytes_6_T_1 ? phv_data_55 : _GEN_2799; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2801 = 8'h38 == _match_key_bytes_6_T_1 ? phv_data_56 : _GEN_2800; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2802 = 8'h39 == _match_key_bytes_6_T_1 ? phv_data_57 : _GEN_2801; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2803 = 8'h3a == _match_key_bytes_6_T_1 ? phv_data_58 : _GEN_2802; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2804 = 8'h3b == _match_key_bytes_6_T_1 ? phv_data_59 : _GEN_2803; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2805 = 8'h3c == _match_key_bytes_6_T_1 ? phv_data_60 : _GEN_2804; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2806 = 8'h3d == _match_key_bytes_6_T_1 ? phv_data_61 : _GEN_2805; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2807 = 8'h3e == _match_key_bytes_6_T_1 ? phv_data_62 : _GEN_2806; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2808 = 8'h3f == _match_key_bytes_6_T_1 ? phv_data_63 : _GEN_2807; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2809 = 8'h40 == _match_key_bytes_6_T_1 ? phv_data_64 : _GEN_2808; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2810 = 8'h41 == _match_key_bytes_6_T_1 ? phv_data_65 : _GEN_2809; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2811 = 8'h42 == _match_key_bytes_6_T_1 ? phv_data_66 : _GEN_2810; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2812 = 8'h43 == _match_key_bytes_6_T_1 ? phv_data_67 : _GEN_2811; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2813 = 8'h44 == _match_key_bytes_6_T_1 ? phv_data_68 : _GEN_2812; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2814 = 8'h45 == _match_key_bytes_6_T_1 ? phv_data_69 : _GEN_2813; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2815 = 8'h46 == _match_key_bytes_6_T_1 ? phv_data_70 : _GEN_2814; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2816 = 8'h47 == _match_key_bytes_6_T_1 ? phv_data_71 : _GEN_2815; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2817 = 8'h48 == _match_key_bytes_6_T_1 ? phv_data_72 : _GEN_2816; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2818 = 8'h49 == _match_key_bytes_6_T_1 ? phv_data_73 : _GEN_2817; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2819 = 8'h4a == _match_key_bytes_6_T_1 ? phv_data_74 : _GEN_2818; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2820 = 8'h4b == _match_key_bytes_6_T_1 ? phv_data_75 : _GEN_2819; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2821 = 8'h4c == _match_key_bytes_6_T_1 ? phv_data_76 : _GEN_2820; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2822 = 8'h4d == _match_key_bytes_6_T_1 ? phv_data_77 : _GEN_2821; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2823 = 8'h4e == _match_key_bytes_6_T_1 ? phv_data_78 : _GEN_2822; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2824 = 8'h4f == _match_key_bytes_6_T_1 ? phv_data_79 : _GEN_2823; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2825 = 8'h50 == _match_key_bytes_6_T_1 ? phv_data_80 : _GEN_2824; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2826 = 8'h51 == _match_key_bytes_6_T_1 ? phv_data_81 : _GEN_2825; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2827 = 8'h52 == _match_key_bytes_6_T_1 ? phv_data_82 : _GEN_2826; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2828 = 8'h53 == _match_key_bytes_6_T_1 ? phv_data_83 : _GEN_2827; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2829 = 8'h54 == _match_key_bytes_6_T_1 ? phv_data_84 : _GEN_2828; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2830 = 8'h55 == _match_key_bytes_6_T_1 ? phv_data_85 : _GEN_2829; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2831 = 8'h56 == _match_key_bytes_6_T_1 ? phv_data_86 : _GEN_2830; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2832 = 8'h57 == _match_key_bytes_6_T_1 ? phv_data_87 : _GEN_2831; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2833 = 8'h58 == _match_key_bytes_6_T_1 ? phv_data_88 : _GEN_2832; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2834 = 8'h59 == _match_key_bytes_6_T_1 ? phv_data_89 : _GEN_2833; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2835 = 8'h5a == _match_key_bytes_6_T_1 ? phv_data_90 : _GEN_2834; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2836 = 8'h5b == _match_key_bytes_6_T_1 ? phv_data_91 : _GEN_2835; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2837 = 8'h5c == _match_key_bytes_6_T_1 ? phv_data_92 : _GEN_2836; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2838 = 8'h5d == _match_key_bytes_6_T_1 ? phv_data_93 : _GEN_2837; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2839 = 8'h5e == _match_key_bytes_6_T_1 ? phv_data_94 : _GEN_2838; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2840 = 8'h5f == _match_key_bytes_6_T_1 ? phv_data_95 : _GEN_2839; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2841 = 8'h60 == _match_key_bytes_6_T_1 ? phv_data_96 : _GEN_2840; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2842 = 8'h61 == _match_key_bytes_6_T_1 ? phv_data_97 : _GEN_2841; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2843 = 8'h62 == _match_key_bytes_6_T_1 ? phv_data_98 : _GEN_2842; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2844 = 8'h63 == _match_key_bytes_6_T_1 ? phv_data_99 : _GEN_2843; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2845 = 8'h64 == _match_key_bytes_6_T_1 ? phv_data_100 : _GEN_2844; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2846 = 8'h65 == _match_key_bytes_6_T_1 ? phv_data_101 : _GEN_2845; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2847 = 8'h66 == _match_key_bytes_6_T_1 ? phv_data_102 : _GEN_2846; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2848 = 8'h67 == _match_key_bytes_6_T_1 ? phv_data_103 : _GEN_2847; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2849 = 8'h68 == _match_key_bytes_6_T_1 ? phv_data_104 : _GEN_2848; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2850 = 8'h69 == _match_key_bytes_6_T_1 ? phv_data_105 : _GEN_2849; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2851 = 8'h6a == _match_key_bytes_6_T_1 ? phv_data_106 : _GEN_2850; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2852 = 8'h6b == _match_key_bytes_6_T_1 ? phv_data_107 : _GEN_2851; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2853 = 8'h6c == _match_key_bytes_6_T_1 ? phv_data_108 : _GEN_2852; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2854 = 8'h6d == _match_key_bytes_6_T_1 ? phv_data_109 : _GEN_2853; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2855 = 8'h6e == _match_key_bytes_6_T_1 ? phv_data_110 : _GEN_2854; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2856 = 8'h6f == _match_key_bytes_6_T_1 ? phv_data_111 : _GEN_2855; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2857 = 8'h70 == _match_key_bytes_6_T_1 ? phv_data_112 : _GEN_2856; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2858 = 8'h71 == _match_key_bytes_6_T_1 ? phv_data_113 : _GEN_2857; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2859 = 8'h72 == _match_key_bytes_6_T_1 ? phv_data_114 : _GEN_2858; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2860 = 8'h73 == _match_key_bytes_6_T_1 ? phv_data_115 : _GEN_2859; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2861 = 8'h74 == _match_key_bytes_6_T_1 ? phv_data_116 : _GEN_2860; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2862 = 8'h75 == _match_key_bytes_6_T_1 ? phv_data_117 : _GEN_2861; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2863 = 8'h76 == _match_key_bytes_6_T_1 ? phv_data_118 : _GEN_2862; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2864 = 8'h77 == _match_key_bytes_6_T_1 ? phv_data_119 : _GEN_2863; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2865 = 8'h78 == _match_key_bytes_6_T_1 ? phv_data_120 : _GEN_2864; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2866 = 8'h79 == _match_key_bytes_6_T_1 ? phv_data_121 : _GEN_2865; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2867 = 8'h7a == _match_key_bytes_6_T_1 ? phv_data_122 : _GEN_2866; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2868 = 8'h7b == _match_key_bytes_6_T_1 ? phv_data_123 : _GEN_2867; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2869 = 8'h7c == _match_key_bytes_6_T_1 ? phv_data_124 : _GEN_2868; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2870 = 8'h7d == _match_key_bytes_6_T_1 ? phv_data_125 : _GEN_2869; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2871 = 8'h7e == _match_key_bytes_6_T_1 ? phv_data_126 : _GEN_2870; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2872 = 8'h7f == _match_key_bytes_6_T_1 ? phv_data_127 : _GEN_2871; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2873 = 8'h80 == _match_key_bytes_6_T_1 ? phv_data_128 : _GEN_2872; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2874 = 8'h81 == _match_key_bytes_6_T_1 ? phv_data_129 : _GEN_2873; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2875 = 8'h82 == _match_key_bytes_6_T_1 ? phv_data_130 : _GEN_2874; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2876 = 8'h83 == _match_key_bytes_6_T_1 ? phv_data_131 : _GEN_2875; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2877 = 8'h84 == _match_key_bytes_6_T_1 ? phv_data_132 : _GEN_2876; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2878 = 8'h85 == _match_key_bytes_6_T_1 ? phv_data_133 : _GEN_2877; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2879 = 8'h86 == _match_key_bytes_6_T_1 ? phv_data_134 : _GEN_2878; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2880 = 8'h87 == _match_key_bytes_6_T_1 ? phv_data_135 : _GEN_2879; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2881 = 8'h88 == _match_key_bytes_6_T_1 ? phv_data_136 : _GEN_2880; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2882 = 8'h89 == _match_key_bytes_6_T_1 ? phv_data_137 : _GEN_2881; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2883 = 8'h8a == _match_key_bytes_6_T_1 ? phv_data_138 : _GEN_2882; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2884 = 8'h8b == _match_key_bytes_6_T_1 ? phv_data_139 : _GEN_2883; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2885 = 8'h8c == _match_key_bytes_6_T_1 ? phv_data_140 : _GEN_2884; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2886 = 8'h8d == _match_key_bytes_6_T_1 ? phv_data_141 : _GEN_2885; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2887 = 8'h8e == _match_key_bytes_6_T_1 ? phv_data_142 : _GEN_2886; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2888 = 8'h8f == _match_key_bytes_6_T_1 ? phv_data_143 : _GEN_2887; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2889 = 8'h90 == _match_key_bytes_6_T_1 ? phv_data_144 : _GEN_2888; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2890 = 8'h91 == _match_key_bytes_6_T_1 ? phv_data_145 : _GEN_2889; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2891 = 8'h92 == _match_key_bytes_6_T_1 ? phv_data_146 : _GEN_2890; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2892 = 8'h93 == _match_key_bytes_6_T_1 ? phv_data_147 : _GEN_2891; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2893 = 8'h94 == _match_key_bytes_6_T_1 ? phv_data_148 : _GEN_2892; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2894 = 8'h95 == _match_key_bytes_6_T_1 ? phv_data_149 : _GEN_2893; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2895 = 8'h96 == _match_key_bytes_6_T_1 ? phv_data_150 : _GEN_2894; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2896 = 8'h97 == _match_key_bytes_6_T_1 ? phv_data_151 : _GEN_2895; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2897 = 8'h98 == _match_key_bytes_6_T_1 ? phv_data_152 : _GEN_2896; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2898 = 8'h99 == _match_key_bytes_6_T_1 ? phv_data_153 : _GEN_2897; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2899 = 8'h9a == _match_key_bytes_6_T_1 ? phv_data_154 : _GEN_2898; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2900 = 8'h9b == _match_key_bytes_6_T_1 ? phv_data_155 : _GEN_2899; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2901 = 8'h9c == _match_key_bytes_6_T_1 ? phv_data_156 : _GEN_2900; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2902 = 8'h9d == _match_key_bytes_6_T_1 ? phv_data_157 : _GEN_2901; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2903 = 8'h9e == _match_key_bytes_6_T_1 ? phv_data_158 : _GEN_2902; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2904 = 8'h9f == _match_key_bytes_6_T_1 ? phv_data_159 : _GEN_2903; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_6 = 8'h11 < _GEN_6 ? _GEN_2904 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_5_T_1 = key_offset + 8'h12; // @[matcher.scala 72:98]
  wire [7:0] _GEN_2907 = 8'h1 == _match_key_bytes_5_T_1 ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2908 = 8'h2 == _match_key_bytes_5_T_1 ? phv_data_2 : _GEN_2907; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2909 = 8'h3 == _match_key_bytes_5_T_1 ? phv_data_3 : _GEN_2908; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2910 = 8'h4 == _match_key_bytes_5_T_1 ? phv_data_4 : _GEN_2909; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2911 = 8'h5 == _match_key_bytes_5_T_1 ? phv_data_5 : _GEN_2910; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2912 = 8'h6 == _match_key_bytes_5_T_1 ? phv_data_6 : _GEN_2911; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2913 = 8'h7 == _match_key_bytes_5_T_1 ? phv_data_7 : _GEN_2912; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2914 = 8'h8 == _match_key_bytes_5_T_1 ? phv_data_8 : _GEN_2913; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2915 = 8'h9 == _match_key_bytes_5_T_1 ? phv_data_9 : _GEN_2914; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2916 = 8'ha == _match_key_bytes_5_T_1 ? phv_data_10 : _GEN_2915; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2917 = 8'hb == _match_key_bytes_5_T_1 ? phv_data_11 : _GEN_2916; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2918 = 8'hc == _match_key_bytes_5_T_1 ? phv_data_12 : _GEN_2917; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2919 = 8'hd == _match_key_bytes_5_T_1 ? phv_data_13 : _GEN_2918; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2920 = 8'he == _match_key_bytes_5_T_1 ? phv_data_14 : _GEN_2919; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2921 = 8'hf == _match_key_bytes_5_T_1 ? phv_data_15 : _GEN_2920; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2922 = 8'h10 == _match_key_bytes_5_T_1 ? phv_data_16 : _GEN_2921; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2923 = 8'h11 == _match_key_bytes_5_T_1 ? phv_data_17 : _GEN_2922; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2924 = 8'h12 == _match_key_bytes_5_T_1 ? phv_data_18 : _GEN_2923; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2925 = 8'h13 == _match_key_bytes_5_T_1 ? phv_data_19 : _GEN_2924; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2926 = 8'h14 == _match_key_bytes_5_T_1 ? phv_data_20 : _GEN_2925; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2927 = 8'h15 == _match_key_bytes_5_T_1 ? phv_data_21 : _GEN_2926; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2928 = 8'h16 == _match_key_bytes_5_T_1 ? phv_data_22 : _GEN_2927; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2929 = 8'h17 == _match_key_bytes_5_T_1 ? phv_data_23 : _GEN_2928; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2930 = 8'h18 == _match_key_bytes_5_T_1 ? phv_data_24 : _GEN_2929; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2931 = 8'h19 == _match_key_bytes_5_T_1 ? phv_data_25 : _GEN_2930; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2932 = 8'h1a == _match_key_bytes_5_T_1 ? phv_data_26 : _GEN_2931; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2933 = 8'h1b == _match_key_bytes_5_T_1 ? phv_data_27 : _GEN_2932; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2934 = 8'h1c == _match_key_bytes_5_T_1 ? phv_data_28 : _GEN_2933; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2935 = 8'h1d == _match_key_bytes_5_T_1 ? phv_data_29 : _GEN_2934; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2936 = 8'h1e == _match_key_bytes_5_T_1 ? phv_data_30 : _GEN_2935; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2937 = 8'h1f == _match_key_bytes_5_T_1 ? phv_data_31 : _GEN_2936; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2938 = 8'h20 == _match_key_bytes_5_T_1 ? phv_data_32 : _GEN_2937; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2939 = 8'h21 == _match_key_bytes_5_T_1 ? phv_data_33 : _GEN_2938; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2940 = 8'h22 == _match_key_bytes_5_T_1 ? phv_data_34 : _GEN_2939; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2941 = 8'h23 == _match_key_bytes_5_T_1 ? phv_data_35 : _GEN_2940; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2942 = 8'h24 == _match_key_bytes_5_T_1 ? phv_data_36 : _GEN_2941; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2943 = 8'h25 == _match_key_bytes_5_T_1 ? phv_data_37 : _GEN_2942; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2944 = 8'h26 == _match_key_bytes_5_T_1 ? phv_data_38 : _GEN_2943; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2945 = 8'h27 == _match_key_bytes_5_T_1 ? phv_data_39 : _GEN_2944; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2946 = 8'h28 == _match_key_bytes_5_T_1 ? phv_data_40 : _GEN_2945; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2947 = 8'h29 == _match_key_bytes_5_T_1 ? phv_data_41 : _GEN_2946; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2948 = 8'h2a == _match_key_bytes_5_T_1 ? phv_data_42 : _GEN_2947; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2949 = 8'h2b == _match_key_bytes_5_T_1 ? phv_data_43 : _GEN_2948; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2950 = 8'h2c == _match_key_bytes_5_T_1 ? phv_data_44 : _GEN_2949; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2951 = 8'h2d == _match_key_bytes_5_T_1 ? phv_data_45 : _GEN_2950; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2952 = 8'h2e == _match_key_bytes_5_T_1 ? phv_data_46 : _GEN_2951; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2953 = 8'h2f == _match_key_bytes_5_T_1 ? phv_data_47 : _GEN_2952; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2954 = 8'h30 == _match_key_bytes_5_T_1 ? phv_data_48 : _GEN_2953; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2955 = 8'h31 == _match_key_bytes_5_T_1 ? phv_data_49 : _GEN_2954; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2956 = 8'h32 == _match_key_bytes_5_T_1 ? phv_data_50 : _GEN_2955; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2957 = 8'h33 == _match_key_bytes_5_T_1 ? phv_data_51 : _GEN_2956; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2958 = 8'h34 == _match_key_bytes_5_T_1 ? phv_data_52 : _GEN_2957; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2959 = 8'h35 == _match_key_bytes_5_T_1 ? phv_data_53 : _GEN_2958; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2960 = 8'h36 == _match_key_bytes_5_T_1 ? phv_data_54 : _GEN_2959; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2961 = 8'h37 == _match_key_bytes_5_T_1 ? phv_data_55 : _GEN_2960; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2962 = 8'h38 == _match_key_bytes_5_T_1 ? phv_data_56 : _GEN_2961; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2963 = 8'h39 == _match_key_bytes_5_T_1 ? phv_data_57 : _GEN_2962; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2964 = 8'h3a == _match_key_bytes_5_T_1 ? phv_data_58 : _GEN_2963; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2965 = 8'h3b == _match_key_bytes_5_T_1 ? phv_data_59 : _GEN_2964; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2966 = 8'h3c == _match_key_bytes_5_T_1 ? phv_data_60 : _GEN_2965; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2967 = 8'h3d == _match_key_bytes_5_T_1 ? phv_data_61 : _GEN_2966; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2968 = 8'h3e == _match_key_bytes_5_T_1 ? phv_data_62 : _GEN_2967; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2969 = 8'h3f == _match_key_bytes_5_T_1 ? phv_data_63 : _GEN_2968; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2970 = 8'h40 == _match_key_bytes_5_T_1 ? phv_data_64 : _GEN_2969; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2971 = 8'h41 == _match_key_bytes_5_T_1 ? phv_data_65 : _GEN_2970; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2972 = 8'h42 == _match_key_bytes_5_T_1 ? phv_data_66 : _GEN_2971; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2973 = 8'h43 == _match_key_bytes_5_T_1 ? phv_data_67 : _GEN_2972; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2974 = 8'h44 == _match_key_bytes_5_T_1 ? phv_data_68 : _GEN_2973; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2975 = 8'h45 == _match_key_bytes_5_T_1 ? phv_data_69 : _GEN_2974; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2976 = 8'h46 == _match_key_bytes_5_T_1 ? phv_data_70 : _GEN_2975; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2977 = 8'h47 == _match_key_bytes_5_T_1 ? phv_data_71 : _GEN_2976; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2978 = 8'h48 == _match_key_bytes_5_T_1 ? phv_data_72 : _GEN_2977; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2979 = 8'h49 == _match_key_bytes_5_T_1 ? phv_data_73 : _GEN_2978; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2980 = 8'h4a == _match_key_bytes_5_T_1 ? phv_data_74 : _GEN_2979; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2981 = 8'h4b == _match_key_bytes_5_T_1 ? phv_data_75 : _GEN_2980; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2982 = 8'h4c == _match_key_bytes_5_T_1 ? phv_data_76 : _GEN_2981; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2983 = 8'h4d == _match_key_bytes_5_T_1 ? phv_data_77 : _GEN_2982; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2984 = 8'h4e == _match_key_bytes_5_T_1 ? phv_data_78 : _GEN_2983; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2985 = 8'h4f == _match_key_bytes_5_T_1 ? phv_data_79 : _GEN_2984; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2986 = 8'h50 == _match_key_bytes_5_T_1 ? phv_data_80 : _GEN_2985; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2987 = 8'h51 == _match_key_bytes_5_T_1 ? phv_data_81 : _GEN_2986; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2988 = 8'h52 == _match_key_bytes_5_T_1 ? phv_data_82 : _GEN_2987; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2989 = 8'h53 == _match_key_bytes_5_T_1 ? phv_data_83 : _GEN_2988; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2990 = 8'h54 == _match_key_bytes_5_T_1 ? phv_data_84 : _GEN_2989; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2991 = 8'h55 == _match_key_bytes_5_T_1 ? phv_data_85 : _GEN_2990; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2992 = 8'h56 == _match_key_bytes_5_T_1 ? phv_data_86 : _GEN_2991; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2993 = 8'h57 == _match_key_bytes_5_T_1 ? phv_data_87 : _GEN_2992; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2994 = 8'h58 == _match_key_bytes_5_T_1 ? phv_data_88 : _GEN_2993; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2995 = 8'h59 == _match_key_bytes_5_T_1 ? phv_data_89 : _GEN_2994; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2996 = 8'h5a == _match_key_bytes_5_T_1 ? phv_data_90 : _GEN_2995; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2997 = 8'h5b == _match_key_bytes_5_T_1 ? phv_data_91 : _GEN_2996; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2998 = 8'h5c == _match_key_bytes_5_T_1 ? phv_data_92 : _GEN_2997; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_2999 = 8'h5d == _match_key_bytes_5_T_1 ? phv_data_93 : _GEN_2998; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3000 = 8'h5e == _match_key_bytes_5_T_1 ? phv_data_94 : _GEN_2999; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3001 = 8'h5f == _match_key_bytes_5_T_1 ? phv_data_95 : _GEN_3000; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3002 = 8'h60 == _match_key_bytes_5_T_1 ? phv_data_96 : _GEN_3001; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3003 = 8'h61 == _match_key_bytes_5_T_1 ? phv_data_97 : _GEN_3002; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3004 = 8'h62 == _match_key_bytes_5_T_1 ? phv_data_98 : _GEN_3003; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3005 = 8'h63 == _match_key_bytes_5_T_1 ? phv_data_99 : _GEN_3004; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3006 = 8'h64 == _match_key_bytes_5_T_1 ? phv_data_100 : _GEN_3005; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3007 = 8'h65 == _match_key_bytes_5_T_1 ? phv_data_101 : _GEN_3006; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3008 = 8'h66 == _match_key_bytes_5_T_1 ? phv_data_102 : _GEN_3007; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3009 = 8'h67 == _match_key_bytes_5_T_1 ? phv_data_103 : _GEN_3008; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3010 = 8'h68 == _match_key_bytes_5_T_1 ? phv_data_104 : _GEN_3009; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3011 = 8'h69 == _match_key_bytes_5_T_1 ? phv_data_105 : _GEN_3010; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3012 = 8'h6a == _match_key_bytes_5_T_1 ? phv_data_106 : _GEN_3011; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3013 = 8'h6b == _match_key_bytes_5_T_1 ? phv_data_107 : _GEN_3012; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3014 = 8'h6c == _match_key_bytes_5_T_1 ? phv_data_108 : _GEN_3013; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3015 = 8'h6d == _match_key_bytes_5_T_1 ? phv_data_109 : _GEN_3014; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3016 = 8'h6e == _match_key_bytes_5_T_1 ? phv_data_110 : _GEN_3015; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3017 = 8'h6f == _match_key_bytes_5_T_1 ? phv_data_111 : _GEN_3016; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3018 = 8'h70 == _match_key_bytes_5_T_1 ? phv_data_112 : _GEN_3017; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3019 = 8'h71 == _match_key_bytes_5_T_1 ? phv_data_113 : _GEN_3018; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3020 = 8'h72 == _match_key_bytes_5_T_1 ? phv_data_114 : _GEN_3019; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3021 = 8'h73 == _match_key_bytes_5_T_1 ? phv_data_115 : _GEN_3020; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3022 = 8'h74 == _match_key_bytes_5_T_1 ? phv_data_116 : _GEN_3021; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3023 = 8'h75 == _match_key_bytes_5_T_1 ? phv_data_117 : _GEN_3022; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3024 = 8'h76 == _match_key_bytes_5_T_1 ? phv_data_118 : _GEN_3023; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3025 = 8'h77 == _match_key_bytes_5_T_1 ? phv_data_119 : _GEN_3024; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3026 = 8'h78 == _match_key_bytes_5_T_1 ? phv_data_120 : _GEN_3025; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3027 = 8'h79 == _match_key_bytes_5_T_1 ? phv_data_121 : _GEN_3026; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3028 = 8'h7a == _match_key_bytes_5_T_1 ? phv_data_122 : _GEN_3027; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3029 = 8'h7b == _match_key_bytes_5_T_1 ? phv_data_123 : _GEN_3028; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3030 = 8'h7c == _match_key_bytes_5_T_1 ? phv_data_124 : _GEN_3029; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3031 = 8'h7d == _match_key_bytes_5_T_1 ? phv_data_125 : _GEN_3030; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3032 = 8'h7e == _match_key_bytes_5_T_1 ? phv_data_126 : _GEN_3031; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3033 = 8'h7f == _match_key_bytes_5_T_1 ? phv_data_127 : _GEN_3032; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3034 = 8'h80 == _match_key_bytes_5_T_1 ? phv_data_128 : _GEN_3033; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3035 = 8'h81 == _match_key_bytes_5_T_1 ? phv_data_129 : _GEN_3034; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3036 = 8'h82 == _match_key_bytes_5_T_1 ? phv_data_130 : _GEN_3035; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3037 = 8'h83 == _match_key_bytes_5_T_1 ? phv_data_131 : _GEN_3036; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3038 = 8'h84 == _match_key_bytes_5_T_1 ? phv_data_132 : _GEN_3037; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3039 = 8'h85 == _match_key_bytes_5_T_1 ? phv_data_133 : _GEN_3038; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3040 = 8'h86 == _match_key_bytes_5_T_1 ? phv_data_134 : _GEN_3039; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3041 = 8'h87 == _match_key_bytes_5_T_1 ? phv_data_135 : _GEN_3040; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3042 = 8'h88 == _match_key_bytes_5_T_1 ? phv_data_136 : _GEN_3041; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3043 = 8'h89 == _match_key_bytes_5_T_1 ? phv_data_137 : _GEN_3042; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3044 = 8'h8a == _match_key_bytes_5_T_1 ? phv_data_138 : _GEN_3043; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3045 = 8'h8b == _match_key_bytes_5_T_1 ? phv_data_139 : _GEN_3044; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3046 = 8'h8c == _match_key_bytes_5_T_1 ? phv_data_140 : _GEN_3045; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3047 = 8'h8d == _match_key_bytes_5_T_1 ? phv_data_141 : _GEN_3046; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3048 = 8'h8e == _match_key_bytes_5_T_1 ? phv_data_142 : _GEN_3047; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3049 = 8'h8f == _match_key_bytes_5_T_1 ? phv_data_143 : _GEN_3048; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3050 = 8'h90 == _match_key_bytes_5_T_1 ? phv_data_144 : _GEN_3049; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3051 = 8'h91 == _match_key_bytes_5_T_1 ? phv_data_145 : _GEN_3050; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3052 = 8'h92 == _match_key_bytes_5_T_1 ? phv_data_146 : _GEN_3051; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3053 = 8'h93 == _match_key_bytes_5_T_1 ? phv_data_147 : _GEN_3052; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3054 = 8'h94 == _match_key_bytes_5_T_1 ? phv_data_148 : _GEN_3053; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3055 = 8'h95 == _match_key_bytes_5_T_1 ? phv_data_149 : _GEN_3054; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3056 = 8'h96 == _match_key_bytes_5_T_1 ? phv_data_150 : _GEN_3055; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3057 = 8'h97 == _match_key_bytes_5_T_1 ? phv_data_151 : _GEN_3056; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3058 = 8'h98 == _match_key_bytes_5_T_1 ? phv_data_152 : _GEN_3057; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3059 = 8'h99 == _match_key_bytes_5_T_1 ? phv_data_153 : _GEN_3058; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3060 = 8'h9a == _match_key_bytes_5_T_1 ? phv_data_154 : _GEN_3059; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3061 = 8'h9b == _match_key_bytes_5_T_1 ? phv_data_155 : _GEN_3060; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3062 = 8'h9c == _match_key_bytes_5_T_1 ? phv_data_156 : _GEN_3061; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3063 = 8'h9d == _match_key_bytes_5_T_1 ? phv_data_157 : _GEN_3062; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3064 = 8'h9e == _match_key_bytes_5_T_1 ? phv_data_158 : _GEN_3063; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3065 = 8'h9f == _match_key_bytes_5_T_1 ? phv_data_159 : _GEN_3064; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_5 = 8'h12 < _GEN_6 ? _GEN_3065 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_4_T_1 = key_offset + 8'h13; // @[matcher.scala 72:98]
  wire [7:0] _GEN_3068 = 8'h1 == _match_key_bytes_4_T_1 ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3069 = 8'h2 == _match_key_bytes_4_T_1 ? phv_data_2 : _GEN_3068; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3070 = 8'h3 == _match_key_bytes_4_T_1 ? phv_data_3 : _GEN_3069; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3071 = 8'h4 == _match_key_bytes_4_T_1 ? phv_data_4 : _GEN_3070; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3072 = 8'h5 == _match_key_bytes_4_T_1 ? phv_data_5 : _GEN_3071; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3073 = 8'h6 == _match_key_bytes_4_T_1 ? phv_data_6 : _GEN_3072; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3074 = 8'h7 == _match_key_bytes_4_T_1 ? phv_data_7 : _GEN_3073; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3075 = 8'h8 == _match_key_bytes_4_T_1 ? phv_data_8 : _GEN_3074; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3076 = 8'h9 == _match_key_bytes_4_T_1 ? phv_data_9 : _GEN_3075; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3077 = 8'ha == _match_key_bytes_4_T_1 ? phv_data_10 : _GEN_3076; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3078 = 8'hb == _match_key_bytes_4_T_1 ? phv_data_11 : _GEN_3077; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3079 = 8'hc == _match_key_bytes_4_T_1 ? phv_data_12 : _GEN_3078; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3080 = 8'hd == _match_key_bytes_4_T_1 ? phv_data_13 : _GEN_3079; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3081 = 8'he == _match_key_bytes_4_T_1 ? phv_data_14 : _GEN_3080; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3082 = 8'hf == _match_key_bytes_4_T_1 ? phv_data_15 : _GEN_3081; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3083 = 8'h10 == _match_key_bytes_4_T_1 ? phv_data_16 : _GEN_3082; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3084 = 8'h11 == _match_key_bytes_4_T_1 ? phv_data_17 : _GEN_3083; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3085 = 8'h12 == _match_key_bytes_4_T_1 ? phv_data_18 : _GEN_3084; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3086 = 8'h13 == _match_key_bytes_4_T_1 ? phv_data_19 : _GEN_3085; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3087 = 8'h14 == _match_key_bytes_4_T_1 ? phv_data_20 : _GEN_3086; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3088 = 8'h15 == _match_key_bytes_4_T_1 ? phv_data_21 : _GEN_3087; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3089 = 8'h16 == _match_key_bytes_4_T_1 ? phv_data_22 : _GEN_3088; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3090 = 8'h17 == _match_key_bytes_4_T_1 ? phv_data_23 : _GEN_3089; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3091 = 8'h18 == _match_key_bytes_4_T_1 ? phv_data_24 : _GEN_3090; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3092 = 8'h19 == _match_key_bytes_4_T_1 ? phv_data_25 : _GEN_3091; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3093 = 8'h1a == _match_key_bytes_4_T_1 ? phv_data_26 : _GEN_3092; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3094 = 8'h1b == _match_key_bytes_4_T_1 ? phv_data_27 : _GEN_3093; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3095 = 8'h1c == _match_key_bytes_4_T_1 ? phv_data_28 : _GEN_3094; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3096 = 8'h1d == _match_key_bytes_4_T_1 ? phv_data_29 : _GEN_3095; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3097 = 8'h1e == _match_key_bytes_4_T_1 ? phv_data_30 : _GEN_3096; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3098 = 8'h1f == _match_key_bytes_4_T_1 ? phv_data_31 : _GEN_3097; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3099 = 8'h20 == _match_key_bytes_4_T_1 ? phv_data_32 : _GEN_3098; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3100 = 8'h21 == _match_key_bytes_4_T_1 ? phv_data_33 : _GEN_3099; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3101 = 8'h22 == _match_key_bytes_4_T_1 ? phv_data_34 : _GEN_3100; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3102 = 8'h23 == _match_key_bytes_4_T_1 ? phv_data_35 : _GEN_3101; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3103 = 8'h24 == _match_key_bytes_4_T_1 ? phv_data_36 : _GEN_3102; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3104 = 8'h25 == _match_key_bytes_4_T_1 ? phv_data_37 : _GEN_3103; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3105 = 8'h26 == _match_key_bytes_4_T_1 ? phv_data_38 : _GEN_3104; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3106 = 8'h27 == _match_key_bytes_4_T_1 ? phv_data_39 : _GEN_3105; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3107 = 8'h28 == _match_key_bytes_4_T_1 ? phv_data_40 : _GEN_3106; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3108 = 8'h29 == _match_key_bytes_4_T_1 ? phv_data_41 : _GEN_3107; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3109 = 8'h2a == _match_key_bytes_4_T_1 ? phv_data_42 : _GEN_3108; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3110 = 8'h2b == _match_key_bytes_4_T_1 ? phv_data_43 : _GEN_3109; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3111 = 8'h2c == _match_key_bytes_4_T_1 ? phv_data_44 : _GEN_3110; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3112 = 8'h2d == _match_key_bytes_4_T_1 ? phv_data_45 : _GEN_3111; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3113 = 8'h2e == _match_key_bytes_4_T_1 ? phv_data_46 : _GEN_3112; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3114 = 8'h2f == _match_key_bytes_4_T_1 ? phv_data_47 : _GEN_3113; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3115 = 8'h30 == _match_key_bytes_4_T_1 ? phv_data_48 : _GEN_3114; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3116 = 8'h31 == _match_key_bytes_4_T_1 ? phv_data_49 : _GEN_3115; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3117 = 8'h32 == _match_key_bytes_4_T_1 ? phv_data_50 : _GEN_3116; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3118 = 8'h33 == _match_key_bytes_4_T_1 ? phv_data_51 : _GEN_3117; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3119 = 8'h34 == _match_key_bytes_4_T_1 ? phv_data_52 : _GEN_3118; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3120 = 8'h35 == _match_key_bytes_4_T_1 ? phv_data_53 : _GEN_3119; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3121 = 8'h36 == _match_key_bytes_4_T_1 ? phv_data_54 : _GEN_3120; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3122 = 8'h37 == _match_key_bytes_4_T_1 ? phv_data_55 : _GEN_3121; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3123 = 8'h38 == _match_key_bytes_4_T_1 ? phv_data_56 : _GEN_3122; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3124 = 8'h39 == _match_key_bytes_4_T_1 ? phv_data_57 : _GEN_3123; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3125 = 8'h3a == _match_key_bytes_4_T_1 ? phv_data_58 : _GEN_3124; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3126 = 8'h3b == _match_key_bytes_4_T_1 ? phv_data_59 : _GEN_3125; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3127 = 8'h3c == _match_key_bytes_4_T_1 ? phv_data_60 : _GEN_3126; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3128 = 8'h3d == _match_key_bytes_4_T_1 ? phv_data_61 : _GEN_3127; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3129 = 8'h3e == _match_key_bytes_4_T_1 ? phv_data_62 : _GEN_3128; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3130 = 8'h3f == _match_key_bytes_4_T_1 ? phv_data_63 : _GEN_3129; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3131 = 8'h40 == _match_key_bytes_4_T_1 ? phv_data_64 : _GEN_3130; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3132 = 8'h41 == _match_key_bytes_4_T_1 ? phv_data_65 : _GEN_3131; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3133 = 8'h42 == _match_key_bytes_4_T_1 ? phv_data_66 : _GEN_3132; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3134 = 8'h43 == _match_key_bytes_4_T_1 ? phv_data_67 : _GEN_3133; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3135 = 8'h44 == _match_key_bytes_4_T_1 ? phv_data_68 : _GEN_3134; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3136 = 8'h45 == _match_key_bytes_4_T_1 ? phv_data_69 : _GEN_3135; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3137 = 8'h46 == _match_key_bytes_4_T_1 ? phv_data_70 : _GEN_3136; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3138 = 8'h47 == _match_key_bytes_4_T_1 ? phv_data_71 : _GEN_3137; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3139 = 8'h48 == _match_key_bytes_4_T_1 ? phv_data_72 : _GEN_3138; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3140 = 8'h49 == _match_key_bytes_4_T_1 ? phv_data_73 : _GEN_3139; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3141 = 8'h4a == _match_key_bytes_4_T_1 ? phv_data_74 : _GEN_3140; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3142 = 8'h4b == _match_key_bytes_4_T_1 ? phv_data_75 : _GEN_3141; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3143 = 8'h4c == _match_key_bytes_4_T_1 ? phv_data_76 : _GEN_3142; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3144 = 8'h4d == _match_key_bytes_4_T_1 ? phv_data_77 : _GEN_3143; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3145 = 8'h4e == _match_key_bytes_4_T_1 ? phv_data_78 : _GEN_3144; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3146 = 8'h4f == _match_key_bytes_4_T_1 ? phv_data_79 : _GEN_3145; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3147 = 8'h50 == _match_key_bytes_4_T_1 ? phv_data_80 : _GEN_3146; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3148 = 8'h51 == _match_key_bytes_4_T_1 ? phv_data_81 : _GEN_3147; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3149 = 8'h52 == _match_key_bytes_4_T_1 ? phv_data_82 : _GEN_3148; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3150 = 8'h53 == _match_key_bytes_4_T_1 ? phv_data_83 : _GEN_3149; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3151 = 8'h54 == _match_key_bytes_4_T_1 ? phv_data_84 : _GEN_3150; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3152 = 8'h55 == _match_key_bytes_4_T_1 ? phv_data_85 : _GEN_3151; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3153 = 8'h56 == _match_key_bytes_4_T_1 ? phv_data_86 : _GEN_3152; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3154 = 8'h57 == _match_key_bytes_4_T_1 ? phv_data_87 : _GEN_3153; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3155 = 8'h58 == _match_key_bytes_4_T_1 ? phv_data_88 : _GEN_3154; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3156 = 8'h59 == _match_key_bytes_4_T_1 ? phv_data_89 : _GEN_3155; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3157 = 8'h5a == _match_key_bytes_4_T_1 ? phv_data_90 : _GEN_3156; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3158 = 8'h5b == _match_key_bytes_4_T_1 ? phv_data_91 : _GEN_3157; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3159 = 8'h5c == _match_key_bytes_4_T_1 ? phv_data_92 : _GEN_3158; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3160 = 8'h5d == _match_key_bytes_4_T_1 ? phv_data_93 : _GEN_3159; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3161 = 8'h5e == _match_key_bytes_4_T_1 ? phv_data_94 : _GEN_3160; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3162 = 8'h5f == _match_key_bytes_4_T_1 ? phv_data_95 : _GEN_3161; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3163 = 8'h60 == _match_key_bytes_4_T_1 ? phv_data_96 : _GEN_3162; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3164 = 8'h61 == _match_key_bytes_4_T_1 ? phv_data_97 : _GEN_3163; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3165 = 8'h62 == _match_key_bytes_4_T_1 ? phv_data_98 : _GEN_3164; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3166 = 8'h63 == _match_key_bytes_4_T_1 ? phv_data_99 : _GEN_3165; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3167 = 8'h64 == _match_key_bytes_4_T_1 ? phv_data_100 : _GEN_3166; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3168 = 8'h65 == _match_key_bytes_4_T_1 ? phv_data_101 : _GEN_3167; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3169 = 8'h66 == _match_key_bytes_4_T_1 ? phv_data_102 : _GEN_3168; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3170 = 8'h67 == _match_key_bytes_4_T_1 ? phv_data_103 : _GEN_3169; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3171 = 8'h68 == _match_key_bytes_4_T_1 ? phv_data_104 : _GEN_3170; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3172 = 8'h69 == _match_key_bytes_4_T_1 ? phv_data_105 : _GEN_3171; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3173 = 8'h6a == _match_key_bytes_4_T_1 ? phv_data_106 : _GEN_3172; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3174 = 8'h6b == _match_key_bytes_4_T_1 ? phv_data_107 : _GEN_3173; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3175 = 8'h6c == _match_key_bytes_4_T_1 ? phv_data_108 : _GEN_3174; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3176 = 8'h6d == _match_key_bytes_4_T_1 ? phv_data_109 : _GEN_3175; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3177 = 8'h6e == _match_key_bytes_4_T_1 ? phv_data_110 : _GEN_3176; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3178 = 8'h6f == _match_key_bytes_4_T_1 ? phv_data_111 : _GEN_3177; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3179 = 8'h70 == _match_key_bytes_4_T_1 ? phv_data_112 : _GEN_3178; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3180 = 8'h71 == _match_key_bytes_4_T_1 ? phv_data_113 : _GEN_3179; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3181 = 8'h72 == _match_key_bytes_4_T_1 ? phv_data_114 : _GEN_3180; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3182 = 8'h73 == _match_key_bytes_4_T_1 ? phv_data_115 : _GEN_3181; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3183 = 8'h74 == _match_key_bytes_4_T_1 ? phv_data_116 : _GEN_3182; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3184 = 8'h75 == _match_key_bytes_4_T_1 ? phv_data_117 : _GEN_3183; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3185 = 8'h76 == _match_key_bytes_4_T_1 ? phv_data_118 : _GEN_3184; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3186 = 8'h77 == _match_key_bytes_4_T_1 ? phv_data_119 : _GEN_3185; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3187 = 8'h78 == _match_key_bytes_4_T_1 ? phv_data_120 : _GEN_3186; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3188 = 8'h79 == _match_key_bytes_4_T_1 ? phv_data_121 : _GEN_3187; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3189 = 8'h7a == _match_key_bytes_4_T_1 ? phv_data_122 : _GEN_3188; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3190 = 8'h7b == _match_key_bytes_4_T_1 ? phv_data_123 : _GEN_3189; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3191 = 8'h7c == _match_key_bytes_4_T_1 ? phv_data_124 : _GEN_3190; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3192 = 8'h7d == _match_key_bytes_4_T_1 ? phv_data_125 : _GEN_3191; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3193 = 8'h7e == _match_key_bytes_4_T_1 ? phv_data_126 : _GEN_3192; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3194 = 8'h7f == _match_key_bytes_4_T_1 ? phv_data_127 : _GEN_3193; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3195 = 8'h80 == _match_key_bytes_4_T_1 ? phv_data_128 : _GEN_3194; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3196 = 8'h81 == _match_key_bytes_4_T_1 ? phv_data_129 : _GEN_3195; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3197 = 8'h82 == _match_key_bytes_4_T_1 ? phv_data_130 : _GEN_3196; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3198 = 8'h83 == _match_key_bytes_4_T_1 ? phv_data_131 : _GEN_3197; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3199 = 8'h84 == _match_key_bytes_4_T_1 ? phv_data_132 : _GEN_3198; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3200 = 8'h85 == _match_key_bytes_4_T_1 ? phv_data_133 : _GEN_3199; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3201 = 8'h86 == _match_key_bytes_4_T_1 ? phv_data_134 : _GEN_3200; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3202 = 8'h87 == _match_key_bytes_4_T_1 ? phv_data_135 : _GEN_3201; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3203 = 8'h88 == _match_key_bytes_4_T_1 ? phv_data_136 : _GEN_3202; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3204 = 8'h89 == _match_key_bytes_4_T_1 ? phv_data_137 : _GEN_3203; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3205 = 8'h8a == _match_key_bytes_4_T_1 ? phv_data_138 : _GEN_3204; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3206 = 8'h8b == _match_key_bytes_4_T_1 ? phv_data_139 : _GEN_3205; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3207 = 8'h8c == _match_key_bytes_4_T_1 ? phv_data_140 : _GEN_3206; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3208 = 8'h8d == _match_key_bytes_4_T_1 ? phv_data_141 : _GEN_3207; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3209 = 8'h8e == _match_key_bytes_4_T_1 ? phv_data_142 : _GEN_3208; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3210 = 8'h8f == _match_key_bytes_4_T_1 ? phv_data_143 : _GEN_3209; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3211 = 8'h90 == _match_key_bytes_4_T_1 ? phv_data_144 : _GEN_3210; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3212 = 8'h91 == _match_key_bytes_4_T_1 ? phv_data_145 : _GEN_3211; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3213 = 8'h92 == _match_key_bytes_4_T_1 ? phv_data_146 : _GEN_3212; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3214 = 8'h93 == _match_key_bytes_4_T_1 ? phv_data_147 : _GEN_3213; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3215 = 8'h94 == _match_key_bytes_4_T_1 ? phv_data_148 : _GEN_3214; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3216 = 8'h95 == _match_key_bytes_4_T_1 ? phv_data_149 : _GEN_3215; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3217 = 8'h96 == _match_key_bytes_4_T_1 ? phv_data_150 : _GEN_3216; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3218 = 8'h97 == _match_key_bytes_4_T_1 ? phv_data_151 : _GEN_3217; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3219 = 8'h98 == _match_key_bytes_4_T_1 ? phv_data_152 : _GEN_3218; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3220 = 8'h99 == _match_key_bytes_4_T_1 ? phv_data_153 : _GEN_3219; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3221 = 8'h9a == _match_key_bytes_4_T_1 ? phv_data_154 : _GEN_3220; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3222 = 8'h9b == _match_key_bytes_4_T_1 ? phv_data_155 : _GEN_3221; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3223 = 8'h9c == _match_key_bytes_4_T_1 ? phv_data_156 : _GEN_3222; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3224 = 8'h9d == _match_key_bytes_4_T_1 ? phv_data_157 : _GEN_3223; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3225 = 8'h9e == _match_key_bytes_4_T_1 ? phv_data_158 : _GEN_3224; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3226 = 8'h9f == _match_key_bytes_4_T_1 ? phv_data_159 : _GEN_3225; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_4 = 8'h13 < _GEN_6 ? _GEN_3226 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_3_T_1 = key_offset + 8'h14; // @[matcher.scala 72:98]
  wire [7:0] _GEN_3229 = 8'h1 == _match_key_bytes_3_T_1 ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3230 = 8'h2 == _match_key_bytes_3_T_1 ? phv_data_2 : _GEN_3229; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3231 = 8'h3 == _match_key_bytes_3_T_1 ? phv_data_3 : _GEN_3230; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3232 = 8'h4 == _match_key_bytes_3_T_1 ? phv_data_4 : _GEN_3231; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3233 = 8'h5 == _match_key_bytes_3_T_1 ? phv_data_5 : _GEN_3232; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3234 = 8'h6 == _match_key_bytes_3_T_1 ? phv_data_6 : _GEN_3233; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3235 = 8'h7 == _match_key_bytes_3_T_1 ? phv_data_7 : _GEN_3234; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3236 = 8'h8 == _match_key_bytes_3_T_1 ? phv_data_8 : _GEN_3235; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3237 = 8'h9 == _match_key_bytes_3_T_1 ? phv_data_9 : _GEN_3236; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3238 = 8'ha == _match_key_bytes_3_T_1 ? phv_data_10 : _GEN_3237; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3239 = 8'hb == _match_key_bytes_3_T_1 ? phv_data_11 : _GEN_3238; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3240 = 8'hc == _match_key_bytes_3_T_1 ? phv_data_12 : _GEN_3239; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3241 = 8'hd == _match_key_bytes_3_T_1 ? phv_data_13 : _GEN_3240; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3242 = 8'he == _match_key_bytes_3_T_1 ? phv_data_14 : _GEN_3241; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3243 = 8'hf == _match_key_bytes_3_T_1 ? phv_data_15 : _GEN_3242; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3244 = 8'h10 == _match_key_bytes_3_T_1 ? phv_data_16 : _GEN_3243; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3245 = 8'h11 == _match_key_bytes_3_T_1 ? phv_data_17 : _GEN_3244; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3246 = 8'h12 == _match_key_bytes_3_T_1 ? phv_data_18 : _GEN_3245; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3247 = 8'h13 == _match_key_bytes_3_T_1 ? phv_data_19 : _GEN_3246; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3248 = 8'h14 == _match_key_bytes_3_T_1 ? phv_data_20 : _GEN_3247; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3249 = 8'h15 == _match_key_bytes_3_T_1 ? phv_data_21 : _GEN_3248; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3250 = 8'h16 == _match_key_bytes_3_T_1 ? phv_data_22 : _GEN_3249; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3251 = 8'h17 == _match_key_bytes_3_T_1 ? phv_data_23 : _GEN_3250; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3252 = 8'h18 == _match_key_bytes_3_T_1 ? phv_data_24 : _GEN_3251; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3253 = 8'h19 == _match_key_bytes_3_T_1 ? phv_data_25 : _GEN_3252; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3254 = 8'h1a == _match_key_bytes_3_T_1 ? phv_data_26 : _GEN_3253; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3255 = 8'h1b == _match_key_bytes_3_T_1 ? phv_data_27 : _GEN_3254; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3256 = 8'h1c == _match_key_bytes_3_T_1 ? phv_data_28 : _GEN_3255; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3257 = 8'h1d == _match_key_bytes_3_T_1 ? phv_data_29 : _GEN_3256; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3258 = 8'h1e == _match_key_bytes_3_T_1 ? phv_data_30 : _GEN_3257; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3259 = 8'h1f == _match_key_bytes_3_T_1 ? phv_data_31 : _GEN_3258; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3260 = 8'h20 == _match_key_bytes_3_T_1 ? phv_data_32 : _GEN_3259; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3261 = 8'h21 == _match_key_bytes_3_T_1 ? phv_data_33 : _GEN_3260; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3262 = 8'h22 == _match_key_bytes_3_T_1 ? phv_data_34 : _GEN_3261; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3263 = 8'h23 == _match_key_bytes_3_T_1 ? phv_data_35 : _GEN_3262; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3264 = 8'h24 == _match_key_bytes_3_T_1 ? phv_data_36 : _GEN_3263; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3265 = 8'h25 == _match_key_bytes_3_T_1 ? phv_data_37 : _GEN_3264; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3266 = 8'h26 == _match_key_bytes_3_T_1 ? phv_data_38 : _GEN_3265; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3267 = 8'h27 == _match_key_bytes_3_T_1 ? phv_data_39 : _GEN_3266; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3268 = 8'h28 == _match_key_bytes_3_T_1 ? phv_data_40 : _GEN_3267; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3269 = 8'h29 == _match_key_bytes_3_T_1 ? phv_data_41 : _GEN_3268; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3270 = 8'h2a == _match_key_bytes_3_T_1 ? phv_data_42 : _GEN_3269; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3271 = 8'h2b == _match_key_bytes_3_T_1 ? phv_data_43 : _GEN_3270; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3272 = 8'h2c == _match_key_bytes_3_T_1 ? phv_data_44 : _GEN_3271; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3273 = 8'h2d == _match_key_bytes_3_T_1 ? phv_data_45 : _GEN_3272; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3274 = 8'h2e == _match_key_bytes_3_T_1 ? phv_data_46 : _GEN_3273; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3275 = 8'h2f == _match_key_bytes_3_T_1 ? phv_data_47 : _GEN_3274; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3276 = 8'h30 == _match_key_bytes_3_T_1 ? phv_data_48 : _GEN_3275; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3277 = 8'h31 == _match_key_bytes_3_T_1 ? phv_data_49 : _GEN_3276; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3278 = 8'h32 == _match_key_bytes_3_T_1 ? phv_data_50 : _GEN_3277; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3279 = 8'h33 == _match_key_bytes_3_T_1 ? phv_data_51 : _GEN_3278; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3280 = 8'h34 == _match_key_bytes_3_T_1 ? phv_data_52 : _GEN_3279; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3281 = 8'h35 == _match_key_bytes_3_T_1 ? phv_data_53 : _GEN_3280; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3282 = 8'h36 == _match_key_bytes_3_T_1 ? phv_data_54 : _GEN_3281; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3283 = 8'h37 == _match_key_bytes_3_T_1 ? phv_data_55 : _GEN_3282; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3284 = 8'h38 == _match_key_bytes_3_T_1 ? phv_data_56 : _GEN_3283; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3285 = 8'h39 == _match_key_bytes_3_T_1 ? phv_data_57 : _GEN_3284; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3286 = 8'h3a == _match_key_bytes_3_T_1 ? phv_data_58 : _GEN_3285; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3287 = 8'h3b == _match_key_bytes_3_T_1 ? phv_data_59 : _GEN_3286; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3288 = 8'h3c == _match_key_bytes_3_T_1 ? phv_data_60 : _GEN_3287; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3289 = 8'h3d == _match_key_bytes_3_T_1 ? phv_data_61 : _GEN_3288; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3290 = 8'h3e == _match_key_bytes_3_T_1 ? phv_data_62 : _GEN_3289; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3291 = 8'h3f == _match_key_bytes_3_T_1 ? phv_data_63 : _GEN_3290; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3292 = 8'h40 == _match_key_bytes_3_T_1 ? phv_data_64 : _GEN_3291; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3293 = 8'h41 == _match_key_bytes_3_T_1 ? phv_data_65 : _GEN_3292; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3294 = 8'h42 == _match_key_bytes_3_T_1 ? phv_data_66 : _GEN_3293; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3295 = 8'h43 == _match_key_bytes_3_T_1 ? phv_data_67 : _GEN_3294; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3296 = 8'h44 == _match_key_bytes_3_T_1 ? phv_data_68 : _GEN_3295; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3297 = 8'h45 == _match_key_bytes_3_T_1 ? phv_data_69 : _GEN_3296; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3298 = 8'h46 == _match_key_bytes_3_T_1 ? phv_data_70 : _GEN_3297; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3299 = 8'h47 == _match_key_bytes_3_T_1 ? phv_data_71 : _GEN_3298; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3300 = 8'h48 == _match_key_bytes_3_T_1 ? phv_data_72 : _GEN_3299; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3301 = 8'h49 == _match_key_bytes_3_T_1 ? phv_data_73 : _GEN_3300; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3302 = 8'h4a == _match_key_bytes_3_T_1 ? phv_data_74 : _GEN_3301; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3303 = 8'h4b == _match_key_bytes_3_T_1 ? phv_data_75 : _GEN_3302; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3304 = 8'h4c == _match_key_bytes_3_T_1 ? phv_data_76 : _GEN_3303; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3305 = 8'h4d == _match_key_bytes_3_T_1 ? phv_data_77 : _GEN_3304; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3306 = 8'h4e == _match_key_bytes_3_T_1 ? phv_data_78 : _GEN_3305; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3307 = 8'h4f == _match_key_bytes_3_T_1 ? phv_data_79 : _GEN_3306; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3308 = 8'h50 == _match_key_bytes_3_T_1 ? phv_data_80 : _GEN_3307; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3309 = 8'h51 == _match_key_bytes_3_T_1 ? phv_data_81 : _GEN_3308; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3310 = 8'h52 == _match_key_bytes_3_T_1 ? phv_data_82 : _GEN_3309; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3311 = 8'h53 == _match_key_bytes_3_T_1 ? phv_data_83 : _GEN_3310; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3312 = 8'h54 == _match_key_bytes_3_T_1 ? phv_data_84 : _GEN_3311; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3313 = 8'h55 == _match_key_bytes_3_T_1 ? phv_data_85 : _GEN_3312; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3314 = 8'h56 == _match_key_bytes_3_T_1 ? phv_data_86 : _GEN_3313; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3315 = 8'h57 == _match_key_bytes_3_T_1 ? phv_data_87 : _GEN_3314; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3316 = 8'h58 == _match_key_bytes_3_T_1 ? phv_data_88 : _GEN_3315; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3317 = 8'h59 == _match_key_bytes_3_T_1 ? phv_data_89 : _GEN_3316; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3318 = 8'h5a == _match_key_bytes_3_T_1 ? phv_data_90 : _GEN_3317; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3319 = 8'h5b == _match_key_bytes_3_T_1 ? phv_data_91 : _GEN_3318; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3320 = 8'h5c == _match_key_bytes_3_T_1 ? phv_data_92 : _GEN_3319; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3321 = 8'h5d == _match_key_bytes_3_T_1 ? phv_data_93 : _GEN_3320; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3322 = 8'h5e == _match_key_bytes_3_T_1 ? phv_data_94 : _GEN_3321; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3323 = 8'h5f == _match_key_bytes_3_T_1 ? phv_data_95 : _GEN_3322; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3324 = 8'h60 == _match_key_bytes_3_T_1 ? phv_data_96 : _GEN_3323; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3325 = 8'h61 == _match_key_bytes_3_T_1 ? phv_data_97 : _GEN_3324; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3326 = 8'h62 == _match_key_bytes_3_T_1 ? phv_data_98 : _GEN_3325; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3327 = 8'h63 == _match_key_bytes_3_T_1 ? phv_data_99 : _GEN_3326; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3328 = 8'h64 == _match_key_bytes_3_T_1 ? phv_data_100 : _GEN_3327; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3329 = 8'h65 == _match_key_bytes_3_T_1 ? phv_data_101 : _GEN_3328; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3330 = 8'h66 == _match_key_bytes_3_T_1 ? phv_data_102 : _GEN_3329; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3331 = 8'h67 == _match_key_bytes_3_T_1 ? phv_data_103 : _GEN_3330; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3332 = 8'h68 == _match_key_bytes_3_T_1 ? phv_data_104 : _GEN_3331; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3333 = 8'h69 == _match_key_bytes_3_T_1 ? phv_data_105 : _GEN_3332; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3334 = 8'h6a == _match_key_bytes_3_T_1 ? phv_data_106 : _GEN_3333; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3335 = 8'h6b == _match_key_bytes_3_T_1 ? phv_data_107 : _GEN_3334; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3336 = 8'h6c == _match_key_bytes_3_T_1 ? phv_data_108 : _GEN_3335; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3337 = 8'h6d == _match_key_bytes_3_T_1 ? phv_data_109 : _GEN_3336; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3338 = 8'h6e == _match_key_bytes_3_T_1 ? phv_data_110 : _GEN_3337; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3339 = 8'h6f == _match_key_bytes_3_T_1 ? phv_data_111 : _GEN_3338; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3340 = 8'h70 == _match_key_bytes_3_T_1 ? phv_data_112 : _GEN_3339; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3341 = 8'h71 == _match_key_bytes_3_T_1 ? phv_data_113 : _GEN_3340; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3342 = 8'h72 == _match_key_bytes_3_T_1 ? phv_data_114 : _GEN_3341; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3343 = 8'h73 == _match_key_bytes_3_T_1 ? phv_data_115 : _GEN_3342; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3344 = 8'h74 == _match_key_bytes_3_T_1 ? phv_data_116 : _GEN_3343; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3345 = 8'h75 == _match_key_bytes_3_T_1 ? phv_data_117 : _GEN_3344; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3346 = 8'h76 == _match_key_bytes_3_T_1 ? phv_data_118 : _GEN_3345; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3347 = 8'h77 == _match_key_bytes_3_T_1 ? phv_data_119 : _GEN_3346; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3348 = 8'h78 == _match_key_bytes_3_T_1 ? phv_data_120 : _GEN_3347; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3349 = 8'h79 == _match_key_bytes_3_T_1 ? phv_data_121 : _GEN_3348; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3350 = 8'h7a == _match_key_bytes_3_T_1 ? phv_data_122 : _GEN_3349; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3351 = 8'h7b == _match_key_bytes_3_T_1 ? phv_data_123 : _GEN_3350; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3352 = 8'h7c == _match_key_bytes_3_T_1 ? phv_data_124 : _GEN_3351; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3353 = 8'h7d == _match_key_bytes_3_T_1 ? phv_data_125 : _GEN_3352; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3354 = 8'h7e == _match_key_bytes_3_T_1 ? phv_data_126 : _GEN_3353; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3355 = 8'h7f == _match_key_bytes_3_T_1 ? phv_data_127 : _GEN_3354; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3356 = 8'h80 == _match_key_bytes_3_T_1 ? phv_data_128 : _GEN_3355; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3357 = 8'h81 == _match_key_bytes_3_T_1 ? phv_data_129 : _GEN_3356; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3358 = 8'h82 == _match_key_bytes_3_T_1 ? phv_data_130 : _GEN_3357; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3359 = 8'h83 == _match_key_bytes_3_T_1 ? phv_data_131 : _GEN_3358; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3360 = 8'h84 == _match_key_bytes_3_T_1 ? phv_data_132 : _GEN_3359; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3361 = 8'h85 == _match_key_bytes_3_T_1 ? phv_data_133 : _GEN_3360; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3362 = 8'h86 == _match_key_bytes_3_T_1 ? phv_data_134 : _GEN_3361; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3363 = 8'h87 == _match_key_bytes_3_T_1 ? phv_data_135 : _GEN_3362; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3364 = 8'h88 == _match_key_bytes_3_T_1 ? phv_data_136 : _GEN_3363; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3365 = 8'h89 == _match_key_bytes_3_T_1 ? phv_data_137 : _GEN_3364; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3366 = 8'h8a == _match_key_bytes_3_T_1 ? phv_data_138 : _GEN_3365; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3367 = 8'h8b == _match_key_bytes_3_T_1 ? phv_data_139 : _GEN_3366; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3368 = 8'h8c == _match_key_bytes_3_T_1 ? phv_data_140 : _GEN_3367; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3369 = 8'h8d == _match_key_bytes_3_T_1 ? phv_data_141 : _GEN_3368; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3370 = 8'h8e == _match_key_bytes_3_T_1 ? phv_data_142 : _GEN_3369; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3371 = 8'h8f == _match_key_bytes_3_T_1 ? phv_data_143 : _GEN_3370; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3372 = 8'h90 == _match_key_bytes_3_T_1 ? phv_data_144 : _GEN_3371; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3373 = 8'h91 == _match_key_bytes_3_T_1 ? phv_data_145 : _GEN_3372; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3374 = 8'h92 == _match_key_bytes_3_T_1 ? phv_data_146 : _GEN_3373; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3375 = 8'h93 == _match_key_bytes_3_T_1 ? phv_data_147 : _GEN_3374; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3376 = 8'h94 == _match_key_bytes_3_T_1 ? phv_data_148 : _GEN_3375; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3377 = 8'h95 == _match_key_bytes_3_T_1 ? phv_data_149 : _GEN_3376; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3378 = 8'h96 == _match_key_bytes_3_T_1 ? phv_data_150 : _GEN_3377; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3379 = 8'h97 == _match_key_bytes_3_T_1 ? phv_data_151 : _GEN_3378; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3380 = 8'h98 == _match_key_bytes_3_T_1 ? phv_data_152 : _GEN_3379; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3381 = 8'h99 == _match_key_bytes_3_T_1 ? phv_data_153 : _GEN_3380; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3382 = 8'h9a == _match_key_bytes_3_T_1 ? phv_data_154 : _GEN_3381; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3383 = 8'h9b == _match_key_bytes_3_T_1 ? phv_data_155 : _GEN_3382; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3384 = 8'h9c == _match_key_bytes_3_T_1 ? phv_data_156 : _GEN_3383; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3385 = 8'h9d == _match_key_bytes_3_T_1 ? phv_data_157 : _GEN_3384; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3386 = 8'h9e == _match_key_bytes_3_T_1 ? phv_data_158 : _GEN_3385; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3387 = 8'h9f == _match_key_bytes_3_T_1 ? phv_data_159 : _GEN_3386; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_3 = 8'h14 < _GEN_6 ? _GEN_3387 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_2_T_1 = key_offset + 8'h15; // @[matcher.scala 72:98]
  wire [7:0] _GEN_3390 = 8'h1 == _match_key_bytes_2_T_1 ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3391 = 8'h2 == _match_key_bytes_2_T_1 ? phv_data_2 : _GEN_3390; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3392 = 8'h3 == _match_key_bytes_2_T_1 ? phv_data_3 : _GEN_3391; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3393 = 8'h4 == _match_key_bytes_2_T_1 ? phv_data_4 : _GEN_3392; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3394 = 8'h5 == _match_key_bytes_2_T_1 ? phv_data_5 : _GEN_3393; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3395 = 8'h6 == _match_key_bytes_2_T_1 ? phv_data_6 : _GEN_3394; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3396 = 8'h7 == _match_key_bytes_2_T_1 ? phv_data_7 : _GEN_3395; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3397 = 8'h8 == _match_key_bytes_2_T_1 ? phv_data_8 : _GEN_3396; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3398 = 8'h9 == _match_key_bytes_2_T_1 ? phv_data_9 : _GEN_3397; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3399 = 8'ha == _match_key_bytes_2_T_1 ? phv_data_10 : _GEN_3398; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3400 = 8'hb == _match_key_bytes_2_T_1 ? phv_data_11 : _GEN_3399; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3401 = 8'hc == _match_key_bytes_2_T_1 ? phv_data_12 : _GEN_3400; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3402 = 8'hd == _match_key_bytes_2_T_1 ? phv_data_13 : _GEN_3401; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3403 = 8'he == _match_key_bytes_2_T_1 ? phv_data_14 : _GEN_3402; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3404 = 8'hf == _match_key_bytes_2_T_1 ? phv_data_15 : _GEN_3403; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3405 = 8'h10 == _match_key_bytes_2_T_1 ? phv_data_16 : _GEN_3404; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3406 = 8'h11 == _match_key_bytes_2_T_1 ? phv_data_17 : _GEN_3405; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3407 = 8'h12 == _match_key_bytes_2_T_1 ? phv_data_18 : _GEN_3406; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3408 = 8'h13 == _match_key_bytes_2_T_1 ? phv_data_19 : _GEN_3407; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3409 = 8'h14 == _match_key_bytes_2_T_1 ? phv_data_20 : _GEN_3408; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3410 = 8'h15 == _match_key_bytes_2_T_1 ? phv_data_21 : _GEN_3409; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3411 = 8'h16 == _match_key_bytes_2_T_1 ? phv_data_22 : _GEN_3410; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3412 = 8'h17 == _match_key_bytes_2_T_1 ? phv_data_23 : _GEN_3411; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3413 = 8'h18 == _match_key_bytes_2_T_1 ? phv_data_24 : _GEN_3412; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3414 = 8'h19 == _match_key_bytes_2_T_1 ? phv_data_25 : _GEN_3413; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3415 = 8'h1a == _match_key_bytes_2_T_1 ? phv_data_26 : _GEN_3414; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3416 = 8'h1b == _match_key_bytes_2_T_1 ? phv_data_27 : _GEN_3415; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3417 = 8'h1c == _match_key_bytes_2_T_1 ? phv_data_28 : _GEN_3416; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3418 = 8'h1d == _match_key_bytes_2_T_1 ? phv_data_29 : _GEN_3417; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3419 = 8'h1e == _match_key_bytes_2_T_1 ? phv_data_30 : _GEN_3418; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3420 = 8'h1f == _match_key_bytes_2_T_1 ? phv_data_31 : _GEN_3419; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3421 = 8'h20 == _match_key_bytes_2_T_1 ? phv_data_32 : _GEN_3420; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3422 = 8'h21 == _match_key_bytes_2_T_1 ? phv_data_33 : _GEN_3421; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3423 = 8'h22 == _match_key_bytes_2_T_1 ? phv_data_34 : _GEN_3422; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3424 = 8'h23 == _match_key_bytes_2_T_1 ? phv_data_35 : _GEN_3423; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3425 = 8'h24 == _match_key_bytes_2_T_1 ? phv_data_36 : _GEN_3424; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3426 = 8'h25 == _match_key_bytes_2_T_1 ? phv_data_37 : _GEN_3425; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3427 = 8'h26 == _match_key_bytes_2_T_1 ? phv_data_38 : _GEN_3426; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3428 = 8'h27 == _match_key_bytes_2_T_1 ? phv_data_39 : _GEN_3427; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3429 = 8'h28 == _match_key_bytes_2_T_1 ? phv_data_40 : _GEN_3428; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3430 = 8'h29 == _match_key_bytes_2_T_1 ? phv_data_41 : _GEN_3429; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3431 = 8'h2a == _match_key_bytes_2_T_1 ? phv_data_42 : _GEN_3430; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3432 = 8'h2b == _match_key_bytes_2_T_1 ? phv_data_43 : _GEN_3431; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3433 = 8'h2c == _match_key_bytes_2_T_1 ? phv_data_44 : _GEN_3432; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3434 = 8'h2d == _match_key_bytes_2_T_1 ? phv_data_45 : _GEN_3433; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3435 = 8'h2e == _match_key_bytes_2_T_1 ? phv_data_46 : _GEN_3434; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3436 = 8'h2f == _match_key_bytes_2_T_1 ? phv_data_47 : _GEN_3435; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3437 = 8'h30 == _match_key_bytes_2_T_1 ? phv_data_48 : _GEN_3436; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3438 = 8'h31 == _match_key_bytes_2_T_1 ? phv_data_49 : _GEN_3437; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3439 = 8'h32 == _match_key_bytes_2_T_1 ? phv_data_50 : _GEN_3438; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3440 = 8'h33 == _match_key_bytes_2_T_1 ? phv_data_51 : _GEN_3439; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3441 = 8'h34 == _match_key_bytes_2_T_1 ? phv_data_52 : _GEN_3440; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3442 = 8'h35 == _match_key_bytes_2_T_1 ? phv_data_53 : _GEN_3441; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3443 = 8'h36 == _match_key_bytes_2_T_1 ? phv_data_54 : _GEN_3442; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3444 = 8'h37 == _match_key_bytes_2_T_1 ? phv_data_55 : _GEN_3443; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3445 = 8'h38 == _match_key_bytes_2_T_1 ? phv_data_56 : _GEN_3444; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3446 = 8'h39 == _match_key_bytes_2_T_1 ? phv_data_57 : _GEN_3445; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3447 = 8'h3a == _match_key_bytes_2_T_1 ? phv_data_58 : _GEN_3446; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3448 = 8'h3b == _match_key_bytes_2_T_1 ? phv_data_59 : _GEN_3447; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3449 = 8'h3c == _match_key_bytes_2_T_1 ? phv_data_60 : _GEN_3448; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3450 = 8'h3d == _match_key_bytes_2_T_1 ? phv_data_61 : _GEN_3449; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3451 = 8'h3e == _match_key_bytes_2_T_1 ? phv_data_62 : _GEN_3450; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3452 = 8'h3f == _match_key_bytes_2_T_1 ? phv_data_63 : _GEN_3451; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3453 = 8'h40 == _match_key_bytes_2_T_1 ? phv_data_64 : _GEN_3452; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3454 = 8'h41 == _match_key_bytes_2_T_1 ? phv_data_65 : _GEN_3453; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3455 = 8'h42 == _match_key_bytes_2_T_1 ? phv_data_66 : _GEN_3454; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3456 = 8'h43 == _match_key_bytes_2_T_1 ? phv_data_67 : _GEN_3455; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3457 = 8'h44 == _match_key_bytes_2_T_1 ? phv_data_68 : _GEN_3456; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3458 = 8'h45 == _match_key_bytes_2_T_1 ? phv_data_69 : _GEN_3457; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3459 = 8'h46 == _match_key_bytes_2_T_1 ? phv_data_70 : _GEN_3458; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3460 = 8'h47 == _match_key_bytes_2_T_1 ? phv_data_71 : _GEN_3459; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3461 = 8'h48 == _match_key_bytes_2_T_1 ? phv_data_72 : _GEN_3460; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3462 = 8'h49 == _match_key_bytes_2_T_1 ? phv_data_73 : _GEN_3461; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3463 = 8'h4a == _match_key_bytes_2_T_1 ? phv_data_74 : _GEN_3462; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3464 = 8'h4b == _match_key_bytes_2_T_1 ? phv_data_75 : _GEN_3463; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3465 = 8'h4c == _match_key_bytes_2_T_1 ? phv_data_76 : _GEN_3464; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3466 = 8'h4d == _match_key_bytes_2_T_1 ? phv_data_77 : _GEN_3465; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3467 = 8'h4e == _match_key_bytes_2_T_1 ? phv_data_78 : _GEN_3466; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3468 = 8'h4f == _match_key_bytes_2_T_1 ? phv_data_79 : _GEN_3467; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3469 = 8'h50 == _match_key_bytes_2_T_1 ? phv_data_80 : _GEN_3468; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3470 = 8'h51 == _match_key_bytes_2_T_1 ? phv_data_81 : _GEN_3469; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3471 = 8'h52 == _match_key_bytes_2_T_1 ? phv_data_82 : _GEN_3470; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3472 = 8'h53 == _match_key_bytes_2_T_1 ? phv_data_83 : _GEN_3471; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3473 = 8'h54 == _match_key_bytes_2_T_1 ? phv_data_84 : _GEN_3472; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3474 = 8'h55 == _match_key_bytes_2_T_1 ? phv_data_85 : _GEN_3473; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3475 = 8'h56 == _match_key_bytes_2_T_1 ? phv_data_86 : _GEN_3474; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3476 = 8'h57 == _match_key_bytes_2_T_1 ? phv_data_87 : _GEN_3475; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3477 = 8'h58 == _match_key_bytes_2_T_1 ? phv_data_88 : _GEN_3476; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3478 = 8'h59 == _match_key_bytes_2_T_1 ? phv_data_89 : _GEN_3477; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3479 = 8'h5a == _match_key_bytes_2_T_1 ? phv_data_90 : _GEN_3478; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3480 = 8'h5b == _match_key_bytes_2_T_1 ? phv_data_91 : _GEN_3479; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3481 = 8'h5c == _match_key_bytes_2_T_1 ? phv_data_92 : _GEN_3480; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3482 = 8'h5d == _match_key_bytes_2_T_1 ? phv_data_93 : _GEN_3481; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3483 = 8'h5e == _match_key_bytes_2_T_1 ? phv_data_94 : _GEN_3482; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3484 = 8'h5f == _match_key_bytes_2_T_1 ? phv_data_95 : _GEN_3483; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3485 = 8'h60 == _match_key_bytes_2_T_1 ? phv_data_96 : _GEN_3484; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3486 = 8'h61 == _match_key_bytes_2_T_1 ? phv_data_97 : _GEN_3485; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3487 = 8'h62 == _match_key_bytes_2_T_1 ? phv_data_98 : _GEN_3486; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3488 = 8'h63 == _match_key_bytes_2_T_1 ? phv_data_99 : _GEN_3487; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3489 = 8'h64 == _match_key_bytes_2_T_1 ? phv_data_100 : _GEN_3488; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3490 = 8'h65 == _match_key_bytes_2_T_1 ? phv_data_101 : _GEN_3489; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3491 = 8'h66 == _match_key_bytes_2_T_1 ? phv_data_102 : _GEN_3490; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3492 = 8'h67 == _match_key_bytes_2_T_1 ? phv_data_103 : _GEN_3491; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3493 = 8'h68 == _match_key_bytes_2_T_1 ? phv_data_104 : _GEN_3492; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3494 = 8'h69 == _match_key_bytes_2_T_1 ? phv_data_105 : _GEN_3493; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3495 = 8'h6a == _match_key_bytes_2_T_1 ? phv_data_106 : _GEN_3494; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3496 = 8'h6b == _match_key_bytes_2_T_1 ? phv_data_107 : _GEN_3495; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3497 = 8'h6c == _match_key_bytes_2_T_1 ? phv_data_108 : _GEN_3496; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3498 = 8'h6d == _match_key_bytes_2_T_1 ? phv_data_109 : _GEN_3497; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3499 = 8'h6e == _match_key_bytes_2_T_1 ? phv_data_110 : _GEN_3498; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3500 = 8'h6f == _match_key_bytes_2_T_1 ? phv_data_111 : _GEN_3499; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3501 = 8'h70 == _match_key_bytes_2_T_1 ? phv_data_112 : _GEN_3500; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3502 = 8'h71 == _match_key_bytes_2_T_1 ? phv_data_113 : _GEN_3501; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3503 = 8'h72 == _match_key_bytes_2_T_1 ? phv_data_114 : _GEN_3502; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3504 = 8'h73 == _match_key_bytes_2_T_1 ? phv_data_115 : _GEN_3503; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3505 = 8'h74 == _match_key_bytes_2_T_1 ? phv_data_116 : _GEN_3504; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3506 = 8'h75 == _match_key_bytes_2_T_1 ? phv_data_117 : _GEN_3505; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3507 = 8'h76 == _match_key_bytes_2_T_1 ? phv_data_118 : _GEN_3506; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3508 = 8'h77 == _match_key_bytes_2_T_1 ? phv_data_119 : _GEN_3507; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3509 = 8'h78 == _match_key_bytes_2_T_1 ? phv_data_120 : _GEN_3508; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3510 = 8'h79 == _match_key_bytes_2_T_1 ? phv_data_121 : _GEN_3509; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3511 = 8'h7a == _match_key_bytes_2_T_1 ? phv_data_122 : _GEN_3510; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3512 = 8'h7b == _match_key_bytes_2_T_1 ? phv_data_123 : _GEN_3511; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3513 = 8'h7c == _match_key_bytes_2_T_1 ? phv_data_124 : _GEN_3512; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3514 = 8'h7d == _match_key_bytes_2_T_1 ? phv_data_125 : _GEN_3513; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3515 = 8'h7e == _match_key_bytes_2_T_1 ? phv_data_126 : _GEN_3514; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3516 = 8'h7f == _match_key_bytes_2_T_1 ? phv_data_127 : _GEN_3515; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3517 = 8'h80 == _match_key_bytes_2_T_1 ? phv_data_128 : _GEN_3516; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3518 = 8'h81 == _match_key_bytes_2_T_1 ? phv_data_129 : _GEN_3517; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3519 = 8'h82 == _match_key_bytes_2_T_1 ? phv_data_130 : _GEN_3518; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3520 = 8'h83 == _match_key_bytes_2_T_1 ? phv_data_131 : _GEN_3519; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3521 = 8'h84 == _match_key_bytes_2_T_1 ? phv_data_132 : _GEN_3520; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3522 = 8'h85 == _match_key_bytes_2_T_1 ? phv_data_133 : _GEN_3521; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3523 = 8'h86 == _match_key_bytes_2_T_1 ? phv_data_134 : _GEN_3522; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3524 = 8'h87 == _match_key_bytes_2_T_1 ? phv_data_135 : _GEN_3523; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3525 = 8'h88 == _match_key_bytes_2_T_1 ? phv_data_136 : _GEN_3524; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3526 = 8'h89 == _match_key_bytes_2_T_1 ? phv_data_137 : _GEN_3525; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3527 = 8'h8a == _match_key_bytes_2_T_1 ? phv_data_138 : _GEN_3526; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3528 = 8'h8b == _match_key_bytes_2_T_1 ? phv_data_139 : _GEN_3527; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3529 = 8'h8c == _match_key_bytes_2_T_1 ? phv_data_140 : _GEN_3528; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3530 = 8'h8d == _match_key_bytes_2_T_1 ? phv_data_141 : _GEN_3529; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3531 = 8'h8e == _match_key_bytes_2_T_1 ? phv_data_142 : _GEN_3530; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3532 = 8'h8f == _match_key_bytes_2_T_1 ? phv_data_143 : _GEN_3531; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3533 = 8'h90 == _match_key_bytes_2_T_1 ? phv_data_144 : _GEN_3532; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3534 = 8'h91 == _match_key_bytes_2_T_1 ? phv_data_145 : _GEN_3533; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3535 = 8'h92 == _match_key_bytes_2_T_1 ? phv_data_146 : _GEN_3534; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3536 = 8'h93 == _match_key_bytes_2_T_1 ? phv_data_147 : _GEN_3535; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3537 = 8'h94 == _match_key_bytes_2_T_1 ? phv_data_148 : _GEN_3536; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3538 = 8'h95 == _match_key_bytes_2_T_1 ? phv_data_149 : _GEN_3537; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3539 = 8'h96 == _match_key_bytes_2_T_1 ? phv_data_150 : _GEN_3538; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3540 = 8'h97 == _match_key_bytes_2_T_1 ? phv_data_151 : _GEN_3539; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3541 = 8'h98 == _match_key_bytes_2_T_1 ? phv_data_152 : _GEN_3540; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3542 = 8'h99 == _match_key_bytes_2_T_1 ? phv_data_153 : _GEN_3541; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3543 = 8'h9a == _match_key_bytes_2_T_1 ? phv_data_154 : _GEN_3542; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3544 = 8'h9b == _match_key_bytes_2_T_1 ? phv_data_155 : _GEN_3543; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3545 = 8'h9c == _match_key_bytes_2_T_1 ? phv_data_156 : _GEN_3544; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3546 = 8'h9d == _match_key_bytes_2_T_1 ? phv_data_157 : _GEN_3545; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3547 = 8'h9e == _match_key_bytes_2_T_1 ? phv_data_158 : _GEN_3546; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3548 = 8'h9f == _match_key_bytes_2_T_1 ? phv_data_159 : _GEN_3547; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_2 = 8'h15 < _GEN_6 ? _GEN_3548 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_1_T_1 = key_offset + 8'h16; // @[matcher.scala 72:98]
  wire [7:0] _GEN_3551 = 8'h1 == _match_key_bytes_1_T_1 ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3552 = 8'h2 == _match_key_bytes_1_T_1 ? phv_data_2 : _GEN_3551; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3553 = 8'h3 == _match_key_bytes_1_T_1 ? phv_data_3 : _GEN_3552; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3554 = 8'h4 == _match_key_bytes_1_T_1 ? phv_data_4 : _GEN_3553; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3555 = 8'h5 == _match_key_bytes_1_T_1 ? phv_data_5 : _GEN_3554; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3556 = 8'h6 == _match_key_bytes_1_T_1 ? phv_data_6 : _GEN_3555; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3557 = 8'h7 == _match_key_bytes_1_T_1 ? phv_data_7 : _GEN_3556; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3558 = 8'h8 == _match_key_bytes_1_T_1 ? phv_data_8 : _GEN_3557; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3559 = 8'h9 == _match_key_bytes_1_T_1 ? phv_data_9 : _GEN_3558; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3560 = 8'ha == _match_key_bytes_1_T_1 ? phv_data_10 : _GEN_3559; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3561 = 8'hb == _match_key_bytes_1_T_1 ? phv_data_11 : _GEN_3560; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3562 = 8'hc == _match_key_bytes_1_T_1 ? phv_data_12 : _GEN_3561; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3563 = 8'hd == _match_key_bytes_1_T_1 ? phv_data_13 : _GEN_3562; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3564 = 8'he == _match_key_bytes_1_T_1 ? phv_data_14 : _GEN_3563; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3565 = 8'hf == _match_key_bytes_1_T_1 ? phv_data_15 : _GEN_3564; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3566 = 8'h10 == _match_key_bytes_1_T_1 ? phv_data_16 : _GEN_3565; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3567 = 8'h11 == _match_key_bytes_1_T_1 ? phv_data_17 : _GEN_3566; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3568 = 8'h12 == _match_key_bytes_1_T_1 ? phv_data_18 : _GEN_3567; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3569 = 8'h13 == _match_key_bytes_1_T_1 ? phv_data_19 : _GEN_3568; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3570 = 8'h14 == _match_key_bytes_1_T_1 ? phv_data_20 : _GEN_3569; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3571 = 8'h15 == _match_key_bytes_1_T_1 ? phv_data_21 : _GEN_3570; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3572 = 8'h16 == _match_key_bytes_1_T_1 ? phv_data_22 : _GEN_3571; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3573 = 8'h17 == _match_key_bytes_1_T_1 ? phv_data_23 : _GEN_3572; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3574 = 8'h18 == _match_key_bytes_1_T_1 ? phv_data_24 : _GEN_3573; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3575 = 8'h19 == _match_key_bytes_1_T_1 ? phv_data_25 : _GEN_3574; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3576 = 8'h1a == _match_key_bytes_1_T_1 ? phv_data_26 : _GEN_3575; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3577 = 8'h1b == _match_key_bytes_1_T_1 ? phv_data_27 : _GEN_3576; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3578 = 8'h1c == _match_key_bytes_1_T_1 ? phv_data_28 : _GEN_3577; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3579 = 8'h1d == _match_key_bytes_1_T_1 ? phv_data_29 : _GEN_3578; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3580 = 8'h1e == _match_key_bytes_1_T_1 ? phv_data_30 : _GEN_3579; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3581 = 8'h1f == _match_key_bytes_1_T_1 ? phv_data_31 : _GEN_3580; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3582 = 8'h20 == _match_key_bytes_1_T_1 ? phv_data_32 : _GEN_3581; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3583 = 8'h21 == _match_key_bytes_1_T_1 ? phv_data_33 : _GEN_3582; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3584 = 8'h22 == _match_key_bytes_1_T_1 ? phv_data_34 : _GEN_3583; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3585 = 8'h23 == _match_key_bytes_1_T_1 ? phv_data_35 : _GEN_3584; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3586 = 8'h24 == _match_key_bytes_1_T_1 ? phv_data_36 : _GEN_3585; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3587 = 8'h25 == _match_key_bytes_1_T_1 ? phv_data_37 : _GEN_3586; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3588 = 8'h26 == _match_key_bytes_1_T_1 ? phv_data_38 : _GEN_3587; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3589 = 8'h27 == _match_key_bytes_1_T_1 ? phv_data_39 : _GEN_3588; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3590 = 8'h28 == _match_key_bytes_1_T_1 ? phv_data_40 : _GEN_3589; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3591 = 8'h29 == _match_key_bytes_1_T_1 ? phv_data_41 : _GEN_3590; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3592 = 8'h2a == _match_key_bytes_1_T_1 ? phv_data_42 : _GEN_3591; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3593 = 8'h2b == _match_key_bytes_1_T_1 ? phv_data_43 : _GEN_3592; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3594 = 8'h2c == _match_key_bytes_1_T_1 ? phv_data_44 : _GEN_3593; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3595 = 8'h2d == _match_key_bytes_1_T_1 ? phv_data_45 : _GEN_3594; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3596 = 8'h2e == _match_key_bytes_1_T_1 ? phv_data_46 : _GEN_3595; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3597 = 8'h2f == _match_key_bytes_1_T_1 ? phv_data_47 : _GEN_3596; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3598 = 8'h30 == _match_key_bytes_1_T_1 ? phv_data_48 : _GEN_3597; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3599 = 8'h31 == _match_key_bytes_1_T_1 ? phv_data_49 : _GEN_3598; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3600 = 8'h32 == _match_key_bytes_1_T_1 ? phv_data_50 : _GEN_3599; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3601 = 8'h33 == _match_key_bytes_1_T_1 ? phv_data_51 : _GEN_3600; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3602 = 8'h34 == _match_key_bytes_1_T_1 ? phv_data_52 : _GEN_3601; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3603 = 8'h35 == _match_key_bytes_1_T_1 ? phv_data_53 : _GEN_3602; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3604 = 8'h36 == _match_key_bytes_1_T_1 ? phv_data_54 : _GEN_3603; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3605 = 8'h37 == _match_key_bytes_1_T_1 ? phv_data_55 : _GEN_3604; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3606 = 8'h38 == _match_key_bytes_1_T_1 ? phv_data_56 : _GEN_3605; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3607 = 8'h39 == _match_key_bytes_1_T_1 ? phv_data_57 : _GEN_3606; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3608 = 8'h3a == _match_key_bytes_1_T_1 ? phv_data_58 : _GEN_3607; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3609 = 8'h3b == _match_key_bytes_1_T_1 ? phv_data_59 : _GEN_3608; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3610 = 8'h3c == _match_key_bytes_1_T_1 ? phv_data_60 : _GEN_3609; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3611 = 8'h3d == _match_key_bytes_1_T_1 ? phv_data_61 : _GEN_3610; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3612 = 8'h3e == _match_key_bytes_1_T_1 ? phv_data_62 : _GEN_3611; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3613 = 8'h3f == _match_key_bytes_1_T_1 ? phv_data_63 : _GEN_3612; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3614 = 8'h40 == _match_key_bytes_1_T_1 ? phv_data_64 : _GEN_3613; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3615 = 8'h41 == _match_key_bytes_1_T_1 ? phv_data_65 : _GEN_3614; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3616 = 8'h42 == _match_key_bytes_1_T_1 ? phv_data_66 : _GEN_3615; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3617 = 8'h43 == _match_key_bytes_1_T_1 ? phv_data_67 : _GEN_3616; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3618 = 8'h44 == _match_key_bytes_1_T_1 ? phv_data_68 : _GEN_3617; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3619 = 8'h45 == _match_key_bytes_1_T_1 ? phv_data_69 : _GEN_3618; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3620 = 8'h46 == _match_key_bytes_1_T_1 ? phv_data_70 : _GEN_3619; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3621 = 8'h47 == _match_key_bytes_1_T_1 ? phv_data_71 : _GEN_3620; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3622 = 8'h48 == _match_key_bytes_1_T_1 ? phv_data_72 : _GEN_3621; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3623 = 8'h49 == _match_key_bytes_1_T_1 ? phv_data_73 : _GEN_3622; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3624 = 8'h4a == _match_key_bytes_1_T_1 ? phv_data_74 : _GEN_3623; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3625 = 8'h4b == _match_key_bytes_1_T_1 ? phv_data_75 : _GEN_3624; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3626 = 8'h4c == _match_key_bytes_1_T_1 ? phv_data_76 : _GEN_3625; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3627 = 8'h4d == _match_key_bytes_1_T_1 ? phv_data_77 : _GEN_3626; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3628 = 8'h4e == _match_key_bytes_1_T_1 ? phv_data_78 : _GEN_3627; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3629 = 8'h4f == _match_key_bytes_1_T_1 ? phv_data_79 : _GEN_3628; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3630 = 8'h50 == _match_key_bytes_1_T_1 ? phv_data_80 : _GEN_3629; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3631 = 8'h51 == _match_key_bytes_1_T_1 ? phv_data_81 : _GEN_3630; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3632 = 8'h52 == _match_key_bytes_1_T_1 ? phv_data_82 : _GEN_3631; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3633 = 8'h53 == _match_key_bytes_1_T_1 ? phv_data_83 : _GEN_3632; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3634 = 8'h54 == _match_key_bytes_1_T_1 ? phv_data_84 : _GEN_3633; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3635 = 8'h55 == _match_key_bytes_1_T_1 ? phv_data_85 : _GEN_3634; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3636 = 8'h56 == _match_key_bytes_1_T_1 ? phv_data_86 : _GEN_3635; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3637 = 8'h57 == _match_key_bytes_1_T_1 ? phv_data_87 : _GEN_3636; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3638 = 8'h58 == _match_key_bytes_1_T_1 ? phv_data_88 : _GEN_3637; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3639 = 8'h59 == _match_key_bytes_1_T_1 ? phv_data_89 : _GEN_3638; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3640 = 8'h5a == _match_key_bytes_1_T_1 ? phv_data_90 : _GEN_3639; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3641 = 8'h5b == _match_key_bytes_1_T_1 ? phv_data_91 : _GEN_3640; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3642 = 8'h5c == _match_key_bytes_1_T_1 ? phv_data_92 : _GEN_3641; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3643 = 8'h5d == _match_key_bytes_1_T_1 ? phv_data_93 : _GEN_3642; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3644 = 8'h5e == _match_key_bytes_1_T_1 ? phv_data_94 : _GEN_3643; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3645 = 8'h5f == _match_key_bytes_1_T_1 ? phv_data_95 : _GEN_3644; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3646 = 8'h60 == _match_key_bytes_1_T_1 ? phv_data_96 : _GEN_3645; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3647 = 8'h61 == _match_key_bytes_1_T_1 ? phv_data_97 : _GEN_3646; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3648 = 8'h62 == _match_key_bytes_1_T_1 ? phv_data_98 : _GEN_3647; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3649 = 8'h63 == _match_key_bytes_1_T_1 ? phv_data_99 : _GEN_3648; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3650 = 8'h64 == _match_key_bytes_1_T_1 ? phv_data_100 : _GEN_3649; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3651 = 8'h65 == _match_key_bytes_1_T_1 ? phv_data_101 : _GEN_3650; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3652 = 8'h66 == _match_key_bytes_1_T_1 ? phv_data_102 : _GEN_3651; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3653 = 8'h67 == _match_key_bytes_1_T_1 ? phv_data_103 : _GEN_3652; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3654 = 8'h68 == _match_key_bytes_1_T_1 ? phv_data_104 : _GEN_3653; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3655 = 8'h69 == _match_key_bytes_1_T_1 ? phv_data_105 : _GEN_3654; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3656 = 8'h6a == _match_key_bytes_1_T_1 ? phv_data_106 : _GEN_3655; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3657 = 8'h6b == _match_key_bytes_1_T_1 ? phv_data_107 : _GEN_3656; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3658 = 8'h6c == _match_key_bytes_1_T_1 ? phv_data_108 : _GEN_3657; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3659 = 8'h6d == _match_key_bytes_1_T_1 ? phv_data_109 : _GEN_3658; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3660 = 8'h6e == _match_key_bytes_1_T_1 ? phv_data_110 : _GEN_3659; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3661 = 8'h6f == _match_key_bytes_1_T_1 ? phv_data_111 : _GEN_3660; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3662 = 8'h70 == _match_key_bytes_1_T_1 ? phv_data_112 : _GEN_3661; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3663 = 8'h71 == _match_key_bytes_1_T_1 ? phv_data_113 : _GEN_3662; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3664 = 8'h72 == _match_key_bytes_1_T_1 ? phv_data_114 : _GEN_3663; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3665 = 8'h73 == _match_key_bytes_1_T_1 ? phv_data_115 : _GEN_3664; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3666 = 8'h74 == _match_key_bytes_1_T_1 ? phv_data_116 : _GEN_3665; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3667 = 8'h75 == _match_key_bytes_1_T_1 ? phv_data_117 : _GEN_3666; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3668 = 8'h76 == _match_key_bytes_1_T_1 ? phv_data_118 : _GEN_3667; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3669 = 8'h77 == _match_key_bytes_1_T_1 ? phv_data_119 : _GEN_3668; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3670 = 8'h78 == _match_key_bytes_1_T_1 ? phv_data_120 : _GEN_3669; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3671 = 8'h79 == _match_key_bytes_1_T_1 ? phv_data_121 : _GEN_3670; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3672 = 8'h7a == _match_key_bytes_1_T_1 ? phv_data_122 : _GEN_3671; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3673 = 8'h7b == _match_key_bytes_1_T_1 ? phv_data_123 : _GEN_3672; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3674 = 8'h7c == _match_key_bytes_1_T_1 ? phv_data_124 : _GEN_3673; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3675 = 8'h7d == _match_key_bytes_1_T_1 ? phv_data_125 : _GEN_3674; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3676 = 8'h7e == _match_key_bytes_1_T_1 ? phv_data_126 : _GEN_3675; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3677 = 8'h7f == _match_key_bytes_1_T_1 ? phv_data_127 : _GEN_3676; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3678 = 8'h80 == _match_key_bytes_1_T_1 ? phv_data_128 : _GEN_3677; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3679 = 8'h81 == _match_key_bytes_1_T_1 ? phv_data_129 : _GEN_3678; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3680 = 8'h82 == _match_key_bytes_1_T_1 ? phv_data_130 : _GEN_3679; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3681 = 8'h83 == _match_key_bytes_1_T_1 ? phv_data_131 : _GEN_3680; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3682 = 8'h84 == _match_key_bytes_1_T_1 ? phv_data_132 : _GEN_3681; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3683 = 8'h85 == _match_key_bytes_1_T_1 ? phv_data_133 : _GEN_3682; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3684 = 8'h86 == _match_key_bytes_1_T_1 ? phv_data_134 : _GEN_3683; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3685 = 8'h87 == _match_key_bytes_1_T_1 ? phv_data_135 : _GEN_3684; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3686 = 8'h88 == _match_key_bytes_1_T_1 ? phv_data_136 : _GEN_3685; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3687 = 8'h89 == _match_key_bytes_1_T_1 ? phv_data_137 : _GEN_3686; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3688 = 8'h8a == _match_key_bytes_1_T_1 ? phv_data_138 : _GEN_3687; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3689 = 8'h8b == _match_key_bytes_1_T_1 ? phv_data_139 : _GEN_3688; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3690 = 8'h8c == _match_key_bytes_1_T_1 ? phv_data_140 : _GEN_3689; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3691 = 8'h8d == _match_key_bytes_1_T_1 ? phv_data_141 : _GEN_3690; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3692 = 8'h8e == _match_key_bytes_1_T_1 ? phv_data_142 : _GEN_3691; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3693 = 8'h8f == _match_key_bytes_1_T_1 ? phv_data_143 : _GEN_3692; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3694 = 8'h90 == _match_key_bytes_1_T_1 ? phv_data_144 : _GEN_3693; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3695 = 8'h91 == _match_key_bytes_1_T_1 ? phv_data_145 : _GEN_3694; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3696 = 8'h92 == _match_key_bytes_1_T_1 ? phv_data_146 : _GEN_3695; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3697 = 8'h93 == _match_key_bytes_1_T_1 ? phv_data_147 : _GEN_3696; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3698 = 8'h94 == _match_key_bytes_1_T_1 ? phv_data_148 : _GEN_3697; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3699 = 8'h95 == _match_key_bytes_1_T_1 ? phv_data_149 : _GEN_3698; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3700 = 8'h96 == _match_key_bytes_1_T_1 ? phv_data_150 : _GEN_3699; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3701 = 8'h97 == _match_key_bytes_1_T_1 ? phv_data_151 : _GEN_3700; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3702 = 8'h98 == _match_key_bytes_1_T_1 ? phv_data_152 : _GEN_3701; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3703 = 8'h99 == _match_key_bytes_1_T_1 ? phv_data_153 : _GEN_3702; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3704 = 8'h9a == _match_key_bytes_1_T_1 ? phv_data_154 : _GEN_3703; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3705 = 8'h9b == _match_key_bytes_1_T_1 ? phv_data_155 : _GEN_3704; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3706 = 8'h9c == _match_key_bytes_1_T_1 ? phv_data_156 : _GEN_3705; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3707 = 8'h9d == _match_key_bytes_1_T_1 ? phv_data_157 : _GEN_3706; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3708 = 8'h9e == _match_key_bytes_1_T_1 ? phv_data_158 : _GEN_3707; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3709 = 8'h9f == _match_key_bytes_1_T_1 ? phv_data_159 : _GEN_3708; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_1 = 8'h16 < _GEN_6 ? _GEN_3709 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_0_T_1 = key_offset + 8'h17; // @[matcher.scala 72:98]
  wire [7:0] _GEN_3712 = 8'h1 == _match_key_bytes_0_T_1 ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3713 = 8'h2 == _match_key_bytes_0_T_1 ? phv_data_2 : _GEN_3712; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3714 = 8'h3 == _match_key_bytes_0_T_1 ? phv_data_3 : _GEN_3713; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3715 = 8'h4 == _match_key_bytes_0_T_1 ? phv_data_4 : _GEN_3714; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3716 = 8'h5 == _match_key_bytes_0_T_1 ? phv_data_5 : _GEN_3715; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3717 = 8'h6 == _match_key_bytes_0_T_1 ? phv_data_6 : _GEN_3716; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3718 = 8'h7 == _match_key_bytes_0_T_1 ? phv_data_7 : _GEN_3717; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3719 = 8'h8 == _match_key_bytes_0_T_1 ? phv_data_8 : _GEN_3718; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3720 = 8'h9 == _match_key_bytes_0_T_1 ? phv_data_9 : _GEN_3719; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3721 = 8'ha == _match_key_bytes_0_T_1 ? phv_data_10 : _GEN_3720; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3722 = 8'hb == _match_key_bytes_0_T_1 ? phv_data_11 : _GEN_3721; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3723 = 8'hc == _match_key_bytes_0_T_1 ? phv_data_12 : _GEN_3722; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3724 = 8'hd == _match_key_bytes_0_T_1 ? phv_data_13 : _GEN_3723; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3725 = 8'he == _match_key_bytes_0_T_1 ? phv_data_14 : _GEN_3724; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3726 = 8'hf == _match_key_bytes_0_T_1 ? phv_data_15 : _GEN_3725; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3727 = 8'h10 == _match_key_bytes_0_T_1 ? phv_data_16 : _GEN_3726; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3728 = 8'h11 == _match_key_bytes_0_T_1 ? phv_data_17 : _GEN_3727; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3729 = 8'h12 == _match_key_bytes_0_T_1 ? phv_data_18 : _GEN_3728; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3730 = 8'h13 == _match_key_bytes_0_T_1 ? phv_data_19 : _GEN_3729; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3731 = 8'h14 == _match_key_bytes_0_T_1 ? phv_data_20 : _GEN_3730; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3732 = 8'h15 == _match_key_bytes_0_T_1 ? phv_data_21 : _GEN_3731; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3733 = 8'h16 == _match_key_bytes_0_T_1 ? phv_data_22 : _GEN_3732; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3734 = 8'h17 == _match_key_bytes_0_T_1 ? phv_data_23 : _GEN_3733; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3735 = 8'h18 == _match_key_bytes_0_T_1 ? phv_data_24 : _GEN_3734; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3736 = 8'h19 == _match_key_bytes_0_T_1 ? phv_data_25 : _GEN_3735; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3737 = 8'h1a == _match_key_bytes_0_T_1 ? phv_data_26 : _GEN_3736; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3738 = 8'h1b == _match_key_bytes_0_T_1 ? phv_data_27 : _GEN_3737; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3739 = 8'h1c == _match_key_bytes_0_T_1 ? phv_data_28 : _GEN_3738; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3740 = 8'h1d == _match_key_bytes_0_T_1 ? phv_data_29 : _GEN_3739; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3741 = 8'h1e == _match_key_bytes_0_T_1 ? phv_data_30 : _GEN_3740; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3742 = 8'h1f == _match_key_bytes_0_T_1 ? phv_data_31 : _GEN_3741; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3743 = 8'h20 == _match_key_bytes_0_T_1 ? phv_data_32 : _GEN_3742; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3744 = 8'h21 == _match_key_bytes_0_T_1 ? phv_data_33 : _GEN_3743; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3745 = 8'h22 == _match_key_bytes_0_T_1 ? phv_data_34 : _GEN_3744; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3746 = 8'h23 == _match_key_bytes_0_T_1 ? phv_data_35 : _GEN_3745; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3747 = 8'h24 == _match_key_bytes_0_T_1 ? phv_data_36 : _GEN_3746; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3748 = 8'h25 == _match_key_bytes_0_T_1 ? phv_data_37 : _GEN_3747; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3749 = 8'h26 == _match_key_bytes_0_T_1 ? phv_data_38 : _GEN_3748; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3750 = 8'h27 == _match_key_bytes_0_T_1 ? phv_data_39 : _GEN_3749; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3751 = 8'h28 == _match_key_bytes_0_T_1 ? phv_data_40 : _GEN_3750; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3752 = 8'h29 == _match_key_bytes_0_T_1 ? phv_data_41 : _GEN_3751; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3753 = 8'h2a == _match_key_bytes_0_T_1 ? phv_data_42 : _GEN_3752; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3754 = 8'h2b == _match_key_bytes_0_T_1 ? phv_data_43 : _GEN_3753; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3755 = 8'h2c == _match_key_bytes_0_T_1 ? phv_data_44 : _GEN_3754; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3756 = 8'h2d == _match_key_bytes_0_T_1 ? phv_data_45 : _GEN_3755; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3757 = 8'h2e == _match_key_bytes_0_T_1 ? phv_data_46 : _GEN_3756; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3758 = 8'h2f == _match_key_bytes_0_T_1 ? phv_data_47 : _GEN_3757; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3759 = 8'h30 == _match_key_bytes_0_T_1 ? phv_data_48 : _GEN_3758; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3760 = 8'h31 == _match_key_bytes_0_T_1 ? phv_data_49 : _GEN_3759; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3761 = 8'h32 == _match_key_bytes_0_T_1 ? phv_data_50 : _GEN_3760; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3762 = 8'h33 == _match_key_bytes_0_T_1 ? phv_data_51 : _GEN_3761; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3763 = 8'h34 == _match_key_bytes_0_T_1 ? phv_data_52 : _GEN_3762; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3764 = 8'h35 == _match_key_bytes_0_T_1 ? phv_data_53 : _GEN_3763; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3765 = 8'h36 == _match_key_bytes_0_T_1 ? phv_data_54 : _GEN_3764; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3766 = 8'h37 == _match_key_bytes_0_T_1 ? phv_data_55 : _GEN_3765; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3767 = 8'h38 == _match_key_bytes_0_T_1 ? phv_data_56 : _GEN_3766; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3768 = 8'h39 == _match_key_bytes_0_T_1 ? phv_data_57 : _GEN_3767; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3769 = 8'h3a == _match_key_bytes_0_T_1 ? phv_data_58 : _GEN_3768; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3770 = 8'h3b == _match_key_bytes_0_T_1 ? phv_data_59 : _GEN_3769; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3771 = 8'h3c == _match_key_bytes_0_T_1 ? phv_data_60 : _GEN_3770; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3772 = 8'h3d == _match_key_bytes_0_T_1 ? phv_data_61 : _GEN_3771; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3773 = 8'h3e == _match_key_bytes_0_T_1 ? phv_data_62 : _GEN_3772; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3774 = 8'h3f == _match_key_bytes_0_T_1 ? phv_data_63 : _GEN_3773; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3775 = 8'h40 == _match_key_bytes_0_T_1 ? phv_data_64 : _GEN_3774; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3776 = 8'h41 == _match_key_bytes_0_T_1 ? phv_data_65 : _GEN_3775; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3777 = 8'h42 == _match_key_bytes_0_T_1 ? phv_data_66 : _GEN_3776; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3778 = 8'h43 == _match_key_bytes_0_T_1 ? phv_data_67 : _GEN_3777; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3779 = 8'h44 == _match_key_bytes_0_T_1 ? phv_data_68 : _GEN_3778; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3780 = 8'h45 == _match_key_bytes_0_T_1 ? phv_data_69 : _GEN_3779; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3781 = 8'h46 == _match_key_bytes_0_T_1 ? phv_data_70 : _GEN_3780; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3782 = 8'h47 == _match_key_bytes_0_T_1 ? phv_data_71 : _GEN_3781; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3783 = 8'h48 == _match_key_bytes_0_T_1 ? phv_data_72 : _GEN_3782; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3784 = 8'h49 == _match_key_bytes_0_T_1 ? phv_data_73 : _GEN_3783; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3785 = 8'h4a == _match_key_bytes_0_T_1 ? phv_data_74 : _GEN_3784; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3786 = 8'h4b == _match_key_bytes_0_T_1 ? phv_data_75 : _GEN_3785; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3787 = 8'h4c == _match_key_bytes_0_T_1 ? phv_data_76 : _GEN_3786; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3788 = 8'h4d == _match_key_bytes_0_T_1 ? phv_data_77 : _GEN_3787; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3789 = 8'h4e == _match_key_bytes_0_T_1 ? phv_data_78 : _GEN_3788; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3790 = 8'h4f == _match_key_bytes_0_T_1 ? phv_data_79 : _GEN_3789; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3791 = 8'h50 == _match_key_bytes_0_T_1 ? phv_data_80 : _GEN_3790; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3792 = 8'h51 == _match_key_bytes_0_T_1 ? phv_data_81 : _GEN_3791; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3793 = 8'h52 == _match_key_bytes_0_T_1 ? phv_data_82 : _GEN_3792; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3794 = 8'h53 == _match_key_bytes_0_T_1 ? phv_data_83 : _GEN_3793; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3795 = 8'h54 == _match_key_bytes_0_T_1 ? phv_data_84 : _GEN_3794; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3796 = 8'h55 == _match_key_bytes_0_T_1 ? phv_data_85 : _GEN_3795; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3797 = 8'h56 == _match_key_bytes_0_T_1 ? phv_data_86 : _GEN_3796; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3798 = 8'h57 == _match_key_bytes_0_T_1 ? phv_data_87 : _GEN_3797; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3799 = 8'h58 == _match_key_bytes_0_T_1 ? phv_data_88 : _GEN_3798; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3800 = 8'h59 == _match_key_bytes_0_T_1 ? phv_data_89 : _GEN_3799; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3801 = 8'h5a == _match_key_bytes_0_T_1 ? phv_data_90 : _GEN_3800; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3802 = 8'h5b == _match_key_bytes_0_T_1 ? phv_data_91 : _GEN_3801; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3803 = 8'h5c == _match_key_bytes_0_T_1 ? phv_data_92 : _GEN_3802; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3804 = 8'h5d == _match_key_bytes_0_T_1 ? phv_data_93 : _GEN_3803; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3805 = 8'h5e == _match_key_bytes_0_T_1 ? phv_data_94 : _GEN_3804; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3806 = 8'h5f == _match_key_bytes_0_T_1 ? phv_data_95 : _GEN_3805; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3807 = 8'h60 == _match_key_bytes_0_T_1 ? phv_data_96 : _GEN_3806; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3808 = 8'h61 == _match_key_bytes_0_T_1 ? phv_data_97 : _GEN_3807; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3809 = 8'h62 == _match_key_bytes_0_T_1 ? phv_data_98 : _GEN_3808; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3810 = 8'h63 == _match_key_bytes_0_T_1 ? phv_data_99 : _GEN_3809; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3811 = 8'h64 == _match_key_bytes_0_T_1 ? phv_data_100 : _GEN_3810; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3812 = 8'h65 == _match_key_bytes_0_T_1 ? phv_data_101 : _GEN_3811; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3813 = 8'h66 == _match_key_bytes_0_T_1 ? phv_data_102 : _GEN_3812; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3814 = 8'h67 == _match_key_bytes_0_T_1 ? phv_data_103 : _GEN_3813; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3815 = 8'h68 == _match_key_bytes_0_T_1 ? phv_data_104 : _GEN_3814; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3816 = 8'h69 == _match_key_bytes_0_T_1 ? phv_data_105 : _GEN_3815; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3817 = 8'h6a == _match_key_bytes_0_T_1 ? phv_data_106 : _GEN_3816; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3818 = 8'h6b == _match_key_bytes_0_T_1 ? phv_data_107 : _GEN_3817; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3819 = 8'h6c == _match_key_bytes_0_T_1 ? phv_data_108 : _GEN_3818; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3820 = 8'h6d == _match_key_bytes_0_T_1 ? phv_data_109 : _GEN_3819; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3821 = 8'h6e == _match_key_bytes_0_T_1 ? phv_data_110 : _GEN_3820; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3822 = 8'h6f == _match_key_bytes_0_T_1 ? phv_data_111 : _GEN_3821; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3823 = 8'h70 == _match_key_bytes_0_T_1 ? phv_data_112 : _GEN_3822; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3824 = 8'h71 == _match_key_bytes_0_T_1 ? phv_data_113 : _GEN_3823; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3825 = 8'h72 == _match_key_bytes_0_T_1 ? phv_data_114 : _GEN_3824; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3826 = 8'h73 == _match_key_bytes_0_T_1 ? phv_data_115 : _GEN_3825; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3827 = 8'h74 == _match_key_bytes_0_T_1 ? phv_data_116 : _GEN_3826; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3828 = 8'h75 == _match_key_bytes_0_T_1 ? phv_data_117 : _GEN_3827; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3829 = 8'h76 == _match_key_bytes_0_T_1 ? phv_data_118 : _GEN_3828; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3830 = 8'h77 == _match_key_bytes_0_T_1 ? phv_data_119 : _GEN_3829; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3831 = 8'h78 == _match_key_bytes_0_T_1 ? phv_data_120 : _GEN_3830; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3832 = 8'h79 == _match_key_bytes_0_T_1 ? phv_data_121 : _GEN_3831; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3833 = 8'h7a == _match_key_bytes_0_T_1 ? phv_data_122 : _GEN_3832; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3834 = 8'h7b == _match_key_bytes_0_T_1 ? phv_data_123 : _GEN_3833; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3835 = 8'h7c == _match_key_bytes_0_T_1 ? phv_data_124 : _GEN_3834; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3836 = 8'h7d == _match_key_bytes_0_T_1 ? phv_data_125 : _GEN_3835; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3837 = 8'h7e == _match_key_bytes_0_T_1 ? phv_data_126 : _GEN_3836; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3838 = 8'h7f == _match_key_bytes_0_T_1 ? phv_data_127 : _GEN_3837; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3839 = 8'h80 == _match_key_bytes_0_T_1 ? phv_data_128 : _GEN_3838; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3840 = 8'h81 == _match_key_bytes_0_T_1 ? phv_data_129 : _GEN_3839; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3841 = 8'h82 == _match_key_bytes_0_T_1 ? phv_data_130 : _GEN_3840; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3842 = 8'h83 == _match_key_bytes_0_T_1 ? phv_data_131 : _GEN_3841; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3843 = 8'h84 == _match_key_bytes_0_T_1 ? phv_data_132 : _GEN_3842; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3844 = 8'h85 == _match_key_bytes_0_T_1 ? phv_data_133 : _GEN_3843; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3845 = 8'h86 == _match_key_bytes_0_T_1 ? phv_data_134 : _GEN_3844; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3846 = 8'h87 == _match_key_bytes_0_T_1 ? phv_data_135 : _GEN_3845; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3847 = 8'h88 == _match_key_bytes_0_T_1 ? phv_data_136 : _GEN_3846; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3848 = 8'h89 == _match_key_bytes_0_T_1 ? phv_data_137 : _GEN_3847; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3849 = 8'h8a == _match_key_bytes_0_T_1 ? phv_data_138 : _GEN_3848; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3850 = 8'h8b == _match_key_bytes_0_T_1 ? phv_data_139 : _GEN_3849; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3851 = 8'h8c == _match_key_bytes_0_T_1 ? phv_data_140 : _GEN_3850; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3852 = 8'h8d == _match_key_bytes_0_T_1 ? phv_data_141 : _GEN_3851; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3853 = 8'h8e == _match_key_bytes_0_T_1 ? phv_data_142 : _GEN_3852; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3854 = 8'h8f == _match_key_bytes_0_T_1 ? phv_data_143 : _GEN_3853; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3855 = 8'h90 == _match_key_bytes_0_T_1 ? phv_data_144 : _GEN_3854; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3856 = 8'h91 == _match_key_bytes_0_T_1 ? phv_data_145 : _GEN_3855; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3857 = 8'h92 == _match_key_bytes_0_T_1 ? phv_data_146 : _GEN_3856; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3858 = 8'h93 == _match_key_bytes_0_T_1 ? phv_data_147 : _GEN_3857; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3859 = 8'h94 == _match_key_bytes_0_T_1 ? phv_data_148 : _GEN_3858; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3860 = 8'h95 == _match_key_bytes_0_T_1 ? phv_data_149 : _GEN_3859; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3861 = 8'h96 == _match_key_bytes_0_T_1 ? phv_data_150 : _GEN_3860; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3862 = 8'h97 == _match_key_bytes_0_T_1 ? phv_data_151 : _GEN_3861; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3863 = 8'h98 == _match_key_bytes_0_T_1 ? phv_data_152 : _GEN_3862; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3864 = 8'h99 == _match_key_bytes_0_T_1 ? phv_data_153 : _GEN_3863; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3865 = 8'h9a == _match_key_bytes_0_T_1 ? phv_data_154 : _GEN_3864; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3866 = 8'h9b == _match_key_bytes_0_T_1 ? phv_data_155 : _GEN_3865; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3867 = 8'h9c == _match_key_bytes_0_T_1 ? phv_data_156 : _GEN_3866; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3868 = 8'h9d == _match_key_bytes_0_T_1 ? phv_data_157 : _GEN_3867; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3869 = 8'h9e == _match_key_bytes_0_T_1 ? phv_data_158 : _GEN_3868; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_3870 = 8'h9f == _match_key_bytes_0_T_1 ? phv_data_159 : _GEN_3869; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_0 = 8'h17 < _GEN_6 ? _GEN_3870 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [79:0] match_key_hi_8 = {match_key_bytes_0,match_key_bytes_1,match_key_bytes_2,match_key_bytes_3,
    match_key_bytes_4,match_key_bytes_5,match_key_bytes_6,match_key_bytes_7,match_key_bytes_8,match_key_bytes_9}; // @[Cat.scala 30:58]
  wire [151:0] match_key_hi_17 = {match_key_hi_8,match_key_bytes_10,match_key_bytes_11,match_key_bytes_12,
    match_key_bytes_13,match_key_bytes_14,match_key_bytes_15,match_key_bytes_16,match_key_bytes_17,match_key_bytes_18}; // @[Cat.scala 30:58]
  wire [191:0] match_key = {match_key_hi_17,match_key_bytes_19,match_key_bytes_20,match_key_bytes_21,match_key_bytes_22,
    match_key_bytes_23}; // @[Cat.scala 30:58]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_96 = phv_data_96; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_97 = phv_data_97; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_98 = phv_data_98; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_99 = phv_data_99; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_100 = phv_data_100; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_101 = phv_data_101; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_102 = phv_data_102; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_103 = phv_data_103; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_104 = phv_data_104; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_105 = phv_data_105; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_106 = phv_data_106; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_107 = phv_data_107; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_108 = phv_data_108; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_109 = phv_data_109; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_110 = phv_data_110; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_111 = phv_data_111; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_112 = phv_data_112; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_113 = phv_data_113; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_114 = phv_data_114; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_115 = phv_data_115; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_116 = phv_data_116; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_117 = phv_data_117; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_118 = phv_data_118; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_119 = phv_data_119; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_120 = phv_data_120; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_121 = phv_data_121; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_122 = phv_data_122; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_123 = phv_data_123; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_124 = phv_data_124; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_125 = phv_data_125; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_126 = phv_data_126; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_127 = phv_data_127; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_128 = phv_data_128; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_129 = phv_data_129; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_130 = phv_data_130; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_131 = phv_data_131; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_132 = phv_data_132; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_133 = phv_data_133; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_134 = phv_data_134; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_135 = phv_data_135; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_136 = phv_data_136; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_137 = phv_data_137; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_138 = phv_data_138; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_139 = phv_data_139; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_140 = phv_data_140; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_141 = phv_data_141; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_142 = phv_data_142; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_143 = phv_data_143; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_144 = phv_data_144; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_145 = phv_data_145; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_146 = phv_data_146; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_147 = phv_data_147; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_148 = phv_data_148; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_149 = phv_data_149; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_150 = phv_data_150; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_151 = phv_data_151; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_152 = phv_data_152; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_153 = phv_data_153; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_154 = phv_data_154; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_155 = phv_data_155; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_156 = phv_data_156; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_157 = phv_data_157; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_158 = phv_data_158; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_159 = phv_data_159; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[matcher.scala 60:25]
  assign io_match_key = phv_is_valid_processor ? match_key : 192'h0; // @[matcher.scala 65:39 matcher.scala 79:26 matcher.scala 81:26]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[matcher.scala 59:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[matcher.scala 59:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[matcher.scala 59:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[matcher.scala 59:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[matcher.scala 59:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[matcher.scala 59:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[matcher.scala 59:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[matcher.scala 59:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[matcher.scala 59:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[matcher.scala 59:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[matcher.scala 59:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[matcher.scala 59:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[matcher.scala 59:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[matcher.scala 59:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[matcher.scala 59:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[matcher.scala 59:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[matcher.scala 59:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[matcher.scala 59:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[matcher.scala 59:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[matcher.scala 59:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[matcher.scala 59:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[matcher.scala 59:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[matcher.scala 59:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[matcher.scala 59:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[matcher.scala 59:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[matcher.scala 59:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[matcher.scala 59:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[matcher.scala 59:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[matcher.scala 59:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[matcher.scala 59:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[matcher.scala 59:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[matcher.scala 59:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[matcher.scala 59:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[matcher.scala 59:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[matcher.scala 59:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[matcher.scala 59:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[matcher.scala 59:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[matcher.scala 59:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[matcher.scala 59:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[matcher.scala 59:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[matcher.scala 59:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[matcher.scala 59:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[matcher.scala 59:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[matcher.scala 59:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[matcher.scala 59:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[matcher.scala 59:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[matcher.scala 59:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[matcher.scala 59:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[matcher.scala 59:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[matcher.scala 59:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[matcher.scala 59:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[matcher.scala 59:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[matcher.scala 59:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[matcher.scala 59:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[matcher.scala 59:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[matcher.scala 59:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[matcher.scala 59:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[matcher.scala 59:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[matcher.scala 59:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[matcher.scala 59:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[matcher.scala 59:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[matcher.scala 59:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[matcher.scala 59:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[matcher.scala 59:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[matcher.scala 59:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[matcher.scala 59:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[matcher.scala 59:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[matcher.scala 59:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[matcher.scala 59:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[matcher.scala 59:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[matcher.scala 59:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[matcher.scala 59:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[matcher.scala 59:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[matcher.scala 59:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[matcher.scala 59:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[matcher.scala 59:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[matcher.scala 59:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[matcher.scala 59:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[matcher.scala 59:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[matcher.scala 59:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[matcher.scala 59:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[matcher.scala 59:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[matcher.scala 59:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[matcher.scala 59:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[matcher.scala 59:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[matcher.scala 59:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[matcher.scala 59:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[matcher.scala 59:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[matcher.scala 59:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[matcher.scala 59:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[matcher.scala 59:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[matcher.scala 59:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[matcher.scala 59:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[matcher.scala 59:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[matcher.scala 59:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[matcher.scala 59:13]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[matcher.scala 59:13]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[matcher.scala 59:13]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[matcher.scala 59:13]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[matcher.scala 59:13]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[matcher.scala 59:13]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[matcher.scala 59:13]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[matcher.scala 59:13]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[matcher.scala 59:13]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[matcher.scala 59:13]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[matcher.scala 59:13]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[matcher.scala 59:13]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[matcher.scala 59:13]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[matcher.scala 59:13]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[matcher.scala 59:13]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[matcher.scala 59:13]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[matcher.scala 59:13]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[matcher.scala 59:13]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[matcher.scala 59:13]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[matcher.scala 59:13]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[matcher.scala 59:13]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[matcher.scala 59:13]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[matcher.scala 59:13]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[matcher.scala 59:13]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[matcher.scala 59:13]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[matcher.scala 59:13]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[matcher.scala 59:13]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[matcher.scala 59:13]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[matcher.scala 59:13]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[matcher.scala 59:13]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[matcher.scala 59:13]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[matcher.scala 59:13]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[matcher.scala 59:13]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[matcher.scala 59:13]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[matcher.scala 59:13]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[matcher.scala 59:13]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[matcher.scala 59:13]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[matcher.scala 59:13]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[matcher.scala 59:13]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[matcher.scala 59:13]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[matcher.scala 59:13]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[matcher.scala 59:13]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[matcher.scala 59:13]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[matcher.scala 59:13]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[matcher.scala 59:13]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[matcher.scala 59:13]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[matcher.scala 59:13]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[matcher.scala 59:13]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[matcher.scala 59:13]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[matcher.scala 59:13]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[matcher.scala 59:13]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[matcher.scala 59:13]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[matcher.scala 59:13]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[matcher.scala 59:13]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[matcher.scala 59:13]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[matcher.scala 59:13]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[matcher.scala 59:13]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[matcher.scala 59:13]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[matcher.scala 59:13]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[matcher.scala 59:13]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[matcher.scala 59:13]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[matcher.scala 59:13]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[matcher.scala 59:13]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[matcher.scala 59:13]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[matcher.scala 59:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[matcher.scala 59:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[matcher.scala 59:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[matcher.scala 59:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[matcher.scala 59:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[matcher.scala 59:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[matcher.scala 59:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[matcher.scala 59:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[matcher.scala 59:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[matcher.scala 59:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[matcher.scala 59:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[matcher.scala 59:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[matcher.scala 59:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[matcher.scala 59:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[matcher.scala 59:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[matcher.scala 59:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[matcher.scala 59:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[matcher.scala 59:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[matcher.scala 59:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[matcher.scala 59:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[matcher.scala 59:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[matcher.scala 59:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[matcher.scala 59:13]
    key_offset <= io_key_offset; // @[matcher.scala 63:20]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_header_0 = _RAND_160[15:0];
  _RAND_161 = {1{`RANDOM}};
  phv_header_1 = _RAND_161[15:0];
  _RAND_162 = {1{`RANDOM}};
  phv_header_2 = _RAND_162[15:0];
  _RAND_163 = {1{`RANDOM}};
  phv_header_3 = _RAND_163[15:0];
  _RAND_164 = {1{`RANDOM}};
  phv_header_4 = _RAND_164[15:0];
  _RAND_165 = {1{`RANDOM}};
  phv_header_5 = _RAND_165[15:0];
  _RAND_166 = {1{`RANDOM}};
  phv_header_6 = _RAND_166[15:0];
  _RAND_167 = {1{`RANDOM}};
  phv_header_7 = _RAND_167[15:0];
  _RAND_168 = {1{`RANDOM}};
  phv_header_8 = _RAND_168[15:0];
  _RAND_169 = {1{`RANDOM}};
  phv_header_9 = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  phv_header_10 = _RAND_170[15:0];
  _RAND_171 = {1{`RANDOM}};
  phv_header_11 = _RAND_171[15:0];
  _RAND_172 = {1{`RANDOM}};
  phv_header_12 = _RAND_172[15:0];
  _RAND_173 = {1{`RANDOM}};
  phv_header_13 = _RAND_173[15:0];
  _RAND_174 = {1{`RANDOM}};
  phv_header_14 = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  phv_header_15 = _RAND_175[15:0];
  _RAND_176 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_178[15:0];
  _RAND_179 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_179[3:0];
  _RAND_180 = {1{`RANDOM}};
  phv_next_config_id = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  key_offset = _RAND_182[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
