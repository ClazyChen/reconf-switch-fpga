module MatchGetKey(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [1:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [1:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input  [3:0]  io_key_config_0_key_length,
  input  [3:0]  io_key_config_1_key_length,
  input  [7:0]  io_key_offset,
  output [63:0] io_match_key
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[matcher.scala 58:22]
  reg [7:0] phv_data_1; // @[matcher.scala 58:22]
  reg [7:0] phv_data_2; // @[matcher.scala 58:22]
  reg [7:0] phv_data_3; // @[matcher.scala 58:22]
  reg [7:0] phv_data_4; // @[matcher.scala 58:22]
  reg [7:0] phv_data_5; // @[matcher.scala 58:22]
  reg [7:0] phv_data_6; // @[matcher.scala 58:22]
  reg [7:0] phv_data_7; // @[matcher.scala 58:22]
  reg [7:0] phv_data_8; // @[matcher.scala 58:22]
  reg [7:0] phv_data_9; // @[matcher.scala 58:22]
  reg [7:0] phv_data_10; // @[matcher.scala 58:22]
  reg [7:0] phv_data_11; // @[matcher.scala 58:22]
  reg [7:0] phv_data_12; // @[matcher.scala 58:22]
  reg [7:0] phv_data_13; // @[matcher.scala 58:22]
  reg [7:0] phv_data_14; // @[matcher.scala 58:22]
  reg [7:0] phv_data_15; // @[matcher.scala 58:22]
  reg [7:0] phv_data_16; // @[matcher.scala 58:22]
  reg [7:0] phv_data_17; // @[matcher.scala 58:22]
  reg [7:0] phv_data_18; // @[matcher.scala 58:22]
  reg [7:0] phv_data_19; // @[matcher.scala 58:22]
  reg [7:0] phv_data_20; // @[matcher.scala 58:22]
  reg [7:0] phv_data_21; // @[matcher.scala 58:22]
  reg [7:0] phv_data_22; // @[matcher.scala 58:22]
  reg [7:0] phv_data_23; // @[matcher.scala 58:22]
  reg [7:0] phv_data_24; // @[matcher.scala 58:22]
  reg [7:0] phv_data_25; // @[matcher.scala 58:22]
  reg [7:0] phv_data_26; // @[matcher.scala 58:22]
  reg [7:0] phv_data_27; // @[matcher.scala 58:22]
  reg [7:0] phv_data_28; // @[matcher.scala 58:22]
  reg [7:0] phv_data_29; // @[matcher.scala 58:22]
  reg [7:0] phv_data_30; // @[matcher.scala 58:22]
  reg [7:0] phv_data_31; // @[matcher.scala 58:22]
  reg [7:0] phv_data_32; // @[matcher.scala 58:22]
  reg [7:0] phv_data_33; // @[matcher.scala 58:22]
  reg [7:0] phv_data_34; // @[matcher.scala 58:22]
  reg [7:0] phv_data_35; // @[matcher.scala 58:22]
  reg [7:0] phv_data_36; // @[matcher.scala 58:22]
  reg [7:0] phv_data_37; // @[matcher.scala 58:22]
  reg [7:0] phv_data_38; // @[matcher.scala 58:22]
  reg [7:0] phv_data_39; // @[matcher.scala 58:22]
  reg [7:0] phv_data_40; // @[matcher.scala 58:22]
  reg [7:0] phv_data_41; // @[matcher.scala 58:22]
  reg [7:0] phv_data_42; // @[matcher.scala 58:22]
  reg [7:0] phv_data_43; // @[matcher.scala 58:22]
  reg [7:0] phv_data_44; // @[matcher.scala 58:22]
  reg [7:0] phv_data_45; // @[matcher.scala 58:22]
  reg [7:0] phv_data_46; // @[matcher.scala 58:22]
  reg [7:0] phv_data_47; // @[matcher.scala 58:22]
  reg [7:0] phv_data_48; // @[matcher.scala 58:22]
  reg [7:0] phv_data_49; // @[matcher.scala 58:22]
  reg [7:0] phv_data_50; // @[matcher.scala 58:22]
  reg [7:0] phv_data_51; // @[matcher.scala 58:22]
  reg [7:0] phv_data_52; // @[matcher.scala 58:22]
  reg [7:0] phv_data_53; // @[matcher.scala 58:22]
  reg [7:0] phv_data_54; // @[matcher.scala 58:22]
  reg [7:0] phv_data_55; // @[matcher.scala 58:22]
  reg [7:0] phv_data_56; // @[matcher.scala 58:22]
  reg [7:0] phv_data_57; // @[matcher.scala 58:22]
  reg [7:0] phv_data_58; // @[matcher.scala 58:22]
  reg [7:0] phv_data_59; // @[matcher.scala 58:22]
  reg [7:0] phv_data_60; // @[matcher.scala 58:22]
  reg [7:0] phv_data_61; // @[matcher.scala 58:22]
  reg [7:0] phv_data_62; // @[matcher.scala 58:22]
  reg [7:0] phv_data_63; // @[matcher.scala 58:22]
  reg [7:0] phv_data_64; // @[matcher.scala 58:22]
  reg [7:0] phv_data_65; // @[matcher.scala 58:22]
  reg [7:0] phv_data_66; // @[matcher.scala 58:22]
  reg [7:0] phv_data_67; // @[matcher.scala 58:22]
  reg [7:0] phv_data_68; // @[matcher.scala 58:22]
  reg [7:0] phv_data_69; // @[matcher.scala 58:22]
  reg [7:0] phv_data_70; // @[matcher.scala 58:22]
  reg [7:0] phv_data_71; // @[matcher.scala 58:22]
  reg [7:0] phv_data_72; // @[matcher.scala 58:22]
  reg [7:0] phv_data_73; // @[matcher.scala 58:22]
  reg [7:0] phv_data_74; // @[matcher.scala 58:22]
  reg [7:0] phv_data_75; // @[matcher.scala 58:22]
  reg [7:0] phv_data_76; // @[matcher.scala 58:22]
  reg [7:0] phv_data_77; // @[matcher.scala 58:22]
  reg [7:0] phv_data_78; // @[matcher.scala 58:22]
  reg [7:0] phv_data_79; // @[matcher.scala 58:22]
  reg [7:0] phv_data_80; // @[matcher.scala 58:22]
  reg [7:0] phv_data_81; // @[matcher.scala 58:22]
  reg [7:0] phv_data_82; // @[matcher.scala 58:22]
  reg [7:0] phv_data_83; // @[matcher.scala 58:22]
  reg [7:0] phv_data_84; // @[matcher.scala 58:22]
  reg [7:0] phv_data_85; // @[matcher.scala 58:22]
  reg [7:0] phv_data_86; // @[matcher.scala 58:22]
  reg [7:0] phv_data_87; // @[matcher.scala 58:22]
  reg [7:0] phv_data_88; // @[matcher.scala 58:22]
  reg [7:0] phv_data_89; // @[matcher.scala 58:22]
  reg [7:0] phv_data_90; // @[matcher.scala 58:22]
  reg [7:0] phv_data_91; // @[matcher.scala 58:22]
  reg [7:0] phv_data_92; // @[matcher.scala 58:22]
  reg [7:0] phv_data_93; // @[matcher.scala 58:22]
  reg [7:0] phv_data_94; // @[matcher.scala 58:22]
  reg [7:0] phv_data_95; // @[matcher.scala 58:22]
  reg [15:0] phv_header_0; // @[matcher.scala 58:22]
  reg [15:0] phv_header_1; // @[matcher.scala 58:22]
  reg [15:0] phv_header_2; // @[matcher.scala 58:22]
  reg [15:0] phv_header_3; // @[matcher.scala 58:22]
  reg [15:0] phv_header_4; // @[matcher.scala 58:22]
  reg [15:0] phv_header_5; // @[matcher.scala 58:22]
  reg [15:0] phv_header_6; // @[matcher.scala 58:22]
  reg [15:0] phv_header_7; // @[matcher.scala 58:22]
  reg [15:0] phv_header_8; // @[matcher.scala 58:22]
  reg [15:0] phv_header_9; // @[matcher.scala 58:22]
  reg [15:0] phv_header_10; // @[matcher.scala 58:22]
  reg [15:0] phv_header_11; // @[matcher.scala 58:22]
  reg [15:0] phv_header_12; // @[matcher.scala 58:22]
  reg [15:0] phv_header_13; // @[matcher.scala 58:22]
  reg [15:0] phv_header_14; // @[matcher.scala 58:22]
  reg [15:0] phv_header_15; // @[matcher.scala 58:22]
  reg [7:0] phv_parse_current_state; // @[matcher.scala 58:22]
  reg [7:0] phv_parse_current_offset; // @[matcher.scala 58:22]
  reg [15:0] phv_parse_transition_field; // @[matcher.scala 58:22]
  reg [1:0] phv_next_processor_id; // @[matcher.scala 58:22]
  reg  phv_next_config_id; // @[matcher.scala 58:22]
  reg  phv_is_valid_processor; // @[matcher.scala 58:22]
  reg [7:0] key_offset; // @[matcher.scala 62:29]
  wire [3:0] _GEN_6 = phv_next_config_id ? io_key_config_1_key_length : io_key_config_0_key_length; // @[matcher.scala 71:36 matcher.scala 71:36]
  wire [8:0] _match_key_bytes_7_T = {{1'd0}, key_offset}; // @[matcher.scala 72:98]
  wire [7:0] _GEN_9 = 7'h1 == _match_key_bytes_7_T[6:0] ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_10 = 7'h2 == _match_key_bytes_7_T[6:0] ? phv_data_2 : _GEN_9; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_11 = 7'h3 == _match_key_bytes_7_T[6:0] ? phv_data_3 : _GEN_10; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_12 = 7'h4 == _match_key_bytes_7_T[6:0] ? phv_data_4 : _GEN_11; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_13 = 7'h5 == _match_key_bytes_7_T[6:0] ? phv_data_5 : _GEN_12; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_14 = 7'h6 == _match_key_bytes_7_T[6:0] ? phv_data_6 : _GEN_13; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_15 = 7'h7 == _match_key_bytes_7_T[6:0] ? phv_data_7 : _GEN_14; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_16 = 7'h8 == _match_key_bytes_7_T[6:0] ? phv_data_8 : _GEN_15; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_17 = 7'h9 == _match_key_bytes_7_T[6:0] ? phv_data_9 : _GEN_16; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_18 = 7'ha == _match_key_bytes_7_T[6:0] ? phv_data_10 : _GEN_17; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_19 = 7'hb == _match_key_bytes_7_T[6:0] ? phv_data_11 : _GEN_18; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_20 = 7'hc == _match_key_bytes_7_T[6:0] ? phv_data_12 : _GEN_19; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_21 = 7'hd == _match_key_bytes_7_T[6:0] ? phv_data_13 : _GEN_20; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_22 = 7'he == _match_key_bytes_7_T[6:0] ? phv_data_14 : _GEN_21; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_23 = 7'hf == _match_key_bytes_7_T[6:0] ? phv_data_15 : _GEN_22; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_24 = 7'h10 == _match_key_bytes_7_T[6:0] ? phv_data_16 : _GEN_23; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_25 = 7'h11 == _match_key_bytes_7_T[6:0] ? phv_data_17 : _GEN_24; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_26 = 7'h12 == _match_key_bytes_7_T[6:0] ? phv_data_18 : _GEN_25; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_27 = 7'h13 == _match_key_bytes_7_T[6:0] ? phv_data_19 : _GEN_26; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_28 = 7'h14 == _match_key_bytes_7_T[6:0] ? phv_data_20 : _GEN_27; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_29 = 7'h15 == _match_key_bytes_7_T[6:0] ? phv_data_21 : _GEN_28; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_30 = 7'h16 == _match_key_bytes_7_T[6:0] ? phv_data_22 : _GEN_29; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_31 = 7'h17 == _match_key_bytes_7_T[6:0] ? phv_data_23 : _GEN_30; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_32 = 7'h18 == _match_key_bytes_7_T[6:0] ? phv_data_24 : _GEN_31; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_33 = 7'h19 == _match_key_bytes_7_T[6:0] ? phv_data_25 : _GEN_32; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_34 = 7'h1a == _match_key_bytes_7_T[6:0] ? phv_data_26 : _GEN_33; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_35 = 7'h1b == _match_key_bytes_7_T[6:0] ? phv_data_27 : _GEN_34; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_36 = 7'h1c == _match_key_bytes_7_T[6:0] ? phv_data_28 : _GEN_35; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_37 = 7'h1d == _match_key_bytes_7_T[6:0] ? phv_data_29 : _GEN_36; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_38 = 7'h1e == _match_key_bytes_7_T[6:0] ? phv_data_30 : _GEN_37; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_39 = 7'h1f == _match_key_bytes_7_T[6:0] ? phv_data_31 : _GEN_38; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_40 = 7'h20 == _match_key_bytes_7_T[6:0] ? phv_data_32 : _GEN_39; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_41 = 7'h21 == _match_key_bytes_7_T[6:0] ? phv_data_33 : _GEN_40; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_42 = 7'h22 == _match_key_bytes_7_T[6:0] ? phv_data_34 : _GEN_41; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_43 = 7'h23 == _match_key_bytes_7_T[6:0] ? phv_data_35 : _GEN_42; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_44 = 7'h24 == _match_key_bytes_7_T[6:0] ? phv_data_36 : _GEN_43; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_45 = 7'h25 == _match_key_bytes_7_T[6:0] ? phv_data_37 : _GEN_44; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_46 = 7'h26 == _match_key_bytes_7_T[6:0] ? phv_data_38 : _GEN_45; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_47 = 7'h27 == _match_key_bytes_7_T[6:0] ? phv_data_39 : _GEN_46; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_48 = 7'h28 == _match_key_bytes_7_T[6:0] ? phv_data_40 : _GEN_47; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_49 = 7'h29 == _match_key_bytes_7_T[6:0] ? phv_data_41 : _GEN_48; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_50 = 7'h2a == _match_key_bytes_7_T[6:0] ? phv_data_42 : _GEN_49; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_51 = 7'h2b == _match_key_bytes_7_T[6:0] ? phv_data_43 : _GEN_50; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_52 = 7'h2c == _match_key_bytes_7_T[6:0] ? phv_data_44 : _GEN_51; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_53 = 7'h2d == _match_key_bytes_7_T[6:0] ? phv_data_45 : _GEN_52; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_54 = 7'h2e == _match_key_bytes_7_T[6:0] ? phv_data_46 : _GEN_53; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_55 = 7'h2f == _match_key_bytes_7_T[6:0] ? phv_data_47 : _GEN_54; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_56 = 7'h30 == _match_key_bytes_7_T[6:0] ? phv_data_48 : _GEN_55; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_57 = 7'h31 == _match_key_bytes_7_T[6:0] ? phv_data_49 : _GEN_56; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_58 = 7'h32 == _match_key_bytes_7_T[6:0] ? phv_data_50 : _GEN_57; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_59 = 7'h33 == _match_key_bytes_7_T[6:0] ? phv_data_51 : _GEN_58; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_60 = 7'h34 == _match_key_bytes_7_T[6:0] ? phv_data_52 : _GEN_59; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_61 = 7'h35 == _match_key_bytes_7_T[6:0] ? phv_data_53 : _GEN_60; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_62 = 7'h36 == _match_key_bytes_7_T[6:0] ? phv_data_54 : _GEN_61; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_63 = 7'h37 == _match_key_bytes_7_T[6:0] ? phv_data_55 : _GEN_62; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_64 = 7'h38 == _match_key_bytes_7_T[6:0] ? phv_data_56 : _GEN_63; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_65 = 7'h39 == _match_key_bytes_7_T[6:0] ? phv_data_57 : _GEN_64; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_66 = 7'h3a == _match_key_bytes_7_T[6:0] ? phv_data_58 : _GEN_65; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_67 = 7'h3b == _match_key_bytes_7_T[6:0] ? phv_data_59 : _GEN_66; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_68 = 7'h3c == _match_key_bytes_7_T[6:0] ? phv_data_60 : _GEN_67; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_69 = 7'h3d == _match_key_bytes_7_T[6:0] ? phv_data_61 : _GEN_68; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_70 = 7'h3e == _match_key_bytes_7_T[6:0] ? phv_data_62 : _GEN_69; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_71 = 7'h3f == _match_key_bytes_7_T[6:0] ? phv_data_63 : _GEN_70; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_72 = 7'h40 == _match_key_bytes_7_T[6:0] ? phv_data_64 : _GEN_71; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_73 = 7'h41 == _match_key_bytes_7_T[6:0] ? phv_data_65 : _GEN_72; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_74 = 7'h42 == _match_key_bytes_7_T[6:0] ? phv_data_66 : _GEN_73; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_75 = 7'h43 == _match_key_bytes_7_T[6:0] ? phv_data_67 : _GEN_74; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_76 = 7'h44 == _match_key_bytes_7_T[6:0] ? phv_data_68 : _GEN_75; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_77 = 7'h45 == _match_key_bytes_7_T[6:0] ? phv_data_69 : _GEN_76; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_78 = 7'h46 == _match_key_bytes_7_T[6:0] ? phv_data_70 : _GEN_77; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_79 = 7'h47 == _match_key_bytes_7_T[6:0] ? phv_data_71 : _GEN_78; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_80 = 7'h48 == _match_key_bytes_7_T[6:0] ? phv_data_72 : _GEN_79; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_81 = 7'h49 == _match_key_bytes_7_T[6:0] ? phv_data_73 : _GEN_80; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_82 = 7'h4a == _match_key_bytes_7_T[6:0] ? phv_data_74 : _GEN_81; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_83 = 7'h4b == _match_key_bytes_7_T[6:0] ? phv_data_75 : _GEN_82; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_84 = 7'h4c == _match_key_bytes_7_T[6:0] ? phv_data_76 : _GEN_83; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_85 = 7'h4d == _match_key_bytes_7_T[6:0] ? phv_data_77 : _GEN_84; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_86 = 7'h4e == _match_key_bytes_7_T[6:0] ? phv_data_78 : _GEN_85; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_87 = 7'h4f == _match_key_bytes_7_T[6:0] ? phv_data_79 : _GEN_86; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_88 = 7'h50 == _match_key_bytes_7_T[6:0] ? phv_data_80 : _GEN_87; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_89 = 7'h51 == _match_key_bytes_7_T[6:0] ? phv_data_81 : _GEN_88; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_90 = 7'h52 == _match_key_bytes_7_T[6:0] ? phv_data_82 : _GEN_89; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_91 = 7'h53 == _match_key_bytes_7_T[6:0] ? phv_data_83 : _GEN_90; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_92 = 7'h54 == _match_key_bytes_7_T[6:0] ? phv_data_84 : _GEN_91; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_93 = 7'h55 == _match_key_bytes_7_T[6:0] ? phv_data_85 : _GEN_92; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_94 = 7'h56 == _match_key_bytes_7_T[6:0] ? phv_data_86 : _GEN_93; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_95 = 7'h57 == _match_key_bytes_7_T[6:0] ? phv_data_87 : _GEN_94; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_96 = 7'h58 == _match_key_bytes_7_T[6:0] ? phv_data_88 : _GEN_95; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_97 = 7'h59 == _match_key_bytes_7_T[6:0] ? phv_data_89 : _GEN_96; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_98 = 7'h5a == _match_key_bytes_7_T[6:0] ? phv_data_90 : _GEN_97; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_99 = 7'h5b == _match_key_bytes_7_T[6:0] ? phv_data_91 : _GEN_98; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_100 = 7'h5c == _match_key_bytes_7_T[6:0] ? phv_data_92 : _GEN_99; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_101 = 7'h5d == _match_key_bytes_7_T[6:0] ? phv_data_93 : _GEN_100; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_102 = 7'h5e == _match_key_bytes_7_T[6:0] ? phv_data_94 : _GEN_101; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_103 = 7'h5f == _match_key_bytes_7_T[6:0] ? phv_data_95 : _GEN_102; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_7 = 4'h0 < _GEN_6 ? _GEN_103 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_6_T_1 = key_offset + 8'h1; // @[matcher.scala 72:98]
  wire [7:0] _GEN_106 = 7'h1 == _match_key_bytes_6_T_1[6:0] ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_107 = 7'h2 == _match_key_bytes_6_T_1[6:0] ? phv_data_2 : _GEN_106; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_108 = 7'h3 == _match_key_bytes_6_T_1[6:0] ? phv_data_3 : _GEN_107; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_109 = 7'h4 == _match_key_bytes_6_T_1[6:0] ? phv_data_4 : _GEN_108; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_110 = 7'h5 == _match_key_bytes_6_T_1[6:0] ? phv_data_5 : _GEN_109; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_111 = 7'h6 == _match_key_bytes_6_T_1[6:0] ? phv_data_6 : _GEN_110; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_112 = 7'h7 == _match_key_bytes_6_T_1[6:0] ? phv_data_7 : _GEN_111; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_113 = 7'h8 == _match_key_bytes_6_T_1[6:0] ? phv_data_8 : _GEN_112; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_114 = 7'h9 == _match_key_bytes_6_T_1[6:0] ? phv_data_9 : _GEN_113; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_115 = 7'ha == _match_key_bytes_6_T_1[6:0] ? phv_data_10 : _GEN_114; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_116 = 7'hb == _match_key_bytes_6_T_1[6:0] ? phv_data_11 : _GEN_115; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_117 = 7'hc == _match_key_bytes_6_T_1[6:0] ? phv_data_12 : _GEN_116; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_118 = 7'hd == _match_key_bytes_6_T_1[6:0] ? phv_data_13 : _GEN_117; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_119 = 7'he == _match_key_bytes_6_T_1[6:0] ? phv_data_14 : _GEN_118; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_120 = 7'hf == _match_key_bytes_6_T_1[6:0] ? phv_data_15 : _GEN_119; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_121 = 7'h10 == _match_key_bytes_6_T_1[6:0] ? phv_data_16 : _GEN_120; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_122 = 7'h11 == _match_key_bytes_6_T_1[6:0] ? phv_data_17 : _GEN_121; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_123 = 7'h12 == _match_key_bytes_6_T_1[6:0] ? phv_data_18 : _GEN_122; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_124 = 7'h13 == _match_key_bytes_6_T_1[6:0] ? phv_data_19 : _GEN_123; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_125 = 7'h14 == _match_key_bytes_6_T_1[6:0] ? phv_data_20 : _GEN_124; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_126 = 7'h15 == _match_key_bytes_6_T_1[6:0] ? phv_data_21 : _GEN_125; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_127 = 7'h16 == _match_key_bytes_6_T_1[6:0] ? phv_data_22 : _GEN_126; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_128 = 7'h17 == _match_key_bytes_6_T_1[6:0] ? phv_data_23 : _GEN_127; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_129 = 7'h18 == _match_key_bytes_6_T_1[6:0] ? phv_data_24 : _GEN_128; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_130 = 7'h19 == _match_key_bytes_6_T_1[6:0] ? phv_data_25 : _GEN_129; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_131 = 7'h1a == _match_key_bytes_6_T_1[6:0] ? phv_data_26 : _GEN_130; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_132 = 7'h1b == _match_key_bytes_6_T_1[6:0] ? phv_data_27 : _GEN_131; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_133 = 7'h1c == _match_key_bytes_6_T_1[6:0] ? phv_data_28 : _GEN_132; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_134 = 7'h1d == _match_key_bytes_6_T_1[6:0] ? phv_data_29 : _GEN_133; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_135 = 7'h1e == _match_key_bytes_6_T_1[6:0] ? phv_data_30 : _GEN_134; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_136 = 7'h1f == _match_key_bytes_6_T_1[6:0] ? phv_data_31 : _GEN_135; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_137 = 7'h20 == _match_key_bytes_6_T_1[6:0] ? phv_data_32 : _GEN_136; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_138 = 7'h21 == _match_key_bytes_6_T_1[6:0] ? phv_data_33 : _GEN_137; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_139 = 7'h22 == _match_key_bytes_6_T_1[6:0] ? phv_data_34 : _GEN_138; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_140 = 7'h23 == _match_key_bytes_6_T_1[6:0] ? phv_data_35 : _GEN_139; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_141 = 7'h24 == _match_key_bytes_6_T_1[6:0] ? phv_data_36 : _GEN_140; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_142 = 7'h25 == _match_key_bytes_6_T_1[6:0] ? phv_data_37 : _GEN_141; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_143 = 7'h26 == _match_key_bytes_6_T_1[6:0] ? phv_data_38 : _GEN_142; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_144 = 7'h27 == _match_key_bytes_6_T_1[6:0] ? phv_data_39 : _GEN_143; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_145 = 7'h28 == _match_key_bytes_6_T_1[6:0] ? phv_data_40 : _GEN_144; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_146 = 7'h29 == _match_key_bytes_6_T_1[6:0] ? phv_data_41 : _GEN_145; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_147 = 7'h2a == _match_key_bytes_6_T_1[6:0] ? phv_data_42 : _GEN_146; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_148 = 7'h2b == _match_key_bytes_6_T_1[6:0] ? phv_data_43 : _GEN_147; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_149 = 7'h2c == _match_key_bytes_6_T_1[6:0] ? phv_data_44 : _GEN_148; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_150 = 7'h2d == _match_key_bytes_6_T_1[6:0] ? phv_data_45 : _GEN_149; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_151 = 7'h2e == _match_key_bytes_6_T_1[6:0] ? phv_data_46 : _GEN_150; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_152 = 7'h2f == _match_key_bytes_6_T_1[6:0] ? phv_data_47 : _GEN_151; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_153 = 7'h30 == _match_key_bytes_6_T_1[6:0] ? phv_data_48 : _GEN_152; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_154 = 7'h31 == _match_key_bytes_6_T_1[6:0] ? phv_data_49 : _GEN_153; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_155 = 7'h32 == _match_key_bytes_6_T_1[6:0] ? phv_data_50 : _GEN_154; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_156 = 7'h33 == _match_key_bytes_6_T_1[6:0] ? phv_data_51 : _GEN_155; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_157 = 7'h34 == _match_key_bytes_6_T_1[6:0] ? phv_data_52 : _GEN_156; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_158 = 7'h35 == _match_key_bytes_6_T_1[6:0] ? phv_data_53 : _GEN_157; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_159 = 7'h36 == _match_key_bytes_6_T_1[6:0] ? phv_data_54 : _GEN_158; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_160 = 7'h37 == _match_key_bytes_6_T_1[6:0] ? phv_data_55 : _GEN_159; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_161 = 7'h38 == _match_key_bytes_6_T_1[6:0] ? phv_data_56 : _GEN_160; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_162 = 7'h39 == _match_key_bytes_6_T_1[6:0] ? phv_data_57 : _GEN_161; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_163 = 7'h3a == _match_key_bytes_6_T_1[6:0] ? phv_data_58 : _GEN_162; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_164 = 7'h3b == _match_key_bytes_6_T_1[6:0] ? phv_data_59 : _GEN_163; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_165 = 7'h3c == _match_key_bytes_6_T_1[6:0] ? phv_data_60 : _GEN_164; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_166 = 7'h3d == _match_key_bytes_6_T_1[6:0] ? phv_data_61 : _GEN_165; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_167 = 7'h3e == _match_key_bytes_6_T_1[6:0] ? phv_data_62 : _GEN_166; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_168 = 7'h3f == _match_key_bytes_6_T_1[6:0] ? phv_data_63 : _GEN_167; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_169 = 7'h40 == _match_key_bytes_6_T_1[6:0] ? phv_data_64 : _GEN_168; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_170 = 7'h41 == _match_key_bytes_6_T_1[6:0] ? phv_data_65 : _GEN_169; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_171 = 7'h42 == _match_key_bytes_6_T_1[6:0] ? phv_data_66 : _GEN_170; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_172 = 7'h43 == _match_key_bytes_6_T_1[6:0] ? phv_data_67 : _GEN_171; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_173 = 7'h44 == _match_key_bytes_6_T_1[6:0] ? phv_data_68 : _GEN_172; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_174 = 7'h45 == _match_key_bytes_6_T_1[6:0] ? phv_data_69 : _GEN_173; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_175 = 7'h46 == _match_key_bytes_6_T_1[6:0] ? phv_data_70 : _GEN_174; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_176 = 7'h47 == _match_key_bytes_6_T_1[6:0] ? phv_data_71 : _GEN_175; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_177 = 7'h48 == _match_key_bytes_6_T_1[6:0] ? phv_data_72 : _GEN_176; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_178 = 7'h49 == _match_key_bytes_6_T_1[6:0] ? phv_data_73 : _GEN_177; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_179 = 7'h4a == _match_key_bytes_6_T_1[6:0] ? phv_data_74 : _GEN_178; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_180 = 7'h4b == _match_key_bytes_6_T_1[6:0] ? phv_data_75 : _GEN_179; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_181 = 7'h4c == _match_key_bytes_6_T_1[6:0] ? phv_data_76 : _GEN_180; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_182 = 7'h4d == _match_key_bytes_6_T_1[6:0] ? phv_data_77 : _GEN_181; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_183 = 7'h4e == _match_key_bytes_6_T_1[6:0] ? phv_data_78 : _GEN_182; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_184 = 7'h4f == _match_key_bytes_6_T_1[6:0] ? phv_data_79 : _GEN_183; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_185 = 7'h50 == _match_key_bytes_6_T_1[6:0] ? phv_data_80 : _GEN_184; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_186 = 7'h51 == _match_key_bytes_6_T_1[6:0] ? phv_data_81 : _GEN_185; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_187 = 7'h52 == _match_key_bytes_6_T_1[6:0] ? phv_data_82 : _GEN_186; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_188 = 7'h53 == _match_key_bytes_6_T_1[6:0] ? phv_data_83 : _GEN_187; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_189 = 7'h54 == _match_key_bytes_6_T_1[6:0] ? phv_data_84 : _GEN_188; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_190 = 7'h55 == _match_key_bytes_6_T_1[6:0] ? phv_data_85 : _GEN_189; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_191 = 7'h56 == _match_key_bytes_6_T_1[6:0] ? phv_data_86 : _GEN_190; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_192 = 7'h57 == _match_key_bytes_6_T_1[6:0] ? phv_data_87 : _GEN_191; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_193 = 7'h58 == _match_key_bytes_6_T_1[6:0] ? phv_data_88 : _GEN_192; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_194 = 7'h59 == _match_key_bytes_6_T_1[6:0] ? phv_data_89 : _GEN_193; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_195 = 7'h5a == _match_key_bytes_6_T_1[6:0] ? phv_data_90 : _GEN_194; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_196 = 7'h5b == _match_key_bytes_6_T_1[6:0] ? phv_data_91 : _GEN_195; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_197 = 7'h5c == _match_key_bytes_6_T_1[6:0] ? phv_data_92 : _GEN_196; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_198 = 7'h5d == _match_key_bytes_6_T_1[6:0] ? phv_data_93 : _GEN_197; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_199 = 7'h5e == _match_key_bytes_6_T_1[6:0] ? phv_data_94 : _GEN_198; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_200 = 7'h5f == _match_key_bytes_6_T_1[6:0] ? phv_data_95 : _GEN_199; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_6 = 4'h1 < _GEN_6 ? _GEN_200 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_5_T_1 = key_offset + 8'h2; // @[matcher.scala 72:98]
  wire [7:0] _GEN_203 = 7'h1 == _match_key_bytes_5_T_1[6:0] ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_204 = 7'h2 == _match_key_bytes_5_T_1[6:0] ? phv_data_2 : _GEN_203; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_205 = 7'h3 == _match_key_bytes_5_T_1[6:0] ? phv_data_3 : _GEN_204; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_206 = 7'h4 == _match_key_bytes_5_T_1[6:0] ? phv_data_4 : _GEN_205; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_207 = 7'h5 == _match_key_bytes_5_T_1[6:0] ? phv_data_5 : _GEN_206; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_208 = 7'h6 == _match_key_bytes_5_T_1[6:0] ? phv_data_6 : _GEN_207; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_209 = 7'h7 == _match_key_bytes_5_T_1[6:0] ? phv_data_7 : _GEN_208; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_210 = 7'h8 == _match_key_bytes_5_T_1[6:0] ? phv_data_8 : _GEN_209; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_211 = 7'h9 == _match_key_bytes_5_T_1[6:0] ? phv_data_9 : _GEN_210; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_212 = 7'ha == _match_key_bytes_5_T_1[6:0] ? phv_data_10 : _GEN_211; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_213 = 7'hb == _match_key_bytes_5_T_1[6:0] ? phv_data_11 : _GEN_212; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_214 = 7'hc == _match_key_bytes_5_T_1[6:0] ? phv_data_12 : _GEN_213; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_215 = 7'hd == _match_key_bytes_5_T_1[6:0] ? phv_data_13 : _GEN_214; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_216 = 7'he == _match_key_bytes_5_T_1[6:0] ? phv_data_14 : _GEN_215; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_217 = 7'hf == _match_key_bytes_5_T_1[6:0] ? phv_data_15 : _GEN_216; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_218 = 7'h10 == _match_key_bytes_5_T_1[6:0] ? phv_data_16 : _GEN_217; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_219 = 7'h11 == _match_key_bytes_5_T_1[6:0] ? phv_data_17 : _GEN_218; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_220 = 7'h12 == _match_key_bytes_5_T_1[6:0] ? phv_data_18 : _GEN_219; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_221 = 7'h13 == _match_key_bytes_5_T_1[6:0] ? phv_data_19 : _GEN_220; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_222 = 7'h14 == _match_key_bytes_5_T_1[6:0] ? phv_data_20 : _GEN_221; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_223 = 7'h15 == _match_key_bytes_5_T_1[6:0] ? phv_data_21 : _GEN_222; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_224 = 7'h16 == _match_key_bytes_5_T_1[6:0] ? phv_data_22 : _GEN_223; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_225 = 7'h17 == _match_key_bytes_5_T_1[6:0] ? phv_data_23 : _GEN_224; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_226 = 7'h18 == _match_key_bytes_5_T_1[6:0] ? phv_data_24 : _GEN_225; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_227 = 7'h19 == _match_key_bytes_5_T_1[6:0] ? phv_data_25 : _GEN_226; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_228 = 7'h1a == _match_key_bytes_5_T_1[6:0] ? phv_data_26 : _GEN_227; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_229 = 7'h1b == _match_key_bytes_5_T_1[6:0] ? phv_data_27 : _GEN_228; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_230 = 7'h1c == _match_key_bytes_5_T_1[6:0] ? phv_data_28 : _GEN_229; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_231 = 7'h1d == _match_key_bytes_5_T_1[6:0] ? phv_data_29 : _GEN_230; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_232 = 7'h1e == _match_key_bytes_5_T_1[6:0] ? phv_data_30 : _GEN_231; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_233 = 7'h1f == _match_key_bytes_5_T_1[6:0] ? phv_data_31 : _GEN_232; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_234 = 7'h20 == _match_key_bytes_5_T_1[6:0] ? phv_data_32 : _GEN_233; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_235 = 7'h21 == _match_key_bytes_5_T_1[6:0] ? phv_data_33 : _GEN_234; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_236 = 7'h22 == _match_key_bytes_5_T_1[6:0] ? phv_data_34 : _GEN_235; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_237 = 7'h23 == _match_key_bytes_5_T_1[6:0] ? phv_data_35 : _GEN_236; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_238 = 7'h24 == _match_key_bytes_5_T_1[6:0] ? phv_data_36 : _GEN_237; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_239 = 7'h25 == _match_key_bytes_5_T_1[6:0] ? phv_data_37 : _GEN_238; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_240 = 7'h26 == _match_key_bytes_5_T_1[6:0] ? phv_data_38 : _GEN_239; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_241 = 7'h27 == _match_key_bytes_5_T_1[6:0] ? phv_data_39 : _GEN_240; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_242 = 7'h28 == _match_key_bytes_5_T_1[6:0] ? phv_data_40 : _GEN_241; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_243 = 7'h29 == _match_key_bytes_5_T_1[6:0] ? phv_data_41 : _GEN_242; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_244 = 7'h2a == _match_key_bytes_5_T_1[6:0] ? phv_data_42 : _GEN_243; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_245 = 7'h2b == _match_key_bytes_5_T_1[6:0] ? phv_data_43 : _GEN_244; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_246 = 7'h2c == _match_key_bytes_5_T_1[6:0] ? phv_data_44 : _GEN_245; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_247 = 7'h2d == _match_key_bytes_5_T_1[6:0] ? phv_data_45 : _GEN_246; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_248 = 7'h2e == _match_key_bytes_5_T_1[6:0] ? phv_data_46 : _GEN_247; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_249 = 7'h2f == _match_key_bytes_5_T_1[6:0] ? phv_data_47 : _GEN_248; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_250 = 7'h30 == _match_key_bytes_5_T_1[6:0] ? phv_data_48 : _GEN_249; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_251 = 7'h31 == _match_key_bytes_5_T_1[6:0] ? phv_data_49 : _GEN_250; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_252 = 7'h32 == _match_key_bytes_5_T_1[6:0] ? phv_data_50 : _GEN_251; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_253 = 7'h33 == _match_key_bytes_5_T_1[6:0] ? phv_data_51 : _GEN_252; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_254 = 7'h34 == _match_key_bytes_5_T_1[6:0] ? phv_data_52 : _GEN_253; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_255 = 7'h35 == _match_key_bytes_5_T_1[6:0] ? phv_data_53 : _GEN_254; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_256 = 7'h36 == _match_key_bytes_5_T_1[6:0] ? phv_data_54 : _GEN_255; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_257 = 7'h37 == _match_key_bytes_5_T_1[6:0] ? phv_data_55 : _GEN_256; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_258 = 7'h38 == _match_key_bytes_5_T_1[6:0] ? phv_data_56 : _GEN_257; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_259 = 7'h39 == _match_key_bytes_5_T_1[6:0] ? phv_data_57 : _GEN_258; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_260 = 7'h3a == _match_key_bytes_5_T_1[6:0] ? phv_data_58 : _GEN_259; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_261 = 7'h3b == _match_key_bytes_5_T_1[6:0] ? phv_data_59 : _GEN_260; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_262 = 7'h3c == _match_key_bytes_5_T_1[6:0] ? phv_data_60 : _GEN_261; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_263 = 7'h3d == _match_key_bytes_5_T_1[6:0] ? phv_data_61 : _GEN_262; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_264 = 7'h3e == _match_key_bytes_5_T_1[6:0] ? phv_data_62 : _GEN_263; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_265 = 7'h3f == _match_key_bytes_5_T_1[6:0] ? phv_data_63 : _GEN_264; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_266 = 7'h40 == _match_key_bytes_5_T_1[6:0] ? phv_data_64 : _GEN_265; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_267 = 7'h41 == _match_key_bytes_5_T_1[6:0] ? phv_data_65 : _GEN_266; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_268 = 7'h42 == _match_key_bytes_5_T_1[6:0] ? phv_data_66 : _GEN_267; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_269 = 7'h43 == _match_key_bytes_5_T_1[6:0] ? phv_data_67 : _GEN_268; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_270 = 7'h44 == _match_key_bytes_5_T_1[6:0] ? phv_data_68 : _GEN_269; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_271 = 7'h45 == _match_key_bytes_5_T_1[6:0] ? phv_data_69 : _GEN_270; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_272 = 7'h46 == _match_key_bytes_5_T_1[6:0] ? phv_data_70 : _GEN_271; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_273 = 7'h47 == _match_key_bytes_5_T_1[6:0] ? phv_data_71 : _GEN_272; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_274 = 7'h48 == _match_key_bytes_5_T_1[6:0] ? phv_data_72 : _GEN_273; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_275 = 7'h49 == _match_key_bytes_5_T_1[6:0] ? phv_data_73 : _GEN_274; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_276 = 7'h4a == _match_key_bytes_5_T_1[6:0] ? phv_data_74 : _GEN_275; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_277 = 7'h4b == _match_key_bytes_5_T_1[6:0] ? phv_data_75 : _GEN_276; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_278 = 7'h4c == _match_key_bytes_5_T_1[6:0] ? phv_data_76 : _GEN_277; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_279 = 7'h4d == _match_key_bytes_5_T_1[6:0] ? phv_data_77 : _GEN_278; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_280 = 7'h4e == _match_key_bytes_5_T_1[6:0] ? phv_data_78 : _GEN_279; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_281 = 7'h4f == _match_key_bytes_5_T_1[6:0] ? phv_data_79 : _GEN_280; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_282 = 7'h50 == _match_key_bytes_5_T_1[6:0] ? phv_data_80 : _GEN_281; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_283 = 7'h51 == _match_key_bytes_5_T_1[6:0] ? phv_data_81 : _GEN_282; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_284 = 7'h52 == _match_key_bytes_5_T_1[6:0] ? phv_data_82 : _GEN_283; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_285 = 7'h53 == _match_key_bytes_5_T_1[6:0] ? phv_data_83 : _GEN_284; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_286 = 7'h54 == _match_key_bytes_5_T_1[6:0] ? phv_data_84 : _GEN_285; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_287 = 7'h55 == _match_key_bytes_5_T_1[6:0] ? phv_data_85 : _GEN_286; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_288 = 7'h56 == _match_key_bytes_5_T_1[6:0] ? phv_data_86 : _GEN_287; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_289 = 7'h57 == _match_key_bytes_5_T_1[6:0] ? phv_data_87 : _GEN_288; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_290 = 7'h58 == _match_key_bytes_5_T_1[6:0] ? phv_data_88 : _GEN_289; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_291 = 7'h59 == _match_key_bytes_5_T_1[6:0] ? phv_data_89 : _GEN_290; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_292 = 7'h5a == _match_key_bytes_5_T_1[6:0] ? phv_data_90 : _GEN_291; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_293 = 7'h5b == _match_key_bytes_5_T_1[6:0] ? phv_data_91 : _GEN_292; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_294 = 7'h5c == _match_key_bytes_5_T_1[6:0] ? phv_data_92 : _GEN_293; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_295 = 7'h5d == _match_key_bytes_5_T_1[6:0] ? phv_data_93 : _GEN_294; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_296 = 7'h5e == _match_key_bytes_5_T_1[6:0] ? phv_data_94 : _GEN_295; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_297 = 7'h5f == _match_key_bytes_5_T_1[6:0] ? phv_data_95 : _GEN_296; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_5 = 4'h2 < _GEN_6 ? _GEN_297 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_4_T_1 = key_offset + 8'h3; // @[matcher.scala 72:98]
  wire [7:0] _GEN_300 = 7'h1 == _match_key_bytes_4_T_1[6:0] ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_301 = 7'h2 == _match_key_bytes_4_T_1[6:0] ? phv_data_2 : _GEN_300; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_302 = 7'h3 == _match_key_bytes_4_T_1[6:0] ? phv_data_3 : _GEN_301; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_303 = 7'h4 == _match_key_bytes_4_T_1[6:0] ? phv_data_4 : _GEN_302; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_304 = 7'h5 == _match_key_bytes_4_T_1[6:0] ? phv_data_5 : _GEN_303; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_305 = 7'h6 == _match_key_bytes_4_T_1[6:0] ? phv_data_6 : _GEN_304; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_306 = 7'h7 == _match_key_bytes_4_T_1[6:0] ? phv_data_7 : _GEN_305; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_307 = 7'h8 == _match_key_bytes_4_T_1[6:0] ? phv_data_8 : _GEN_306; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_308 = 7'h9 == _match_key_bytes_4_T_1[6:0] ? phv_data_9 : _GEN_307; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_309 = 7'ha == _match_key_bytes_4_T_1[6:0] ? phv_data_10 : _GEN_308; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_310 = 7'hb == _match_key_bytes_4_T_1[6:0] ? phv_data_11 : _GEN_309; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_311 = 7'hc == _match_key_bytes_4_T_1[6:0] ? phv_data_12 : _GEN_310; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_312 = 7'hd == _match_key_bytes_4_T_1[6:0] ? phv_data_13 : _GEN_311; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_313 = 7'he == _match_key_bytes_4_T_1[6:0] ? phv_data_14 : _GEN_312; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_314 = 7'hf == _match_key_bytes_4_T_1[6:0] ? phv_data_15 : _GEN_313; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_315 = 7'h10 == _match_key_bytes_4_T_1[6:0] ? phv_data_16 : _GEN_314; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_316 = 7'h11 == _match_key_bytes_4_T_1[6:0] ? phv_data_17 : _GEN_315; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_317 = 7'h12 == _match_key_bytes_4_T_1[6:0] ? phv_data_18 : _GEN_316; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_318 = 7'h13 == _match_key_bytes_4_T_1[6:0] ? phv_data_19 : _GEN_317; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_319 = 7'h14 == _match_key_bytes_4_T_1[6:0] ? phv_data_20 : _GEN_318; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_320 = 7'h15 == _match_key_bytes_4_T_1[6:0] ? phv_data_21 : _GEN_319; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_321 = 7'h16 == _match_key_bytes_4_T_1[6:0] ? phv_data_22 : _GEN_320; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_322 = 7'h17 == _match_key_bytes_4_T_1[6:0] ? phv_data_23 : _GEN_321; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_323 = 7'h18 == _match_key_bytes_4_T_1[6:0] ? phv_data_24 : _GEN_322; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_324 = 7'h19 == _match_key_bytes_4_T_1[6:0] ? phv_data_25 : _GEN_323; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_325 = 7'h1a == _match_key_bytes_4_T_1[6:0] ? phv_data_26 : _GEN_324; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_326 = 7'h1b == _match_key_bytes_4_T_1[6:0] ? phv_data_27 : _GEN_325; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_327 = 7'h1c == _match_key_bytes_4_T_1[6:0] ? phv_data_28 : _GEN_326; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_328 = 7'h1d == _match_key_bytes_4_T_1[6:0] ? phv_data_29 : _GEN_327; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_329 = 7'h1e == _match_key_bytes_4_T_1[6:0] ? phv_data_30 : _GEN_328; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_330 = 7'h1f == _match_key_bytes_4_T_1[6:0] ? phv_data_31 : _GEN_329; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_331 = 7'h20 == _match_key_bytes_4_T_1[6:0] ? phv_data_32 : _GEN_330; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_332 = 7'h21 == _match_key_bytes_4_T_1[6:0] ? phv_data_33 : _GEN_331; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_333 = 7'h22 == _match_key_bytes_4_T_1[6:0] ? phv_data_34 : _GEN_332; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_334 = 7'h23 == _match_key_bytes_4_T_1[6:0] ? phv_data_35 : _GEN_333; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_335 = 7'h24 == _match_key_bytes_4_T_1[6:0] ? phv_data_36 : _GEN_334; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_336 = 7'h25 == _match_key_bytes_4_T_1[6:0] ? phv_data_37 : _GEN_335; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_337 = 7'h26 == _match_key_bytes_4_T_1[6:0] ? phv_data_38 : _GEN_336; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_338 = 7'h27 == _match_key_bytes_4_T_1[6:0] ? phv_data_39 : _GEN_337; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_339 = 7'h28 == _match_key_bytes_4_T_1[6:0] ? phv_data_40 : _GEN_338; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_340 = 7'h29 == _match_key_bytes_4_T_1[6:0] ? phv_data_41 : _GEN_339; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_341 = 7'h2a == _match_key_bytes_4_T_1[6:0] ? phv_data_42 : _GEN_340; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_342 = 7'h2b == _match_key_bytes_4_T_1[6:0] ? phv_data_43 : _GEN_341; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_343 = 7'h2c == _match_key_bytes_4_T_1[6:0] ? phv_data_44 : _GEN_342; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_344 = 7'h2d == _match_key_bytes_4_T_1[6:0] ? phv_data_45 : _GEN_343; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_345 = 7'h2e == _match_key_bytes_4_T_1[6:0] ? phv_data_46 : _GEN_344; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_346 = 7'h2f == _match_key_bytes_4_T_1[6:0] ? phv_data_47 : _GEN_345; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_347 = 7'h30 == _match_key_bytes_4_T_1[6:0] ? phv_data_48 : _GEN_346; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_348 = 7'h31 == _match_key_bytes_4_T_1[6:0] ? phv_data_49 : _GEN_347; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_349 = 7'h32 == _match_key_bytes_4_T_1[6:0] ? phv_data_50 : _GEN_348; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_350 = 7'h33 == _match_key_bytes_4_T_1[6:0] ? phv_data_51 : _GEN_349; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_351 = 7'h34 == _match_key_bytes_4_T_1[6:0] ? phv_data_52 : _GEN_350; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_352 = 7'h35 == _match_key_bytes_4_T_1[6:0] ? phv_data_53 : _GEN_351; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_353 = 7'h36 == _match_key_bytes_4_T_1[6:0] ? phv_data_54 : _GEN_352; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_354 = 7'h37 == _match_key_bytes_4_T_1[6:0] ? phv_data_55 : _GEN_353; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_355 = 7'h38 == _match_key_bytes_4_T_1[6:0] ? phv_data_56 : _GEN_354; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_356 = 7'h39 == _match_key_bytes_4_T_1[6:0] ? phv_data_57 : _GEN_355; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_357 = 7'h3a == _match_key_bytes_4_T_1[6:0] ? phv_data_58 : _GEN_356; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_358 = 7'h3b == _match_key_bytes_4_T_1[6:0] ? phv_data_59 : _GEN_357; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_359 = 7'h3c == _match_key_bytes_4_T_1[6:0] ? phv_data_60 : _GEN_358; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_360 = 7'h3d == _match_key_bytes_4_T_1[6:0] ? phv_data_61 : _GEN_359; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_361 = 7'h3e == _match_key_bytes_4_T_1[6:0] ? phv_data_62 : _GEN_360; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_362 = 7'h3f == _match_key_bytes_4_T_1[6:0] ? phv_data_63 : _GEN_361; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_363 = 7'h40 == _match_key_bytes_4_T_1[6:0] ? phv_data_64 : _GEN_362; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_364 = 7'h41 == _match_key_bytes_4_T_1[6:0] ? phv_data_65 : _GEN_363; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_365 = 7'h42 == _match_key_bytes_4_T_1[6:0] ? phv_data_66 : _GEN_364; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_366 = 7'h43 == _match_key_bytes_4_T_1[6:0] ? phv_data_67 : _GEN_365; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_367 = 7'h44 == _match_key_bytes_4_T_1[6:0] ? phv_data_68 : _GEN_366; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_368 = 7'h45 == _match_key_bytes_4_T_1[6:0] ? phv_data_69 : _GEN_367; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_369 = 7'h46 == _match_key_bytes_4_T_1[6:0] ? phv_data_70 : _GEN_368; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_370 = 7'h47 == _match_key_bytes_4_T_1[6:0] ? phv_data_71 : _GEN_369; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_371 = 7'h48 == _match_key_bytes_4_T_1[6:0] ? phv_data_72 : _GEN_370; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_372 = 7'h49 == _match_key_bytes_4_T_1[6:0] ? phv_data_73 : _GEN_371; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_373 = 7'h4a == _match_key_bytes_4_T_1[6:0] ? phv_data_74 : _GEN_372; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_374 = 7'h4b == _match_key_bytes_4_T_1[6:0] ? phv_data_75 : _GEN_373; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_375 = 7'h4c == _match_key_bytes_4_T_1[6:0] ? phv_data_76 : _GEN_374; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_376 = 7'h4d == _match_key_bytes_4_T_1[6:0] ? phv_data_77 : _GEN_375; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_377 = 7'h4e == _match_key_bytes_4_T_1[6:0] ? phv_data_78 : _GEN_376; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_378 = 7'h4f == _match_key_bytes_4_T_1[6:0] ? phv_data_79 : _GEN_377; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_379 = 7'h50 == _match_key_bytes_4_T_1[6:0] ? phv_data_80 : _GEN_378; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_380 = 7'h51 == _match_key_bytes_4_T_1[6:0] ? phv_data_81 : _GEN_379; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_381 = 7'h52 == _match_key_bytes_4_T_1[6:0] ? phv_data_82 : _GEN_380; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_382 = 7'h53 == _match_key_bytes_4_T_1[6:0] ? phv_data_83 : _GEN_381; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_383 = 7'h54 == _match_key_bytes_4_T_1[6:0] ? phv_data_84 : _GEN_382; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_384 = 7'h55 == _match_key_bytes_4_T_1[6:0] ? phv_data_85 : _GEN_383; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_385 = 7'h56 == _match_key_bytes_4_T_1[6:0] ? phv_data_86 : _GEN_384; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_386 = 7'h57 == _match_key_bytes_4_T_1[6:0] ? phv_data_87 : _GEN_385; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_387 = 7'h58 == _match_key_bytes_4_T_1[6:0] ? phv_data_88 : _GEN_386; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_388 = 7'h59 == _match_key_bytes_4_T_1[6:0] ? phv_data_89 : _GEN_387; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_389 = 7'h5a == _match_key_bytes_4_T_1[6:0] ? phv_data_90 : _GEN_388; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_390 = 7'h5b == _match_key_bytes_4_T_1[6:0] ? phv_data_91 : _GEN_389; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_391 = 7'h5c == _match_key_bytes_4_T_1[6:0] ? phv_data_92 : _GEN_390; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_392 = 7'h5d == _match_key_bytes_4_T_1[6:0] ? phv_data_93 : _GEN_391; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_393 = 7'h5e == _match_key_bytes_4_T_1[6:0] ? phv_data_94 : _GEN_392; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_394 = 7'h5f == _match_key_bytes_4_T_1[6:0] ? phv_data_95 : _GEN_393; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_4 = 4'h3 < _GEN_6 ? _GEN_394 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_3_T_1 = key_offset + 8'h4; // @[matcher.scala 72:98]
  wire [7:0] _GEN_397 = 7'h1 == _match_key_bytes_3_T_1[6:0] ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_398 = 7'h2 == _match_key_bytes_3_T_1[6:0] ? phv_data_2 : _GEN_397; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_399 = 7'h3 == _match_key_bytes_3_T_1[6:0] ? phv_data_3 : _GEN_398; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_400 = 7'h4 == _match_key_bytes_3_T_1[6:0] ? phv_data_4 : _GEN_399; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_401 = 7'h5 == _match_key_bytes_3_T_1[6:0] ? phv_data_5 : _GEN_400; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_402 = 7'h6 == _match_key_bytes_3_T_1[6:0] ? phv_data_6 : _GEN_401; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_403 = 7'h7 == _match_key_bytes_3_T_1[6:0] ? phv_data_7 : _GEN_402; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_404 = 7'h8 == _match_key_bytes_3_T_1[6:0] ? phv_data_8 : _GEN_403; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_405 = 7'h9 == _match_key_bytes_3_T_1[6:0] ? phv_data_9 : _GEN_404; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_406 = 7'ha == _match_key_bytes_3_T_1[6:0] ? phv_data_10 : _GEN_405; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_407 = 7'hb == _match_key_bytes_3_T_1[6:0] ? phv_data_11 : _GEN_406; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_408 = 7'hc == _match_key_bytes_3_T_1[6:0] ? phv_data_12 : _GEN_407; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_409 = 7'hd == _match_key_bytes_3_T_1[6:0] ? phv_data_13 : _GEN_408; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_410 = 7'he == _match_key_bytes_3_T_1[6:0] ? phv_data_14 : _GEN_409; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_411 = 7'hf == _match_key_bytes_3_T_1[6:0] ? phv_data_15 : _GEN_410; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_412 = 7'h10 == _match_key_bytes_3_T_1[6:0] ? phv_data_16 : _GEN_411; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_413 = 7'h11 == _match_key_bytes_3_T_1[6:0] ? phv_data_17 : _GEN_412; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_414 = 7'h12 == _match_key_bytes_3_T_1[6:0] ? phv_data_18 : _GEN_413; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_415 = 7'h13 == _match_key_bytes_3_T_1[6:0] ? phv_data_19 : _GEN_414; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_416 = 7'h14 == _match_key_bytes_3_T_1[6:0] ? phv_data_20 : _GEN_415; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_417 = 7'h15 == _match_key_bytes_3_T_1[6:0] ? phv_data_21 : _GEN_416; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_418 = 7'h16 == _match_key_bytes_3_T_1[6:0] ? phv_data_22 : _GEN_417; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_419 = 7'h17 == _match_key_bytes_3_T_1[6:0] ? phv_data_23 : _GEN_418; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_420 = 7'h18 == _match_key_bytes_3_T_1[6:0] ? phv_data_24 : _GEN_419; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_421 = 7'h19 == _match_key_bytes_3_T_1[6:0] ? phv_data_25 : _GEN_420; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_422 = 7'h1a == _match_key_bytes_3_T_1[6:0] ? phv_data_26 : _GEN_421; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_423 = 7'h1b == _match_key_bytes_3_T_1[6:0] ? phv_data_27 : _GEN_422; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_424 = 7'h1c == _match_key_bytes_3_T_1[6:0] ? phv_data_28 : _GEN_423; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_425 = 7'h1d == _match_key_bytes_3_T_1[6:0] ? phv_data_29 : _GEN_424; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_426 = 7'h1e == _match_key_bytes_3_T_1[6:0] ? phv_data_30 : _GEN_425; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_427 = 7'h1f == _match_key_bytes_3_T_1[6:0] ? phv_data_31 : _GEN_426; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_428 = 7'h20 == _match_key_bytes_3_T_1[6:0] ? phv_data_32 : _GEN_427; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_429 = 7'h21 == _match_key_bytes_3_T_1[6:0] ? phv_data_33 : _GEN_428; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_430 = 7'h22 == _match_key_bytes_3_T_1[6:0] ? phv_data_34 : _GEN_429; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_431 = 7'h23 == _match_key_bytes_3_T_1[6:0] ? phv_data_35 : _GEN_430; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_432 = 7'h24 == _match_key_bytes_3_T_1[6:0] ? phv_data_36 : _GEN_431; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_433 = 7'h25 == _match_key_bytes_3_T_1[6:0] ? phv_data_37 : _GEN_432; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_434 = 7'h26 == _match_key_bytes_3_T_1[6:0] ? phv_data_38 : _GEN_433; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_435 = 7'h27 == _match_key_bytes_3_T_1[6:0] ? phv_data_39 : _GEN_434; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_436 = 7'h28 == _match_key_bytes_3_T_1[6:0] ? phv_data_40 : _GEN_435; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_437 = 7'h29 == _match_key_bytes_3_T_1[6:0] ? phv_data_41 : _GEN_436; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_438 = 7'h2a == _match_key_bytes_3_T_1[6:0] ? phv_data_42 : _GEN_437; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_439 = 7'h2b == _match_key_bytes_3_T_1[6:0] ? phv_data_43 : _GEN_438; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_440 = 7'h2c == _match_key_bytes_3_T_1[6:0] ? phv_data_44 : _GEN_439; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_441 = 7'h2d == _match_key_bytes_3_T_1[6:0] ? phv_data_45 : _GEN_440; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_442 = 7'h2e == _match_key_bytes_3_T_1[6:0] ? phv_data_46 : _GEN_441; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_443 = 7'h2f == _match_key_bytes_3_T_1[6:0] ? phv_data_47 : _GEN_442; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_444 = 7'h30 == _match_key_bytes_3_T_1[6:0] ? phv_data_48 : _GEN_443; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_445 = 7'h31 == _match_key_bytes_3_T_1[6:0] ? phv_data_49 : _GEN_444; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_446 = 7'h32 == _match_key_bytes_3_T_1[6:0] ? phv_data_50 : _GEN_445; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_447 = 7'h33 == _match_key_bytes_3_T_1[6:0] ? phv_data_51 : _GEN_446; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_448 = 7'h34 == _match_key_bytes_3_T_1[6:0] ? phv_data_52 : _GEN_447; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_449 = 7'h35 == _match_key_bytes_3_T_1[6:0] ? phv_data_53 : _GEN_448; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_450 = 7'h36 == _match_key_bytes_3_T_1[6:0] ? phv_data_54 : _GEN_449; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_451 = 7'h37 == _match_key_bytes_3_T_1[6:0] ? phv_data_55 : _GEN_450; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_452 = 7'h38 == _match_key_bytes_3_T_1[6:0] ? phv_data_56 : _GEN_451; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_453 = 7'h39 == _match_key_bytes_3_T_1[6:0] ? phv_data_57 : _GEN_452; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_454 = 7'h3a == _match_key_bytes_3_T_1[6:0] ? phv_data_58 : _GEN_453; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_455 = 7'h3b == _match_key_bytes_3_T_1[6:0] ? phv_data_59 : _GEN_454; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_456 = 7'h3c == _match_key_bytes_3_T_1[6:0] ? phv_data_60 : _GEN_455; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_457 = 7'h3d == _match_key_bytes_3_T_1[6:0] ? phv_data_61 : _GEN_456; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_458 = 7'h3e == _match_key_bytes_3_T_1[6:0] ? phv_data_62 : _GEN_457; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_459 = 7'h3f == _match_key_bytes_3_T_1[6:0] ? phv_data_63 : _GEN_458; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_460 = 7'h40 == _match_key_bytes_3_T_1[6:0] ? phv_data_64 : _GEN_459; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_461 = 7'h41 == _match_key_bytes_3_T_1[6:0] ? phv_data_65 : _GEN_460; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_462 = 7'h42 == _match_key_bytes_3_T_1[6:0] ? phv_data_66 : _GEN_461; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_463 = 7'h43 == _match_key_bytes_3_T_1[6:0] ? phv_data_67 : _GEN_462; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_464 = 7'h44 == _match_key_bytes_3_T_1[6:0] ? phv_data_68 : _GEN_463; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_465 = 7'h45 == _match_key_bytes_3_T_1[6:0] ? phv_data_69 : _GEN_464; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_466 = 7'h46 == _match_key_bytes_3_T_1[6:0] ? phv_data_70 : _GEN_465; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_467 = 7'h47 == _match_key_bytes_3_T_1[6:0] ? phv_data_71 : _GEN_466; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_468 = 7'h48 == _match_key_bytes_3_T_1[6:0] ? phv_data_72 : _GEN_467; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_469 = 7'h49 == _match_key_bytes_3_T_1[6:0] ? phv_data_73 : _GEN_468; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_470 = 7'h4a == _match_key_bytes_3_T_1[6:0] ? phv_data_74 : _GEN_469; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_471 = 7'h4b == _match_key_bytes_3_T_1[6:0] ? phv_data_75 : _GEN_470; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_472 = 7'h4c == _match_key_bytes_3_T_1[6:0] ? phv_data_76 : _GEN_471; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_473 = 7'h4d == _match_key_bytes_3_T_1[6:0] ? phv_data_77 : _GEN_472; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_474 = 7'h4e == _match_key_bytes_3_T_1[6:0] ? phv_data_78 : _GEN_473; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_475 = 7'h4f == _match_key_bytes_3_T_1[6:0] ? phv_data_79 : _GEN_474; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_476 = 7'h50 == _match_key_bytes_3_T_1[6:0] ? phv_data_80 : _GEN_475; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_477 = 7'h51 == _match_key_bytes_3_T_1[6:0] ? phv_data_81 : _GEN_476; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_478 = 7'h52 == _match_key_bytes_3_T_1[6:0] ? phv_data_82 : _GEN_477; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_479 = 7'h53 == _match_key_bytes_3_T_1[6:0] ? phv_data_83 : _GEN_478; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_480 = 7'h54 == _match_key_bytes_3_T_1[6:0] ? phv_data_84 : _GEN_479; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_481 = 7'h55 == _match_key_bytes_3_T_1[6:0] ? phv_data_85 : _GEN_480; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_482 = 7'h56 == _match_key_bytes_3_T_1[6:0] ? phv_data_86 : _GEN_481; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_483 = 7'h57 == _match_key_bytes_3_T_1[6:0] ? phv_data_87 : _GEN_482; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_484 = 7'h58 == _match_key_bytes_3_T_1[6:0] ? phv_data_88 : _GEN_483; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_485 = 7'h59 == _match_key_bytes_3_T_1[6:0] ? phv_data_89 : _GEN_484; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_486 = 7'h5a == _match_key_bytes_3_T_1[6:0] ? phv_data_90 : _GEN_485; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_487 = 7'h5b == _match_key_bytes_3_T_1[6:0] ? phv_data_91 : _GEN_486; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_488 = 7'h5c == _match_key_bytes_3_T_1[6:0] ? phv_data_92 : _GEN_487; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_489 = 7'h5d == _match_key_bytes_3_T_1[6:0] ? phv_data_93 : _GEN_488; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_490 = 7'h5e == _match_key_bytes_3_T_1[6:0] ? phv_data_94 : _GEN_489; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_491 = 7'h5f == _match_key_bytes_3_T_1[6:0] ? phv_data_95 : _GEN_490; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_3 = 4'h4 < _GEN_6 ? _GEN_491 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_2_T_1 = key_offset + 8'h5; // @[matcher.scala 72:98]
  wire [7:0] _GEN_494 = 7'h1 == _match_key_bytes_2_T_1[6:0] ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_495 = 7'h2 == _match_key_bytes_2_T_1[6:0] ? phv_data_2 : _GEN_494; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_496 = 7'h3 == _match_key_bytes_2_T_1[6:0] ? phv_data_3 : _GEN_495; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_497 = 7'h4 == _match_key_bytes_2_T_1[6:0] ? phv_data_4 : _GEN_496; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_498 = 7'h5 == _match_key_bytes_2_T_1[6:0] ? phv_data_5 : _GEN_497; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_499 = 7'h6 == _match_key_bytes_2_T_1[6:0] ? phv_data_6 : _GEN_498; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_500 = 7'h7 == _match_key_bytes_2_T_1[6:0] ? phv_data_7 : _GEN_499; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_501 = 7'h8 == _match_key_bytes_2_T_1[6:0] ? phv_data_8 : _GEN_500; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_502 = 7'h9 == _match_key_bytes_2_T_1[6:0] ? phv_data_9 : _GEN_501; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_503 = 7'ha == _match_key_bytes_2_T_1[6:0] ? phv_data_10 : _GEN_502; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_504 = 7'hb == _match_key_bytes_2_T_1[6:0] ? phv_data_11 : _GEN_503; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_505 = 7'hc == _match_key_bytes_2_T_1[6:0] ? phv_data_12 : _GEN_504; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_506 = 7'hd == _match_key_bytes_2_T_1[6:0] ? phv_data_13 : _GEN_505; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_507 = 7'he == _match_key_bytes_2_T_1[6:0] ? phv_data_14 : _GEN_506; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_508 = 7'hf == _match_key_bytes_2_T_1[6:0] ? phv_data_15 : _GEN_507; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_509 = 7'h10 == _match_key_bytes_2_T_1[6:0] ? phv_data_16 : _GEN_508; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_510 = 7'h11 == _match_key_bytes_2_T_1[6:0] ? phv_data_17 : _GEN_509; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_511 = 7'h12 == _match_key_bytes_2_T_1[6:0] ? phv_data_18 : _GEN_510; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_512 = 7'h13 == _match_key_bytes_2_T_1[6:0] ? phv_data_19 : _GEN_511; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_513 = 7'h14 == _match_key_bytes_2_T_1[6:0] ? phv_data_20 : _GEN_512; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_514 = 7'h15 == _match_key_bytes_2_T_1[6:0] ? phv_data_21 : _GEN_513; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_515 = 7'h16 == _match_key_bytes_2_T_1[6:0] ? phv_data_22 : _GEN_514; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_516 = 7'h17 == _match_key_bytes_2_T_1[6:0] ? phv_data_23 : _GEN_515; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_517 = 7'h18 == _match_key_bytes_2_T_1[6:0] ? phv_data_24 : _GEN_516; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_518 = 7'h19 == _match_key_bytes_2_T_1[6:0] ? phv_data_25 : _GEN_517; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_519 = 7'h1a == _match_key_bytes_2_T_1[6:0] ? phv_data_26 : _GEN_518; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_520 = 7'h1b == _match_key_bytes_2_T_1[6:0] ? phv_data_27 : _GEN_519; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_521 = 7'h1c == _match_key_bytes_2_T_1[6:0] ? phv_data_28 : _GEN_520; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_522 = 7'h1d == _match_key_bytes_2_T_1[6:0] ? phv_data_29 : _GEN_521; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_523 = 7'h1e == _match_key_bytes_2_T_1[6:0] ? phv_data_30 : _GEN_522; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_524 = 7'h1f == _match_key_bytes_2_T_1[6:0] ? phv_data_31 : _GEN_523; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_525 = 7'h20 == _match_key_bytes_2_T_1[6:0] ? phv_data_32 : _GEN_524; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_526 = 7'h21 == _match_key_bytes_2_T_1[6:0] ? phv_data_33 : _GEN_525; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_527 = 7'h22 == _match_key_bytes_2_T_1[6:0] ? phv_data_34 : _GEN_526; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_528 = 7'h23 == _match_key_bytes_2_T_1[6:0] ? phv_data_35 : _GEN_527; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_529 = 7'h24 == _match_key_bytes_2_T_1[6:0] ? phv_data_36 : _GEN_528; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_530 = 7'h25 == _match_key_bytes_2_T_1[6:0] ? phv_data_37 : _GEN_529; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_531 = 7'h26 == _match_key_bytes_2_T_1[6:0] ? phv_data_38 : _GEN_530; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_532 = 7'h27 == _match_key_bytes_2_T_1[6:0] ? phv_data_39 : _GEN_531; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_533 = 7'h28 == _match_key_bytes_2_T_1[6:0] ? phv_data_40 : _GEN_532; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_534 = 7'h29 == _match_key_bytes_2_T_1[6:0] ? phv_data_41 : _GEN_533; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_535 = 7'h2a == _match_key_bytes_2_T_1[6:0] ? phv_data_42 : _GEN_534; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_536 = 7'h2b == _match_key_bytes_2_T_1[6:0] ? phv_data_43 : _GEN_535; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_537 = 7'h2c == _match_key_bytes_2_T_1[6:0] ? phv_data_44 : _GEN_536; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_538 = 7'h2d == _match_key_bytes_2_T_1[6:0] ? phv_data_45 : _GEN_537; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_539 = 7'h2e == _match_key_bytes_2_T_1[6:0] ? phv_data_46 : _GEN_538; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_540 = 7'h2f == _match_key_bytes_2_T_1[6:0] ? phv_data_47 : _GEN_539; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_541 = 7'h30 == _match_key_bytes_2_T_1[6:0] ? phv_data_48 : _GEN_540; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_542 = 7'h31 == _match_key_bytes_2_T_1[6:0] ? phv_data_49 : _GEN_541; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_543 = 7'h32 == _match_key_bytes_2_T_1[6:0] ? phv_data_50 : _GEN_542; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_544 = 7'h33 == _match_key_bytes_2_T_1[6:0] ? phv_data_51 : _GEN_543; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_545 = 7'h34 == _match_key_bytes_2_T_1[6:0] ? phv_data_52 : _GEN_544; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_546 = 7'h35 == _match_key_bytes_2_T_1[6:0] ? phv_data_53 : _GEN_545; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_547 = 7'h36 == _match_key_bytes_2_T_1[6:0] ? phv_data_54 : _GEN_546; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_548 = 7'h37 == _match_key_bytes_2_T_1[6:0] ? phv_data_55 : _GEN_547; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_549 = 7'h38 == _match_key_bytes_2_T_1[6:0] ? phv_data_56 : _GEN_548; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_550 = 7'h39 == _match_key_bytes_2_T_1[6:0] ? phv_data_57 : _GEN_549; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_551 = 7'h3a == _match_key_bytes_2_T_1[6:0] ? phv_data_58 : _GEN_550; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_552 = 7'h3b == _match_key_bytes_2_T_1[6:0] ? phv_data_59 : _GEN_551; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_553 = 7'h3c == _match_key_bytes_2_T_1[6:0] ? phv_data_60 : _GEN_552; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_554 = 7'h3d == _match_key_bytes_2_T_1[6:0] ? phv_data_61 : _GEN_553; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_555 = 7'h3e == _match_key_bytes_2_T_1[6:0] ? phv_data_62 : _GEN_554; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_556 = 7'h3f == _match_key_bytes_2_T_1[6:0] ? phv_data_63 : _GEN_555; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_557 = 7'h40 == _match_key_bytes_2_T_1[6:0] ? phv_data_64 : _GEN_556; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_558 = 7'h41 == _match_key_bytes_2_T_1[6:0] ? phv_data_65 : _GEN_557; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_559 = 7'h42 == _match_key_bytes_2_T_1[6:0] ? phv_data_66 : _GEN_558; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_560 = 7'h43 == _match_key_bytes_2_T_1[6:0] ? phv_data_67 : _GEN_559; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_561 = 7'h44 == _match_key_bytes_2_T_1[6:0] ? phv_data_68 : _GEN_560; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_562 = 7'h45 == _match_key_bytes_2_T_1[6:0] ? phv_data_69 : _GEN_561; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_563 = 7'h46 == _match_key_bytes_2_T_1[6:0] ? phv_data_70 : _GEN_562; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_564 = 7'h47 == _match_key_bytes_2_T_1[6:0] ? phv_data_71 : _GEN_563; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_565 = 7'h48 == _match_key_bytes_2_T_1[6:0] ? phv_data_72 : _GEN_564; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_566 = 7'h49 == _match_key_bytes_2_T_1[6:0] ? phv_data_73 : _GEN_565; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_567 = 7'h4a == _match_key_bytes_2_T_1[6:0] ? phv_data_74 : _GEN_566; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_568 = 7'h4b == _match_key_bytes_2_T_1[6:0] ? phv_data_75 : _GEN_567; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_569 = 7'h4c == _match_key_bytes_2_T_1[6:0] ? phv_data_76 : _GEN_568; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_570 = 7'h4d == _match_key_bytes_2_T_1[6:0] ? phv_data_77 : _GEN_569; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_571 = 7'h4e == _match_key_bytes_2_T_1[6:0] ? phv_data_78 : _GEN_570; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_572 = 7'h4f == _match_key_bytes_2_T_1[6:0] ? phv_data_79 : _GEN_571; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_573 = 7'h50 == _match_key_bytes_2_T_1[6:0] ? phv_data_80 : _GEN_572; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_574 = 7'h51 == _match_key_bytes_2_T_1[6:0] ? phv_data_81 : _GEN_573; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_575 = 7'h52 == _match_key_bytes_2_T_1[6:0] ? phv_data_82 : _GEN_574; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_576 = 7'h53 == _match_key_bytes_2_T_1[6:0] ? phv_data_83 : _GEN_575; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_577 = 7'h54 == _match_key_bytes_2_T_1[6:0] ? phv_data_84 : _GEN_576; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_578 = 7'h55 == _match_key_bytes_2_T_1[6:0] ? phv_data_85 : _GEN_577; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_579 = 7'h56 == _match_key_bytes_2_T_1[6:0] ? phv_data_86 : _GEN_578; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_580 = 7'h57 == _match_key_bytes_2_T_1[6:0] ? phv_data_87 : _GEN_579; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_581 = 7'h58 == _match_key_bytes_2_T_1[6:0] ? phv_data_88 : _GEN_580; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_582 = 7'h59 == _match_key_bytes_2_T_1[6:0] ? phv_data_89 : _GEN_581; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_583 = 7'h5a == _match_key_bytes_2_T_1[6:0] ? phv_data_90 : _GEN_582; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_584 = 7'h5b == _match_key_bytes_2_T_1[6:0] ? phv_data_91 : _GEN_583; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_585 = 7'h5c == _match_key_bytes_2_T_1[6:0] ? phv_data_92 : _GEN_584; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_586 = 7'h5d == _match_key_bytes_2_T_1[6:0] ? phv_data_93 : _GEN_585; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_587 = 7'h5e == _match_key_bytes_2_T_1[6:0] ? phv_data_94 : _GEN_586; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_588 = 7'h5f == _match_key_bytes_2_T_1[6:0] ? phv_data_95 : _GEN_587; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_2 = 4'h5 < _GEN_6 ? _GEN_588 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_1_T_1 = key_offset + 8'h6; // @[matcher.scala 72:98]
  wire [7:0] _GEN_591 = 7'h1 == _match_key_bytes_1_T_1[6:0] ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_592 = 7'h2 == _match_key_bytes_1_T_1[6:0] ? phv_data_2 : _GEN_591; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_593 = 7'h3 == _match_key_bytes_1_T_1[6:0] ? phv_data_3 : _GEN_592; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_594 = 7'h4 == _match_key_bytes_1_T_1[6:0] ? phv_data_4 : _GEN_593; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_595 = 7'h5 == _match_key_bytes_1_T_1[6:0] ? phv_data_5 : _GEN_594; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_596 = 7'h6 == _match_key_bytes_1_T_1[6:0] ? phv_data_6 : _GEN_595; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_597 = 7'h7 == _match_key_bytes_1_T_1[6:0] ? phv_data_7 : _GEN_596; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_598 = 7'h8 == _match_key_bytes_1_T_1[6:0] ? phv_data_8 : _GEN_597; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_599 = 7'h9 == _match_key_bytes_1_T_1[6:0] ? phv_data_9 : _GEN_598; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_600 = 7'ha == _match_key_bytes_1_T_1[6:0] ? phv_data_10 : _GEN_599; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_601 = 7'hb == _match_key_bytes_1_T_1[6:0] ? phv_data_11 : _GEN_600; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_602 = 7'hc == _match_key_bytes_1_T_1[6:0] ? phv_data_12 : _GEN_601; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_603 = 7'hd == _match_key_bytes_1_T_1[6:0] ? phv_data_13 : _GEN_602; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_604 = 7'he == _match_key_bytes_1_T_1[6:0] ? phv_data_14 : _GEN_603; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_605 = 7'hf == _match_key_bytes_1_T_1[6:0] ? phv_data_15 : _GEN_604; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_606 = 7'h10 == _match_key_bytes_1_T_1[6:0] ? phv_data_16 : _GEN_605; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_607 = 7'h11 == _match_key_bytes_1_T_1[6:0] ? phv_data_17 : _GEN_606; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_608 = 7'h12 == _match_key_bytes_1_T_1[6:0] ? phv_data_18 : _GEN_607; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_609 = 7'h13 == _match_key_bytes_1_T_1[6:0] ? phv_data_19 : _GEN_608; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_610 = 7'h14 == _match_key_bytes_1_T_1[6:0] ? phv_data_20 : _GEN_609; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_611 = 7'h15 == _match_key_bytes_1_T_1[6:0] ? phv_data_21 : _GEN_610; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_612 = 7'h16 == _match_key_bytes_1_T_1[6:0] ? phv_data_22 : _GEN_611; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_613 = 7'h17 == _match_key_bytes_1_T_1[6:0] ? phv_data_23 : _GEN_612; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_614 = 7'h18 == _match_key_bytes_1_T_1[6:0] ? phv_data_24 : _GEN_613; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_615 = 7'h19 == _match_key_bytes_1_T_1[6:0] ? phv_data_25 : _GEN_614; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_616 = 7'h1a == _match_key_bytes_1_T_1[6:0] ? phv_data_26 : _GEN_615; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_617 = 7'h1b == _match_key_bytes_1_T_1[6:0] ? phv_data_27 : _GEN_616; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_618 = 7'h1c == _match_key_bytes_1_T_1[6:0] ? phv_data_28 : _GEN_617; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_619 = 7'h1d == _match_key_bytes_1_T_1[6:0] ? phv_data_29 : _GEN_618; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_620 = 7'h1e == _match_key_bytes_1_T_1[6:0] ? phv_data_30 : _GEN_619; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_621 = 7'h1f == _match_key_bytes_1_T_1[6:0] ? phv_data_31 : _GEN_620; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_622 = 7'h20 == _match_key_bytes_1_T_1[6:0] ? phv_data_32 : _GEN_621; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_623 = 7'h21 == _match_key_bytes_1_T_1[6:0] ? phv_data_33 : _GEN_622; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_624 = 7'h22 == _match_key_bytes_1_T_1[6:0] ? phv_data_34 : _GEN_623; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_625 = 7'h23 == _match_key_bytes_1_T_1[6:0] ? phv_data_35 : _GEN_624; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_626 = 7'h24 == _match_key_bytes_1_T_1[6:0] ? phv_data_36 : _GEN_625; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_627 = 7'h25 == _match_key_bytes_1_T_1[6:0] ? phv_data_37 : _GEN_626; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_628 = 7'h26 == _match_key_bytes_1_T_1[6:0] ? phv_data_38 : _GEN_627; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_629 = 7'h27 == _match_key_bytes_1_T_1[6:0] ? phv_data_39 : _GEN_628; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_630 = 7'h28 == _match_key_bytes_1_T_1[6:0] ? phv_data_40 : _GEN_629; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_631 = 7'h29 == _match_key_bytes_1_T_1[6:0] ? phv_data_41 : _GEN_630; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_632 = 7'h2a == _match_key_bytes_1_T_1[6:0] ? phv_data_42 : _GEN_631; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_633 = 7'h2b == _match_key_bytes_1_T_1[6:0] ? phv_data_43 : _GEN_632; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_634 = 7'h2c == _match_key_bytes_1_T_1[6:0] ? phv_data_44 : _GEN_633; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_635 = 7'h2d == _match_key_bytes_1_T_1[6:0] ? phv_data_45 : _GEN_634; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_636 = 7'h2e == _match_key_bytes_1_T_1[6:0] ? phv_data_46 : _GEN_635; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_637 = 7'h2f == _match_key_bytes_1_T_1[6:0] ? phv_data_47 : _GEN_636; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_638 = 7'h30 == _match_key_bytes_1_T_1[6:0] ? phv_data_48 : _GEN_637; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_639 = 7'h31 == _match_key_bytes_1_T_1[6:0] ? phv_data_49 : _GEN_638; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_640 = 7'h32 == _match_key_bytes_1_T_1[6:0] ? phv_data_50 : _GEN_639; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_641 = 7'h33 == _match_key_bytes_1_T_1[6:0] ? phv_data_51 : _GEN_640; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_642 = 7'h34 == _match_key_bytes_1_T_1[6:0] ? phv_data_52 : _GEN_641; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_643 = 7'h35 == _match_key_bytes_1_T_1[6:0] ? phv_data_53 : _GEN_642; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_644 = 7'h36 == _match_key_bytes_1_T_1[6:0] ? phv_data_54 : _GEN_643; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_645 = 7'h37 == _match_key_bytes_1_T_1[6:0] ? phv_data_55 : _GEN_644; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_646 = 7'h38 == _match_key_bytes_1_T_1[6:0] ? phv_data_56 : _GEN_645; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_647 = 7'h39 == _match_key_bytes_1_T_1[6:0] ? phv_data_57 : _GEN_646; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_648 = 7'h3a == _match_key_bytes_1_T_1[6:0] ? phv_data_58 : _GEN_647; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_649 = 7'h3b == _match_key_bytes_1_T_1[6:0] ? phv_data_59 : _GEN_648; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_650 = 7'h3c == _match_key_bytes_1_T_1[6:0] ? phv_data_60 : _GEN_649; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_651 = 7'h3d == _match_key_bytes_1_T_1[6:0] ? phv_data_61 : _GEN_650; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_652 = 7'h3e == _match_key_bytes_1_T_1[6:0] ? phv_data_62 : _GEN_651; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_653 = 7'h3f == _match_key_bytes_1_T_1[6:0] ? phv_data_63 : _GEN_652; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_654 = 7'h40 == _match_key_bytes_1_T_1[6:0] ? phv_data_64 : _GEN_653; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_655 = 7'h41 == _match_key_bytes_1_T_1[6:0] ? phv_data_65 : _GEN_654; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_656 = 7'h42 == _match_key_bytes_1_T_1[6:0] ? phv_data_66 : _GEN_655; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_657 = 7'h43 == _match_key_bytes_1_T_1[6:0] ? phv_data_67 : _GEN_656; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_658 = 7'h44 == _match_key_bytes_1_T_1[6:0] ? phv_data_68 : _GEN_657; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_659 = 7'h45 == _match_key_bytes_1_T_1[6:0] ? phv_data_69 : _GEN_658; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_660 = 7'h46 == _match_key_bytes_1_T_1[6:0] ? phv_data_70 : _GEN_659; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_661 = 7'h47 == _match_key_bytes_1_T_1[6:0] ? phv_data_71 : _GEN_660; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_662 = 7'h48 == _match_key_bytes_1_T_1[6:0] ? phv_data_72 : _GEN_661; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_663 = 7'h49 == _match_key_bytes_1_T_1[6:0] ? phv_data_73 : _GEN_662; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_664 = 7'h4a == _match_key_bytes_1_T_1[6:0] ? phv_data_74 : _GEN_663; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_665 = 7'h4b == _match_key_bytes_1_T_1[6:0] ? phv_data_75 : _GEN_664; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_666 = 7'h4c == _match_key_bytes_1_T_1[6:0] ? phv_data_76 : _GEN_665; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_667 = 7'h4d == _match_key_bytes_1_T_1[6:0] ? phv_data_77 : _GEN_666; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_668 = 7'h4e == _match_key_bytes_1_T_1[6:0] ? phv_data_78 : _GEN_667; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_669 = 7'h4f == _match_key_bytes_1_T_1[6:0] ? phv_data_79 : _GEN_668; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_670 = 7'h50 == _match_key_bytes_1_T_1[6:0] ? phv_data_80 : _GEN_669; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_671 = 7'h51 == _match_key_bytes_1_T_1[6:0] ? phv_data_81 : _GEN_670; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_672 = 7'h52 == _match_key_bytes_1_T_1[6:0] ? phv_data_82 : _GEN_671; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_673 = 7'h53 == _match_key_bytes_1_T_1[6:0] ? phv_data_83 : _GEN_672; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_674 = 7'h54 == _match_key_bytes_1_T_1[6:0] ? phv_data_84 : _GEN_673; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_675 = 7'h55 == _match_key_bytes_1_T_1[6:0] ? phv_data_85 : _GEN_674; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_676 = 7'h56 == _match_key_bytes_1_T_1[6:0] ? phv_data_86 : _GEN_675; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_677 = 7'h57 == _match_key_bytes_1_T_1[6:0] ? phv_data_87 : _GEN_676; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_678 = 7'h58 == _match_key_bytes_1_T_1[6:0] ? phv_data_88 : _GEN_677; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_679 = 7'h59 == _match_key_bytes_1_T_1[6:0] ? phv_data_89 : _GEN_678; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_680 = 7'h5a == _match_key_bytes_1_T_1[6:0] ? phv_data_90 : _GEN_679; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_681 = 7'h5b == _match_key_bytes_1_T_1[6:0] ? phv_data_91 : _GEN_680; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_682 = 7'h5c == _match_key_bytes_1_T_1[6:0] ? phv_data_92 : _GEN_681; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_683 = 7'h5d == _match_key_bytes_1_T_1[6:0] ? phv_data_93 : _GEN_682; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_684 = 7'h5e == _match_key_bytes_1_T_1[6:0] ? phv_data_94 : _GEN_683; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_685 = 7'h5f == _match_key_bytes_1_T_1[6:0] ? phv_data_95 : _GEN_684; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_1 = 4'h6 < _GEN_6 ? _GEN_685 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_0_T_1 = key_offset + 8'h7; // @[matcher.scala 72:98]
  wire [7:0] _GEN_688 = 7'h1 == _match_key_bytes_0_T_1[6:0] ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_689 = 7'h2 == _match_key_bytes_0_T_1[6:0] ? phv_data_2 : _GEN_688; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_690 = 7'h3 == _match_key_bytes_0_T_1[6:0] ? phv_data_3 : _GEN_689; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_691 = 7'h4 == _match_key_bytes_0_T_1[6:0] ? phv_data_4 : _GEN_690; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_692 = 7'h5 == _match_key_bytes_0_T_1[6:0] ? phv_data_5 : _GEN_691; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_693 = 7'h6 == _match_key_bytes_0_T_1[6:0] ? phv_data_6 : _GEN_692; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_694 = 7'h7 == _match_key_bytes_0_T_1[6:0] ? phv_data_7 : _GEN_693; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_695 = 7'h8 == _match_key_bytes_0_T_1[6:0] ? phv_data_8 : _GEN_694; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_696 = 7'h9 == _match_key_bytes_0_T_1[6:0] ? phv_data_9 : _GEN_695; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_697 = 7'ha == _match_key_bytes_0_T_1[6:0] ? phv_data_10 : _GEN_696; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_698 = 7'hb == _match_key_bytes_0_T_1[6:0] ? phv_data_11 : _GEN_697; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_699 = 7'hc == _match_key_bytes_0_T_1[6:0] ? phv_data_12 : _GEN_698; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_700 = 7'hd == _match_key_bytes_0_T_1[6:0] ? phv_data_13 : _GEN_699; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_701 = 7'he == _match_key_bytes_0_T_1[6:0] ? phv_data_14 : _GEN_700; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_702 = 7'hf == _match_key_bytes_0_T_1[6:0] ? phv_data_15 : _GEN_701; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_703 = 7'h10 == _match_key_bytes_0_T_1[6:0] ? phv_data_16 : _GEN_702; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_704 = 7'h11 == _match_key_bytes_0_T_1[6:0] ? phv_data_17 : _GEN_703; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_705 = 7'h12 == _match_key_bytes_0_T_1[6:0] ? phv_data_18 : _GEN_704; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_706 = 7'h13 == _match_key_bytes_0_T_1[6:0] ? phv_data_19 : _GEN_705; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_707 = 7'h14 == _match_key_bytes_0_T_1[6:0] ? phv_data_20 : _GEN_706; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_708 = 7'h15 == _match_key_bytes_0_T_1[6:0] ? phv_data_21 : _GEN_707; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_709 = 7'h16 == _match_key_bytes_0_T_1[6:0] ? phv_data_22 : _GEN_708; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_710 = 7'h17 == _match_key_bytes_0_T_1[6:0] ? phv_data_23 : _GEN_709; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_711 = 7'h18 == _match_key_bytes_0_T_1[6:0] ? phv_data_24 : _GEN_710; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_712 = 7'h19 == _match_key_bytes_0_T_1[6:0] ? phv_data_25 : _GEN_711; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_713 = 7'h1a == _match_key_bytes_0_T_1[6:0] ? phv_data_26 : _GEN_712; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_714 = 7'h1b == _match_key_bytes_0_T_1[6:0] ? phv_data_27 : _GEN_713; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_715 = 7'h1c == _match_key_bytes_0_T_1[6:0] ? phv_data_28 : _GEN_714; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_716 = 7'h1d == _match_key_bytes_0_T_1[6:0] ? phv_data_29 : _GEN_715; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_717 = 7'h1e == _match_key_bytes_0_T_1[6:0] ? phv_data_30 : _GEN_716; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_718 = 7'h1f == _match_key_bytes_0_T_1[6:0] ? phv_data_31 : _GEN_717; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_719 = 7'h20 == _match_key_bytes_0_T_1[6:0] ? phv_data_32 : _GEN_718; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_720 = 7'h21 == _match_key_bytes_0_T_1[6:0] ? phv_data_33 : _GEN_719; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_721 = 7'h22 == _match_key_bytes_0_T_1[6:0] ? phv_data_34 : _GEN_720; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_722 = 7'h23 == _match_key_bytes_0_T_1[6:0] ? phv_data_35 : _GEN_721; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_723 = 7'h24 == _match_key_bytes_0_T_1[6:0] ? phv_data_36 : _GEN_722; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_724 = 7'h25 == _match_key_bytes_0_T_1[6:0] ? phv_data_37 : _GEN_723; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_725 = 7'h26 == _match_key_bytes_0_T_1[6:0] ? phv_data_38 : _GEN_724; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_726 = 7'h27 == _match_key_bytes_0_T_1[6:0] ? phv_data_39 : _GEN_725; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_727 = 7'h28 == _match_key_bytes_0_T_1[6:0] ? phv_data_40 : _GEN_726; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_728 = 7'h29 == _match_key_bytes_0_T_1[6:0] ? phv_data_41 : _GEN_727; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_729 = 7'h2a == _match_key_bytes_0_T_1[6:0] ? phv_data_42 : _GEN_728; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_730 = 7'h2b == _match_key_bytes_0_T_1[6:0] ? phv_data_43 : _GEN_729; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_731 = 7'h2c == _match_key_bytes_0_T_1[6:0] ? phv_data_44 : _GEN_730; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_732 = 7'h2d == _match_key_bytes_0_T_1[6:0] ? phv_data_45 : _GEN_731; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_733 = 7'h2e == _match_key_bytes_0_T_1[6:0] ? phv_data_46 : _GEN_732; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_734 = 7'h2f == _match_key_bytes_0_T_1[6:0] ? phv_data_47 : _GEN_733; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_735 = 7'h30 == _match_key_bytes_0_T_1[6:0] ? phv_data_48 : _GEN_734; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_736 = 7'h31 == _match_key_bytes_0_T_1[6:0] ? phv_data_49 : _GEN_735; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_737 = 7'h32 == _match_key_bytes_0_T_1[6:0] ? phv_data_50 : _GEN_736; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_738 = 7'h33 == _match_key_bytes_0_T_1[6:0] ? phv_data_51 : _GEN_737; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_739 = 7'h34 == _match_key_bytes_0_T_1[6:0] ? phv_data_52 : _GEN_738; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_740 = 7'h35 == _match_key_bytes_0_T_1[6:0] ? phv_data_53 : _GEN_739; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_741 = 7'h36 == _match_key_bytes_0_T_1[6:0] ? phv_data_54 : _GEN_740; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_742 = 7'h37 == _match_key_bytes_0_T_1[6:0] ? phv_data_55 : _GEN_741; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_743 = 7'h38 == _match_key_bytes_0_T_1[6:0] ? phv_data_56 : _GEN_742; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_744 = 7'h39 == _match_key_bytes_0_T_1[6:0] ? phv_data_57 : _GEN_743; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_745 = 7'h3a == _match_key_bytes_0_T_1[6:0] ? phv_data_58 : _GEN_744; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_746 = 7'h3b == _match_key_bytes_0_T_1[6:0] ? phv_data_59 : _GEN_745; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_747 = 7'h3c == _match_key_bytes_0_T_1[6:0] ? phv_data_60 : _GEN_746; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_748 = 7'h3d == _match_key_bytes_0_T_1[6:0] ? phv_data_61 : _GEN_747; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_749 = 7'h3e == _match_key_bytes_0_T_1[6:0] ? phv_data_62 : _GEN_748; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_750 = 7'h3f == _match_key_bytes_0_T_1[6:0] ? phv_data_63 : _GEN_749; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_751 = 7'h40 == _match_key_bytes_0_T_1[6:0] ? phv_data_64 : _GEN_750; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_752 = 7'h41 == _match_key_bytes_0_T_1[6:0] ? phv_data_65 : _GEN_751; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_753 = 7'h42 == _match_key_bytes_0_T_1[6:0] ? phv_data_66 : _GEN_752; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_754 = 7'h43 == _match_key_bytes_0_T_1[6:0] ? phv_data_67 : _GEN_753; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_755 = 7'h44 == _match_key_bytes_0_T_1[6:0] ? phv_data_68 : _GEN_754; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_756 = 7'h45 == _match_key_bytes_0_T_1[6:0] ? phv_data_69 : _GEN_755; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_757 = 7'h46 == _match_key_bytes_0_T_1[6:0] ? phv_data_70 : _GEN_756; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_758 = 7'h47 == _match_key_bytes_0_T_1[6:0] ? phv_data_71 : _GEN_757; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_759 = 7'h48 == _match_key_bytes_0_T_1[6:0] ? phv_data_72 : _GEN_758; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_760 = 7'h49 == _match_key_bytes_0_T_1[6:0] ? phv_data_73 : _GEN_759; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_761 = 7'h4a == _match_key_bytes_0_T_1[6:0] ? phv_data_74 : _GEN_760; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_762 = 7'h4b == _match_key_bytes_0_T_1[6:0] ? phv_data_75 : _GEN_761; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_763 = 7'h4c == _match_key_bytes_0_T_1[6:0] ? phv_data_76 : _GEN_762; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_764 = 7'h4d == _match_key_bytes_0_T_1[6:0] ? phv_data_77 : _GEN_763; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_765 = 7'h4e == _match_key_bytes_0_T_1[6:0] ? phv_data_78 : _GEN_764; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_766 = 7'h4f == _match_key_bytes_0_T_1[6:0] ? phv_data_79 : _GEN_765; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_767 = 7'h50 == _match_key_bytes_0_T_1[6:0] ? phv_data_80 : _GEN_766; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_768 = 7'h51 == _match_key_bytes_0_T_1[6:0] ? phv_data_81 : _GEN_767; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_769 = 7'h52 == _match_key_bytes_0_T_1[6:0] ? phv_data_82 : _GEN_768; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_770 = 7'h53 == _match_key_bytes_0_T_1[6:0] ? phv_data_83 : _GEN_769; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_771 = 7'h54 == _match_key_bytes_0_T_1[6:0] ? phv_data_84 : _GEN_770; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_772 = 7'h55 == _match_key_bytes_0_T_1[6:0] ? phv_data_85 : _GEN_771; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_773 = 7'h56 == _match_key_bytes_0_T_1[6:0] ? phv_data_86 : _GEN_772; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_774 = 7'h57 == _match_key_bytes_0_T_1[6:0] ? phv_data_87 : _GEN_773; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_775 = 7'h58 == _match_key_bytes_0_T_1[6:0] ? phv_data_88 : _GEN_774; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_776 = 7'h59 == _match_key_bytes_0_T_1[6:0] ? phv_data_89 : _GEN_775; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_777 = 7'h5a == _match_key_bytes_0_T_1[6:0] ? phv_data_90 : _GEN_776; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_778 = 7'h5b == _match_key_bytes_0_T_1[6:0] ? phv_data_91 : _GEN_777; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_779 = 7'h5c == _match_key_bytes_0_T_1[6:0] ? phv_data_92 : _GEN_778; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_780 = 7'h5d == _match_key_bytes_0_T_1[6:0] ? phv_data_93 : _GEN_779; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_781 = 7'h5e == _match_key_bytes_0_T_1[6:0] ? phv_data_94 : _GEN_780; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_782 = 7'h5f == _match_key_bytes_0_T_1[6:0] ? phv_data_95 : _GEN_781; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_0 = 4'h7 < _GEN_6 ? _GEN_782 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [63:0] match_key = {match_key_bytes_0,match_key_bytes_1,match_key_bytes_2,match_key_bytes_3,match_key_bytes_4,
    match_key_bytes_5,match_key_bytes_6,match_key_bytes_7}; // @[Cat.scala 30:58]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[matcher.scala 60:25]
  assign io_match_key = phv_is_valid_processor ? match_key : 64'h0; // @[matcher.scala 65:39 matcher.scala 79:26 matcher.scala 81:26]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[matcher.scala 59:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[matcher.scala 59:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[matcher.scala 59:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[matcher.scala 59:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[matcher.scala 59:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[matcher.scala 59:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[matcher.scala 59:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[matcher.scala 59:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[matcher.scala 59:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[matcher.scala 59:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[matcher.scala 59:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[matcher.scala 59:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[matcher.scala 59:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[matcher.scala 59:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[matcher.scala 59:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[matcher.scala 59:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[matcher.scala 59:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[matcher.scala 59:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[matcher.scala 59:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[matcher.scala 59:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[matcher.scala 59:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[matcher.scala 59:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[matcher.scala 59:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[matcher.scala 59:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[matcher.scala 59:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[matcher.scala 59:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[matcher.scala 59:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[matcher.scala 59:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[matcher.scala 59:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[matcher.scala 59:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[matcher.scala 59:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[matcher.scala 59:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[matcher.scala 59:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[matcher.scala 59:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[matcher.scala 59:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[matcher.scala 59:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[matcher.scala 59:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[matcher.scala 59:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[matcher.scala 59:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[matcher.scala 59:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[matcher.scala 59:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[matcher.scala 59:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[matcher.scala 59:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[matcher.scala 59:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[matcher.scala 59:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[matcher.scala 59:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[matcher.scala 59:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[matcher.scala 59:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[matcher.scala 59:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[matcher.scala 59:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[matcher.scala 59:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[matcher.scala 59:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[matcher.scala 59:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[matcher.scala 59:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[matcher.scala 59:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[matcher.scala 59:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[matcher.scala 59:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[matcher.scala 59:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[matcher.scala 59:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[matcher.scala 59:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[matcher.scala 59:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[matcher.scala 59:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[matcher.scala 59:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[matcher.scala 59:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[matcher.scala 59:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[matcher.scala 59:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[matcher.scala 59:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[matcher.scala 59:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[matcher.scala 59:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[matcher.scala 59:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[matcher.scala 59:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[matcher.scala 59:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[matcher.scala 59:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[matcher.scala 59:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[matcher.scala 59:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[matcher.scala 59:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[matcher.scala 59:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[matcher.scala 59:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[matcher.scala 59:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[matcher.scala 59:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[matcher.scala 59:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[matcher.scala 59:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[matcher.scala 59:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[matcher.scala 59:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[matcher.scala 59:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[matcher.scala 59:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[matcher.scala 59:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[matcher.scala 59:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[matcher.scala 59:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[matcher.scala 59:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[matcher.scala 59:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[matcher.scala 59:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[matcher.scala 59:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[matcher.scala 59:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[matcher.scala 59:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[matcher.scala 59:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[matcher.scala 59:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[matcher.scala 59:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[matcher.scala 59:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[matcher.scala 59:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[matcher.scala 59:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[matcher.scala 59:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[matcher.scala 59:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[matcher.scala 59:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[matcher.scala 59:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[matcher.scala 59:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[matcher.scala 59:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[matcher.scala 59:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[matcher.scala 59:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[matcher.scala 59:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[matcher.scala 59:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[matcher.scala 59:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[matcher.scala 59:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[matcher.scala 59:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[matcher.scala 59:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[matcher.scala 59:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[matcher.scala 59:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[matcher.scala 59:13]
    key_offset <= io_key_offset; // @[matcher.scala 63:20]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_header_0 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  phv_header_1 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  phv_header_2 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  phv_header_3 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  phv_header_4 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  phv_header_5 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  phv_header_6 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  phv_header_7 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  phv_header_8 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  phv_header_9 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  phv_header_10 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  phv_header_11 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  phv_header_12 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  phv_header_13 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  phv_header_14 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  phv_header_15 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  phv_next_config_id = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  key_offset = _RAND_118[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
