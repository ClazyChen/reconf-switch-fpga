module ExecutorPISA(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input         io_hit,
  input  [63:0] io_match_value,
  input         io_action_mod_en_0,
  input         io_action_mod_en_1,
  input  [7:0]  io_action_mod_addr,
  input  [63:0] io_action_mod_data_0,
  input  [63:0] io_action_mod_data_1
);
  wire  pipe1_clock; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_0; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_1; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_2; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_3; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_4; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_5; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_6; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_7; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_8; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_9; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_10; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_11; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_12; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_13; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_14; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_15; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_16; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_17; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_18; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_19; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_20; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_21; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_22; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_23; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_24; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_25; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_26; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_27; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_28; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_29; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_30; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_31; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_32; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_33; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_34; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_35; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_36; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_37; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_38; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_39; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_40; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_41; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_42; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_43; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_44; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_45; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_46; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_47; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_48; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_49; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_50; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_51; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_52; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_53; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_54; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_55; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_56; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_57; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_58; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_59; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_60; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_61; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_62; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_63; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_64; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_65; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_66; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_67; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_68; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_69; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_70; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_71; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_72; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_73; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_74; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_75; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_76; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_77; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_78; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_79; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_80; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_81; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_82; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_83; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_84; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_85; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_86; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_87; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_88; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_89; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_90; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_91; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_92; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_93; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_94; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_95; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_96; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_97; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_98; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_99; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_100; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_101; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_102; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_103; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_104; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_105; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_106; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_107; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_108; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_109; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_110; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_111; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_112; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_113; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_114; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_115; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_116; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_117; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_118; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_119; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_120; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_121; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_122; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_123; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_124; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_125; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_126; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_127; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_128; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_129; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_130; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_131; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_132; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_133; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_134; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_135; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_136; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_137; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_138; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_139; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_140; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_141; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_142; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_143; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_144; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_145; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_146; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_147; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_148; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_149; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_150; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_151; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_152; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_153; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_154; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_155; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_156; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_157; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_158; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_159; // @[executor_pisa.scala 286:23]
  wire  pipe1_io_pipe_phv_in_next_config_id; // @[executor_pisa.scala 286:23]
  wire  pipe1_io_pipe_phv_in_is_valid_processor; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_0; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_1; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_2; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_3; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_4; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_5; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_6; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_7; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_8; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_9; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_10; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_11; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_12; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_13; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_14; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_15; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_16; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_17; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_18; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_19; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_20; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_21; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_22; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_23; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_24; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_25; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_26; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_27; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_28; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_29; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_30; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_31; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_32; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_33; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_34; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_35; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_36; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_37; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_38; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_39; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_40; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_41; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_42; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_43; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_44; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_45; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_46; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_47; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_48; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_49; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_50; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_51; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_52; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_53; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_54; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_55; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_56; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_57; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_58; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_59; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_60; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_61; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_62; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_63; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_64; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_65; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_66; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_67; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_68; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_69; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_70; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_71; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_72; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_73; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_74; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_75; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_76; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_77; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_78; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_79; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_80; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_81; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_82; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_83; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_84; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_85; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_86; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_87; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_88; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_89; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_90; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_91; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_92; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_93; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_94; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_95; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_96; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_97; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_98; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_99; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_100; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_101; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_102; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_103; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_104; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_105; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_106; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_107; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_108; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_109; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_110; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_111; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_112; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_113; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_114; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_115; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_116; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_117; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_118; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_119; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_120; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_121; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_122; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_123; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_124; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_125; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_126; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_127; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_128; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_129; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_130; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_131; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_132; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_133; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_134; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_135; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_136; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_137; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_138; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_139; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_140; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_141; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_142; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_143; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_144; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_145; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_146; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_147; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_148; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_149; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_150; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_151; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_152; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_153; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_154; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_155; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_156; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_157; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_158; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_159; // @[executor_pisa.scala 286:23]
  wire  pipe1_io_pipe_phv_out_next_config_id; // @[executor_pisa.scala 286:23]
  wire  pipe1_io_pipe_phv_out_is_valid_processor; // @[executor_pisa.scala 286:23]
  wire  pipe1_io_hit; // @[executor_pisa.scala 286:23]
  wire [63:0] pipe1_io_match_value; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_args_out_0; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_args_out_1; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_args_out_2; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_args_out_3; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_args_out_4; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_args_out_5; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_args_out_6; // @[executor_pisa.scala 286:23]
  wire [31:0] pipe1_io_vliw_out_0; // @[executor_pisa.scala 286:23]
  wire [31:0] pipe1_io_vliw_out_1; // @[executor_pisa.scala 286:23]
  wire [31:0] pipe1_io_vliw_out_2; // @[executor_pisa.scala 286:23]
  wire [31:0] pipe1_io_vliw_out_3; // @[executor_pisa.scala 286:23]
  wire  pipe1_io_action_mod_en_0; // @[executor_pisa.scala 286:23]
  wire  pipe1_io_action_mod_en_1; // @[executor_pisa.scala 286:23]
  wire [7:0] pipe1_io_action_mod_addr; // @[executor_pisa.scala 286:23]
  wire [63:0] pipe1_io_action_mod_data_0; // @[executor_pisa.scala 286:23]
  wire [63:0] pipe1_io_action_mod_data_1; // @[executor_pisa.scala 286:23]
  wire  pipe2_clock; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_0; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_1; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_2; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_3; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_4; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_5; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_6; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_7; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_8; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_9; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_10; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_11; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_12; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_13; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_14; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_15; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_16; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_17; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_18; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_19; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_20; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_21; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_22; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_23; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_24; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_25; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_26; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_27; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_28; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_29; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_30; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_31; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_32; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_33; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_34; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_35; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_36; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_37; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_38; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_39; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_40; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_41; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_42; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_43; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_44; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_45; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_46; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_47; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_48; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_49; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_50; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_51; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_52; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_53; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_54; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_55; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_56; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_57; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_58; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_59; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_60; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_61; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_62; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_63; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_64; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_65; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_66; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_67; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_68; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_69; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_70; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_71; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_72; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_73; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_74; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_75; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_76; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_77; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_78; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_79; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_80; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_81; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_82; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_83; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_84; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_85; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_86; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_87; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_88; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_89; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_90; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_91; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_92; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_93; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_94; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_95; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_96; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_97; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_98; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_99; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_100; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_101; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_102; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_103; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_104; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_105; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_106; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_107; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_108; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_109; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_110; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_111; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_112; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_113; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_114; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_115; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_116; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_117; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_118; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_119; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_120; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_121; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_122; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_123; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_124; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_125; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_126; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_127; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_128; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_129; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_130; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_131; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_132; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_133; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_134; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_135; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_136; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_137; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_138; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_139; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_140; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_141; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_142; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_143; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_144; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_145; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_146; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_147; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_148; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_149; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_150; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_151; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_152; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_153; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_154; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_155; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_156; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_157; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_158; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_159; // @[executor_pisa.scala 287:23]
  wire  pipe2_io_pipe_phv_in_next_config_id; // @[executor_pisa.scala 287:23]
  wire  pipe2_io_pipe_phv_in_is_valid_processor; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_0; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_1; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_2; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_3; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_4; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_5; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_6; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_7; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_8; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_9; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_10; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_11; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_12; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_13; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_14; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_15; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_16; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_17; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_18; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_19; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_20; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_21; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_22; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_23; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_24; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_25; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_26; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_27; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_28; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_29; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_30; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_31; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_32; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_33; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_34; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_35; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_36; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_37; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_38; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_39; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_40; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_41; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_42; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_43; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_44; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_45; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_46; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_47; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_48; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_49; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_50; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_51; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_52; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_53; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_54; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_55; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_56; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_57; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_58; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_59; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_60; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_61; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_62; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_63; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_64; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_65; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_66; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_67; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_68; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_69; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_70; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_71; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_72; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_73; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_74; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_75; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_76; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_77; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_78; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_79; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_80; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_81; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_82; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_83; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_84; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_85; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_86; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_87; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_88; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_89; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_90; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_91; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_92; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_93; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_94; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_95; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_96; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_97; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_98; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_99; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_100; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_101; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_102; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_103; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_104; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_105; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_106; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_107; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_108; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_109; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_110; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_111; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_112; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_113; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_114; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_115; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_116; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_117; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_118; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_119; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_120; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_121; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_122; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_123; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_124; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_125; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_126; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_127; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_128; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_129; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_130; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_131; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_132; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_133; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_134; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_135; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_136; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_137; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_138; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_139; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_140; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_141; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_142; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_143; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_144; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_145; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_146; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_147; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_148; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_149; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_150; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_151; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_152; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_153; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_154; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_155; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_156; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_157; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_158; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_159; // @[executor_pisa.scala 287:23]
  wire  pipe2_io_pipe_phv_out_next_config_id; // @[executor_pisa.scala 287:23]
  wire  pipe2_io_pipe_phv_out_is_valid_processor; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_args_in_0; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_args_in_1; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_args_in_2; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_args_in_3; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_args_in_4; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_args_in_5; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_args_in_6; // @[executor_pisa.scala 287:23]
  wire [31:0] pipe2_io_vliw_in_0; // @[executor_pisa.scala 287:23]
  wire [31:0] pipe2_io_vliw_in_1; // @[executor_pisa.scala 287:23]
  wire [31:0] pipe2_io_vliw_in_2; // @[executor_pisa.scala 287:23]
  wire [31:0] pipe2_io_vliw_in_3; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_args_out_0; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_args_out_1; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_args_out_2; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_args_out_3; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_args_out_4; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_args_out_5; // @[executor_pisa.scala 287:23]
  wire [7:0] pipe2_io_args_out_6; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_0; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_1; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_2; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_3; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_4; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_5; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_6; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_7; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_8; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_9; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_10; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_11; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_12; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_13; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_14; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_15; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_16; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_17; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_18; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_19; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_20; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_21; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_22; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_23; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_24; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_25; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_26; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_27; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_28; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_29; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_30; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_31; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_32; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_33; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_34; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_35; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_36; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_37; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_38; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_39; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_40; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_41; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_42; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_43; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_44; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_45; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_46; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_47; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_48; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_49; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_50; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_51; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_52; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_53; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_54; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_55; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_56; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_57; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_58; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_59; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_60; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_61; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_62; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_63; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_64; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_65; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_66; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_67; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_68; // @[executor_pisa.scala 287:23]
  wire [17:0] pipe2_io_vliw_out_69; // @[executor_pisa.scala 287:23]
  wire [14:0] pipe2_io_nid_out; // @[executor_pisa.scala 287:23]
  wire  pipe3_clock; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_0; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_1; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_2; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_3; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_4; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_5; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_6; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_7; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_8; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_9; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_10; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_11; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_12; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_13; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_14; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_15; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_16; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_17; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_18; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_19; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_20; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_21; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_22; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_23; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_24; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_25; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_26; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_27; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_28; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_29; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_30; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_31; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_32; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_33; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_34; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_35; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_36; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_37; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_38; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_39; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_40; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_41; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_42; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_43; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_44; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_45; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_46; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_47; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_48; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_49; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_50; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_51; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_52; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_53; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_54; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_55; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_56; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_57; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_58; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_59; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_60; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_61; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_62; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_63; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_64; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_65; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_66; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_67; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_68; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_69; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_70; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_71; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_72; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_73; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_74; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_75; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_76; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_77; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_78; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_79; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_80; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_81; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_82; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_83; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_84; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_85; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_86; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_87; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_88; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_89; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_90; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_91; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_92; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_93; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_94; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_95; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_96; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_97; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_98; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_99; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_100; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_101; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_102; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_103; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_104; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_105; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_106; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_107; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_108; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_109; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_110; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_111; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_112; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_113; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_114; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_115; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_116; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_117; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_118; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_119; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_120; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_121; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_122; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_123; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_124; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_125; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_126; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_127; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_128; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_129; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_130; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_131; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_132; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_133; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_134; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_135; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_136; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_137; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_138; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_139; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_140; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_141; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_142; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_143; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_144; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_145; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_146; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_147; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_148; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_149; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_150; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_151; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_152; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_153; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_154; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_155; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_156; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_157; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_158; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_159; // @[executor_pisa.scala 288:23]
  wire  pipe3_io_pipe_phv_in_next_config_id; // @[executor_pisa.scala 288:23]
  wire  pipe3_io_pipe_phv_in_is_valid_processor; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_0; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_1; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_2; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_3; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_4; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_5; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_6; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_7; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_8; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_9; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_10; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_11; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_12; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_13; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_14; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_15; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_16; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_17; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_18; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_19; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_20; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_21; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_22; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_23; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_24; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_25; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_26; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_27; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_28; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_29; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_30; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_31; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_32; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_33; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_34; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_35; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_36; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_37; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_38; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_39; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_40; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_41; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_42; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_43; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_44; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_45; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_46; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_47; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_48; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_49; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_50; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_51; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_52; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_53; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_54; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_55; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_56; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_57; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_58; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_59; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_60; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_61; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_62; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_63; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_64; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_65; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_66; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_67; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_68; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_69; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_70; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_71; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_72; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_73; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_74; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_75; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_76; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_77; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_78; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_79; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_80; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_81; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_82; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_83; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_84; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_85; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_86; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_87; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_88; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_89; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_90; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_91; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_92; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_93; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_94; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_95; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_96; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_97; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_98; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_99; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_100; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_101; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_102; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_103; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_104; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_105; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_106; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_107; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_108; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_109; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_110; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_111; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_112; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_113; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_114; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_115; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_116; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_117; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_118; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_119; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_120; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_121; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_122; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_123; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_124; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_125; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_126; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_127; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_128; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_129; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_130; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_131; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_132; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_133; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_134; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_135; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_136; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_137; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_138; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_139; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_140; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_141; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_142; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_143; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_144; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_145; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_146; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_147; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_148; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_149; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_150; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_151; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_152; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_153; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_154; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_155; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_156; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_157; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_158; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_159; // @[executor_pisa.scala 288:23]
  wire  pipe3_io_pipe_phv_out_next_config_id; // @[executor_pisa.scala 288:23]
  wire  pipe3_io_pipe_phv_out_is_valid_processor; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_args_in_0; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_args_in_1; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_args_in_2; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_args_in_3; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_args_in_4; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_args_in_5; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_args_in_6; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_0; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_1; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_2; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_3; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_4; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_5; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_6; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_7; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_8; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_9; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_10; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_11; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_12; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_13; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_14; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_15; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_16; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_17; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_18; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_19; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_20; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_21; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_22; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_23; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_24; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_25; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_26; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_27; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_28; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_29; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_30; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_31; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_32; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_33; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_34; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_35; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_36; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_37; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_38; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_39; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_40; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_41; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_42; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_43; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_44; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_45; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_46; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_47; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_48; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_49; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_50; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_51; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_52; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_53; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_54; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_55; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_56; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_57; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_58; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_59; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_60; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_61; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_62; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_63; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_64; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_65; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_66; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_67; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_68; // @[executor_pisa.scala 288:23]
  wire [17:0] pipe3_io_vliw_in_69; // @[executor_pisa.scala 288:23]
  wire [14:0] pipe3_io_nid_in; // @[executor_pisa.scala 288:23]
  wire [14:0] pipe3_io_nid_out; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_0; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_1; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_2; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_3; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_4; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_5; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_6; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_7; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_8; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_9; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_10; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_11; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_12; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_13; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_14; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_15; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_16; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_17; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_18; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_19; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_20; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_21; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_22; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_23; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_24; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_25; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_26; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_27; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_28; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_29; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_30; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_31; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_32; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_33; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_34; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_35; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_36; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_37; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_38; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_39; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_40; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_41; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_42; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_43; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_44; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_45; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_46; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_47; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_48; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_49; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_50; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_51; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_52; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_53; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_54; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_55; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_56; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_57; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_58; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_59; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_60; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_61; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_62; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_63; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_64; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_65; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_66; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_67; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_68; // @[executor_pisa.scala 288:23]
  wire [1:0] pipe3_io_tag_out_69; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_field_set_field8_0; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_field_set_field8_1; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_field_set_field8_2; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_field_set_field8_3; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_field_set_field8_4; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_field_set_field8_5; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_field_set_field8_6; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_field_set_field8_7; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_field_set_field8_8; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_field_set_field8_9; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_field_set_field8_10; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_field_set_field8_11; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_field_set_field8_12; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_field_set_field8_13; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_field_set_field8_14; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_field_set_field8_15; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_field_set_field8_16; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_field_set_field8_17; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_field_set_field8_18; // @[executor_pisa.scala 288:23]
  wire [7:0] pipe3_io_field_set_field8_19; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_0; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_1; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_2; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_3; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_4; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_5; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_6; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_7; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_8; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_9; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_10; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_11; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_12; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_13; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_14; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_15; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_16; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_17; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_18; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_19; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_20; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_21; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_22; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_23; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_24; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_25; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_26; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_27; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_28; // @[executor_pisa.scala 288:23]
  wire [15:0] pipe3_io_field_set_field16_29; // @[executor_pisa.scala 288:23]
  wire [31:0] pipe3_io_field_set_field32_0; // @[executor_pisa.scala 288:23]
  wire [31:0] pipe3_io_field_set_field32_1; // @[executor_pisa.scala 288:23]
  wire [31:0] pipe3_io_field_set_field32_2; // @[executor_pisa.scala 288:23]
  wire [31:0] pipe3_io_field_set_field32_3; // @[executor_pisa.scala 288:23]
  wire [31:0] pipe3_io_field_set_field32_4; // @[executor_pisa.scala 288:23]
  wire [31:0] pipe3_io_field_set_field32_5; // @[executor_pisa.scala 288:23]
  wire [31:0] pipe3_io_field_set_field32_6; // @[executor_pisa.scala 288:23]
  wire [31:0] pipe3_io_field_set_field32_7; // @[executor_pisa.scala 288:23]
  wire [31:0] pipe3_io_field_set_field32_8; // @[executor_pisa.scala 288:23]
  wire [31:0] pipe3_io_field_set_field32_9; // @[executor_pisa.scala 288:23]
  wire [31:0] pipe3_io_field_set_field32_10; // @[executor_pisa.scala 288:23]
  wire [31:0] pipe3_io_field_set_field32_11; // @[executor_pisa.scala 288:23]
  wire [31:0] pipe3_io_field_set_field32_12; // @[executor_pisa.scala 288:23]
  wire [31:0] pipe3_io_field_set_field32_13; // @[executor_pisa.scala 288:23]
  wire [31:0] pipe3_io_field_set_field32_14; // @[executor_pisa.scala 288:23]
  wire [31:0] pipe3_io_field_set_field32_15; // @[executor_pisa.scala 288:23]
  wire [31:0] pipe3_io_field_set_field32_16; // @[executor_pisa.scala 288:23]
  wire [31:0] pipe3_io_field_set_field32_17; // @[executor_pisa.scala 288:23]
  wire [31:0] pipe3_io_field_set_field32_18; // @[executor_pisa.scala 288:23]
  wire [31:0] pipe3_io_field_set_field32_19; // @[executor_pisa.scala 288:23]
  wire  pipe4_clock; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_0; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_1; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_2; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_3; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_4; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_5; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_6; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_7; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_8; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_9; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_10; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_11; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_12; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_13; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_14; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_15; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_16; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_17; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_18; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_19; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_20; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_21; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_22; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_23; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_24; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_25; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_26; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_27; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_28; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_29; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_30; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_31; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_32; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_33; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_34; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_35; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_36; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_37; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_38; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_39; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_40; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_41; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_42; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_43; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_44; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_45; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_46; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_47; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_48; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_49; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_50; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_51; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_52; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_53; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_54; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_55; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_56; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_57; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_58; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_59; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_60; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_61; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_62; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_63; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_64; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_65; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_66; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_67; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_68; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_69; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_70; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_71; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_72; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_73; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_74; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_75; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_76; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_77; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_78; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_79; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_80; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_81; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_82; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_83; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_84; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_85; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_86; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_87; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_88; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_89; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_90; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_91; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_92; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_93; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_94; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_95; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_96; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_97; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_98; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_99; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_100; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_101; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_102; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_103; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_104; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_105; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_106; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_107; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_108; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_109; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_110; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_111; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_112; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_113; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_114; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_115; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_116; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_117; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_118; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_119; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_120; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_121; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_122; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_123; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_124; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_125; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_126; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_127; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_128; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_129; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_130; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_131; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_132; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_133; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_134; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_135; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_136; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_137; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_138; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_139; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_140; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_141; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_142; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_143; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_144; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_145; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_146; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_147; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_148; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_149; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_150; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_151; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_152; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_153; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_154; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_155; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_156; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_157; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_158; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_159; // @[executor_pisa.scala 289:23]
  wire  pipe4_io_pipe_phv_in_next_config_id; // @[executor_pisa.scala 289:23]
  wire  pipe4_io_pipe_phv_in_is_valid_processor; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_0; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_1; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_2; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_3; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_4; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_5; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_6; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_7; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_8; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_9; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_10; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_11; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_12; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_13; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_14; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_15; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_16; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_17; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_18; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_19; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_20; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_21; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_22; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_23; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_24; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_25; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_26; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_27; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_28; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_29; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_30; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_31; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_32; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_33; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_34; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_35; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_36; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_37; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_38; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_39; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_40; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_41; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_42; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_43; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_44; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_45; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_46; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_47; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_48; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_49; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_50; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_51; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_52; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_53; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_54; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_55; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_56; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_57; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_58; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_59; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_60; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_61; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_62; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_63; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_64; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_65; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_66; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_67; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_68; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_69; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_70; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_71; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_72; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_73; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_74; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_75; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_76; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_77; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_78; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_79; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_80; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_81; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_82; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_83; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_84; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_85; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_86; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_87; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_88; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_89; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_90; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_91; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_92; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_93; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_94; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_95; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_96; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_97; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_98; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_99; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_100; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_101; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_102; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_103; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_104; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_105; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_106; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_107; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_108; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_109; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_110; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_111; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_112; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_113; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_114; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_115; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_116; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_117; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_118; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_119; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_120; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_121; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_122; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_123; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_124; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_125; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_126; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_127; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_128; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_129; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_130; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_131; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_132; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_133; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_134; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_135; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_136; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_137; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_138; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_139; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_140; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_141; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_142; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_143; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_144; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_145; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_146; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_147; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_148; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_149; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_150; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_151; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_152; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_153; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_154; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_155; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_156; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_157; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_158; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_159; // @[executor_pisa.scala 289:23]
  wire  pipe4_io_pipe_phv_out_next_config_id; // @[executor_pisa.scala 289:23]
  wire  pipe4_io_pipe_phv_out_is_valid_processor; // @[executor_pisa.scala 289:23]
  wire [14:0] pipe4_io_nid_in; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_0; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_1; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_2; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_3; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_4; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_5; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_6; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_7; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_8; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_9; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_10; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_11; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_12; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_13; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_14; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_15; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_16; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_17; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_18; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_19; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_20; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_21; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_22; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_23; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_24; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_25; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_26; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_27; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_28; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_29; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_30; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_31; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_32; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_33; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_34; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_35; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_36; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_37; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_38; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_39; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_40; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_41; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_42; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_43; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_44; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_45; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_46; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_47; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_48; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_49; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_50; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_51; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_52; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_53; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_54; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_55; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_56; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_57; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_58; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_59; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_60; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_61; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_62; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_63; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_64; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_65; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_66; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_67; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_68; // @[executor_pisa.scala 289:23]
  wire [1:0] pipe4_io_tag_in_69; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_field_set_field8_0; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_field_set_field8_1; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_field_set_field8_2; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_field_set_field8_3; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_field_set_field8_4; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_field_set_field8_5; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_field_set_field8_6; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_field_set_field8_7; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_field_set_field8_8; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_field_set_field8_9; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_field_set_field8_10; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_field_set_field8_11; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_field_set_field8_12; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_field_set_field8_13; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_field_set_field8_14; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_field_set_field8_15; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_field_set_field8_16; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_field_set_field8_17; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_field_set_field8_18; // @[executor_pisa.scala 289:23]
  wire [7:0] pipe4_io_field_set_field8_19; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_0; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_1; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_2; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_3; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_4; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_5; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_6; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_7; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_8; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_9; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_10; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_11; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_12; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_13; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_14; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_15; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_16; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_17; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_18; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_19; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_20; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_21; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_22; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_23; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_24; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_25; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_26; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_27; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_28; // @[executor_pisa.scala 289:23]
  wire [15:0] pipe4_io_field_set_field16_29; // @[executor_pisa.scala 289:23]
  wire [31:0] pipe4_io_field_set_field32_0; // @[executor_pisa.scala 289:23]
  wire [31:0] pipe4_io_field_set_field32_1; // @[executor_pisa.scala 289:23]
  wire [31:0] pipe4_io_field_set_field32_2; // @[executor_pisa.scala 289:23]
  wire [31:0] pipe4_io_field_set_field32_3; // @[executor_pisa.scala 289:23]
  wire [31:0] pipe4_io_field_set_field32_4; // @[executor_pisa.scala 289:23]
  wire [31:0] pipe4_io_field_set_field32_5; // @[executor_pisa.scala 289:23]
  wire [31:0] pipe4_io_field_set_field32_6; // @[executor_pisa.scala 289:23]
  wire [31:0] pipe4_io_field_set_field32_7; // @[executor_pisa.scala 289:23]
  wire [31:0] pipe4_io_field_set_field32_8; // @[executor_pisa.scala 289:23]
  wire [31:0] pipe4_io_field_set_field32_9; // @[executor_pisa.scala 289:23]
  wire [31:0] pipe4_io_field_set_field32_10; // @[executor_pisa.scala 289:23]
  wire [31:0] pipe4_io_field_set_field32_11; // @[executor_pisa.scala 289:23]
  wire [31:0] pipe4_io_field_set_field32_12; // @[executor_pisa.scala 289:23]
  wire [31:0] pipe4_io_field_set_field32_13; // @[executor_pisa.scala 289:23]
  wire [31:0] pipe4_io_field_set_field32_14; // @[executor_pisa.scala 289:23]
  wire [31:0] pipe4_io_field_set_field32_15; // @[executor_pisa.scala 289:23]
  wire [31:0] pipe4_io_field_set_field32_16; // @[executor_pisa.scala 289:23]
  wire [31:0] pipe4_io_field_set_field32_17; // @[executor_pisa.scala 289:23]
  wire [31:0] pipe4_io_field_set_field32_18; // @[executor_pisa.scala 289:23]
  wire [31:0] pipe4_io_field_set_field32_19; // @[executor_pisa.scala 289:23]
  ActionReaderPISA pipe1 ( // @[executor_pisa.scala 286:23]
    .clock(pipe1_clock),
    .io_pipe_phv_in_data_0(pipe1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe1_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe1_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe1_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe1_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe1_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe1_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe1_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe1_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe1_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe1_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe1_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe1_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe1_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe1_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe1_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe1_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe1_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe1_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe1_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe1_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe1_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe1_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe1_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe1_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe1_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe1_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe1_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe1_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe1_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe1_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe1_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe1_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe1_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe1_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe1_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe1_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe1_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe1_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe1_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe1_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe1_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe1_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe1_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe1_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe1_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe1_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe1_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe1_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe1_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe1_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe1_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe1_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe1_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe1_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe1_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe1_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe1_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe1_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe1_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe1_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe1_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe1_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe1_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe1_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_next_config_id(pipe1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe1_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe1_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe1_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe1_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe1_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe1_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe1_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe1_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe1_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe1_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe1_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe1_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe1_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe1_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe1_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe1_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe1_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe1_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe1_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe1_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe1_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe1_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe1_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe1_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe1_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe1_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe1_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe1_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe1_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe1_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe1_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe1_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe1_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe1_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe1_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe1_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe1_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe1_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe1_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe1_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe1_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe1_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe1_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe1_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe1_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe1_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe1_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe1_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe1_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe1_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe1_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe1_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe1_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe1_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe1_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe1_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe1_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe1_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe1_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe1_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe1_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe1_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe1_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe1_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe1_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_next_config_id(pipe1_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe1_io_pipe_phv_out_is_valid_processor),
    .io_hit(pipe1_io_hit),
    .io_match_value(pipe1_io_match_value),
    .io_args_out_0(pipe1_io_args_out_0),
    .io_args_out_1(pipe1_io_args_out_1),
    .io_args_out_2(pipe1_io_args_out_2),
    .io_args_out_3(pipe1_io_args_out_3),
    .io_args_out_4(pipe1_io_args_out_4),
    .io_args_out_5(pipe1_io_args_out_5),
    .io_args_out_6(pipe1_io_args_out_6),
    .io_vliw_out_0(pipe1_io_vliw_out_0),
    .io_vliw_out_1(pipe1_io_vliw_out_1),
    .io_vliw_out_2(pipe1_io_vliw_out_2),
    .io_vliw_out_3(pipe1_io_vliw_out_3),
    .io_action_mod_en_0(pipe1_io_action_mod_en_0),
    .io_action_mod_en_1(pipe1_io_action_mod_en_1),
    .io_action_mod_addr(pipe1_io_action_mod_addr),
    .io_action_mod_data_0(pipe1_io_action_mod_data_0),
    .io_action_mod_data_1(pipe1_io_action_mod_data_1)
  );
  PrimitiveDistributionPISA pipe2 ( // @[executor_pisa.scala 287:23]
    .clock(pipe2_clock),
    .io_pipe_phv_in_data_0(pipe2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe2_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe2_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe2_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe2_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe2_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe2_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe2_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe2_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe2_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe2_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe2_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe2_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe2_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe2_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe2_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe2_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe2_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe2_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe2_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe2_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe2_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe2_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe2_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe2_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe2_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe2_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe2_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe2_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe2_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe2_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe2_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe2_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe2_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe2_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe2_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe2_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe2_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe2_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe2_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe2_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe2_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe2_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe2_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe2_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe2_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe2_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe2_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe2_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe2_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe2_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe2_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe2_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe2_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe2_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe2_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe2_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe2_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe2_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe2_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe2_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe2_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe2_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe2_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe2_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_next_config_id(pipe2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe2_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe2_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe2_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe2_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe2_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe2_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe2_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe2_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe2_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe2_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe2_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe2_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe2_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe2_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe2_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe2_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe2_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe2_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe2_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe2_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe2_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe2_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe2_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe2_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe2_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe2_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe2_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe2_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe2_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe2_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe2_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe2_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe2_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe2_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe2_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe2_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe2_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe2_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe2_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe2_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe2_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe2_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe2_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe2_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe2_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe2_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe2_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe2_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe2_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe2_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe2_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe2_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe2_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe2_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe2_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe2_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe2_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe2_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe2_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe2_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe2_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe2_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe2_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe2_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe2_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_next_config_id(pipe2_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe2_io_pipe_phv_out_is_valid_processor),
    .io_args_in_0(pipe2_io_args_in_0),
    .io_args_in_1(pipe2_io_args_in_1),
    .io_args_in_2(pipe2_io_args_in_2),
    .io_args_in_3(pipe2_io_args_in_3),
    .io_args_in_4(pipe2_io_args_in_4),
    .io_args_in_5(pipe2_io_args_in_5),
    .io_args_in_6(pipe2_io_args_in_6),
    .io_vliw_in_0(pipe2_io_vliw_in_0),
    .io_vliw_in_1(pipe2_io_vliw_in_1),
    .io_vliw_in_2(pipe2_io_vliw_in_2),
    .io_vliw_in_3(pipe2_io_vliw_in_3),
    .io_args_out_0(pipe2_io_args_out_0),
    .io_args_out_1(pipe2_io_args_out_1),
    .io_args_out_2(pipe2_io_args_out_2),
    .io_args_out_3(pipe2_io_args_out_3),
    .io_args_out_4(pipe2_io_args_out_4),
    .io_args_out_5(pipe2_io_args_out_5),
    .io_args_out_6(pipe2_io_args_out_6),
    .io_vliw_out_0(pipe2_io_vliw_out_0),
    .io_vliw_out_1(pipe2_io_vliw_out_1),
    .io_vliw_out_2(pipe2_io_vliw_out_2),
    .io_vliw_out_3(pipe2_io_vliw_out_3),
    .io_vliw_out_4(pipe2_io_vliw_out_4),
    .io_vliw_out_5(pipe2_io_vliw_out_5),
    .io_vliw_out_6(pipe2_io_vliw_out_6),
    .io_vliw_out_7(pipe2_io_vliw_out_7),
    .io_vliw_out_8(pipe2_io_vliw_out_8),
    .io_vliw_out_9(pipe2_io_vliw_out_9),
    .io_vliw_out_10(pipe2_io_vliw_out_10),
    .io_vliw_out_11(pipe2_io_vliw_out_11),
    .io_vliw_out_12(pipe2_io_vliw_out_12),
    .io_vliw_out_13(pipe2_io_vliw_out_13),
    .io_vliw_out_14(pipe2_io_vliw_out_14),
    .io_vliw_out_15(pipe2_io_vliw_out_15),
    .io_vliw_out_16(pipe2_io_vliw_out_16),
    .io_vliw_out_17(pipe2_io_vliw_out_17),
    .io_vliw_out_18(pipe2_io_vliw_out_18),
    .io_vliw_out_19(pipe2_io_vliw_out_19),
    .io_vliw_out_20(pipe2_io_vliw_out_20),
    .io_vliw_out_21(pipe2_io_vliw_out_21),
    .io_vliw_out_22(pipe2_io_vliw_out_22),
    .io_vliw_out_23(pipe2_io_vliw_out_23),
    .io_vliw_out_24(pipe2_io_vliw_out_24),
    .io_vliw_out_25(pipe2_io_vliw_out_25),
    .io_vliw_out_26(pipe2_io_vliw_out_26),
    .io_vliw_out_27(pipe2_io_vliw_out_27),
    .io_vliw_out_28(pipe2_io_vliw_out_28),
    .io_vliw_out_29(pipe2_io_vliw_out_29),
    .io_vliw_out_30(pipe2_io_vliw_out_30),
    .io_vliw_out_31(pipe2_io_vliw_out_31),
    .io_vliw_out_32(pipe2_io_vliw_out_32),
    .io_vliw_out_33(pipe2_io_vliw_out_33),
    .io_vliw_out_34(pipe2_io_vliw_out_34),
    .io_vliw_out_35(pipe2_io_vliw_out_35),
    .io_vliw_out_36(pipe2_io_vliw_out_36),
    .io_vliw_out_37(pipe2_io_vliw_out_37),
    .io_vliw_out_38(pipe2_io_vliw_out_38),
    .io_vliw_out_39(pipe2_io_vliw_out_39),
    .io_vliw_out_40(pipe2_io_vliw_out_40),
    .io_vliw_out_41(pipe2_io_vliw_out_41),
    .io_vliw_out_42(pipe2_io_vliw_out_42),
    .io_vliw_out_43(pipe2_io_vliw_out_43),
    .io_vliw_out_44(pipe2_io_vliw_out_44),
    .io_vliw_out_45(pipe2_io_vliw_out_45),
    .io_vliw_out_46(pipe2_io_vliw_out_46),
    .io_vliw_out_47(pipe2_io_vliw_out_47),
    .io_vliw_out_48(pipe2_io_vliw_out_48),
    .io_vliw_out_49(pipe2_io_vliw_out_49),
    .io_vliw_out_50(pipe2_io_vliw_out_50),
    .io_vliw_out_51(pipe2_io_vliw_out_51),
    .io_vliw_out_52(pipe2_io_vliw_out_52),
    .io_vliw_out_53(pipe2_io_vliw_out_53),
    .io_vliw_out_54(pipe2_io_vliw_out_54),
    .io_vliw_out_55(pipe2_io_vliw_out_55),
    .io_vliw_out_56(pipe2_io_vliw_out_56),
    .io_vliw_out_57(pipe2_io_vliw_out_57),
    .io_vliw_out_58(pipe2_io_vliw_out_58),
    .io_vliw_out_59(pipe2_io_vliw_out_59),
    .io_vliw_out_60(pipe2_io_vliw_out_60),
    .io_vliw_out_61(pipe2_io_vliw_out_61),
    .io_vliw_out_62(pipe2_io_vliw_out_62),
    .io_vliw_out_63(pipe2_io_vliw_out_63),
    .io_vliw_out_64(pipe2_io_vliw_out_64),
    .io_vliw_out_65(pipe2_io_vliw_out_65),
    .io_vliw_out_66(pipe2_io_vliw_out_66),
    .io_vliw_out_67(pipe2_io_vliw_out_67),
    .io_vliw_out_68(pipe2_io_vliw_out_68),
    .io_vliw_out_69(pipe2_io_vliw_out_69),
    .io_nid_out(pipe2_io_nid_out)
  );
  PrimitiveGetSourcePISA pipe3 ( // @[executor_pisa.scala 288:23]
    .clock(pipe3_clock),
    .io_pipe_phv_in_data_0(pipe3_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe3_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe3_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe3_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe3_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe3_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe3_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe3_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe3_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe3_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe3_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe3_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe3_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe3_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe3_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe3_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe3_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe3_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe3_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe3_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe3_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe3_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe3_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe3_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe3_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe3_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe3_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe3_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe3_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe3_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe3_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe3_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe3_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe3_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe3_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe3_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe3_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe3_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe3_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe3_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe3_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe3_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe3_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe3_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe3_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe3_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe3_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe3_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe3_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe3_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe3_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe3_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe3_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe3_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe3_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe3_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe3_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe3_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe3_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe3_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe3_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe3_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe3_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe3_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe3_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe3_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe3_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe3_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe3_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe3_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe3_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe3_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe3_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe3_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe3_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe3_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe3_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe3_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe3_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe3_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe3_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe3_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe3_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe3_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe3_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe3_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe3_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe3_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe3_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe3_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe3_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe3_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe3_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe3_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe3_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe3_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe3_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe3_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe3_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe3_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe3_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe3_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe3_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe3_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe3_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe3_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe3_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe3_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe3_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe3_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe3_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe3_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe3_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe3_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe3_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe3_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe3_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe3_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe3_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe3_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe3_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe3_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe3_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe3_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe3_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe3_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe3_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe3_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe3_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe3_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe3_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe3_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe3_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe3_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe3_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe3_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe3_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe3_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe3_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe3_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe3_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe3_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe3_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe3_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe3_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe3_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe3_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe3_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe3_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe3_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe3_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe3_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe3_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe3_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe3_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe3_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe3_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe3_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe3_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe3_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_next_config_id(pipe3_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe3_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe3_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe3_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe3_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe3_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe3_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe3_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe3_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe3_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe3_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe3_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe3_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe3_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe3_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe3_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe3_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe3_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe3_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe3_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe3_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe3_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe3_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe3_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe3_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe3_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe3_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe3_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe3_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe3_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe3_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe3_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe3_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe3_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe3_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe3_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe3_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe3_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe3_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe3_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe3_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe3_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe3_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe3_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe3_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe3_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe3_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe3_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe3_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe3_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe3_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe3_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe3_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe3_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe3_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe3_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe3_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe3_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe3_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe3_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe3_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe3_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe3_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe3_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe3_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe3_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe3_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe3_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe3_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe3_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe3_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe3_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe3_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe3_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe3_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe3_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe3_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe3_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe3_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe3_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe3_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe3_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe3_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe3_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe3_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe3_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe3_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe3_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe3_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe3_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe3_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe3_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe3_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe3_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe3_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe3_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe3_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe3_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe3_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe3_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe3_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe3_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe3_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe3_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe3_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe3_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe3_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe3_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe3_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe3_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe3_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe3_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe3_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe3_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe3_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe3_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe3_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe3_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe3_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe3_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe3_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe3_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe3_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe3_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe3_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe3_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe3_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe3_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe3_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe3_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe3_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe3_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe3_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe3_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe3_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe3_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe3_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe3_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe3_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe3_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe3_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe3_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe3_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe3_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe3_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe3_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe3_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe3_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe3_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe3_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe3_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe3_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe3_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe3_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe3_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe3_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe3_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe3_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe3_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe3_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe3_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe3_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_next_config_id(pipe3_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe3_io_pipe_phv_out_is_valid_processor),
    .io_args_in_0(pipe3_io_args_in_0),
    .io_args_in_1(pipe3_io_args_in_1),
    .io_args_in_2(pipe3_io_args_in_2),
    .io_args_in_3(pipe3_io_args_in_3),
    .io_args_in_4(pipe3_io_args_in_4),
    .io_args_in_5(pipe3_io_args_in_5),
    .io_args_in_6(pipe3_io_args_in_6),
    .io_vliw_in_0(pipe3_io_vliw_in_0),
    .io_vliw_in_1(pipe3_io_vliw_in_1),
    .io_vliw_in_2(pipe3_io_vliw_in_2),
    .io_vliw_in_3(pipe3_io_vliw_in_3),
    .io_vliw_in_4(pipe3_io_vliw_in_4),
    .io_vliw_in_5(pipe3_io_vliw_in_5),
    .io_vliw_in_6(pipe3_io_vliw_in_6),
    .io_vliw_in_7(pipe3_io_vliw_in_7),
    .io_vliw_in_8(pipe3_io_vliw_in_8),
    .io_vliw_in_9(pipe3_io_vliw_in_9),
    .io_vliw_in_10(pipe3_io_vliw_in_10),
    .io_vliw_in_11(pipe3_io_vliw_in_11),
    .io_vliw_in_12(pipe3_io_vliw_in_12),
    .io_vliw_in_13(pipe3_io_vliw_in_13),
    .io_vliw_in_14(pipe3_io_vliw_in_14),
    .io_vliw_in_15(pipe3_io_vliw_in_15),
    .io_vliw_in_16(pipe3_io_vliw_in_16),
    .io_vliw_in_17(pipe3_io_vliw_in_17),
    .io_vliw_in_18(pipe3_io_vliw_in_18),
    .io_vliw_in_19(pipe3_io_vliw_in_19),
    .io_vliw_in_20(pipe3_io_vliw_in_20),
    .io_vliw_in_21(pipe3_io_vliw_in_21),
    .io_vliw_in_22(pipe3_io_vliw_in_22),
    .io_vliw_in_23(pipe3_io_vliw_in_23),
    .io_vliw_in_24(pipe3_io_vliw_in_24),
    .io_vliw_in_25(pipe3_io_vliw_in_25),
    .io_vliw_in_26(pipe3_io_vliw_in_26),
    .io_vliw_in_27(pipe3_io_vliw_in_27),
    .io_vliw_in_28(pipe3_io_vliw_in_28),
    .io_vliw_in_29(pipe3_io_vliw_in_29),
    .io_vliw_in_30(pipe3_io_vliw_in_30),
    .io_vliw_in_31(pipe3_io_vliw_in_31),
    .io_vliw_in_32(pipe3_io_vliw_in_32),
    .io_vliw_in_33(pipe3_io_vliw_in_33),
    .io_vliw_in_34(pipe3_io_vliw_in_34),
    .io_vliw_in_35(pipe3_io_vliw_in_35),
    .io_vliw_in_36(pipe3_io_vliw_in_36),
    .io_vliw_in_37(pipe3_io_vliw_in_37),
    .io_vliw_in_38(pipe3_io_vliw_in_38),
    .io_vliw_in_39(pipe3_io_vliw_in_39),
    .io_vliw_in_40(pipe3_io_vliw_in_40),
    .io_vliw_in_41(pipe3_io_vliw_in_41),
    .io_vliw_in_42(pipe3_io_vliw_in_42),
    .io_vliw_in_43(pipe3_io_vliw_in_43),
    .io_vliw_in_44(pipe3_io_vliw_in_44),
    .io_vliw_in_45(pipe3_io_vliw_in_45),
    .io_vliw_in_46(pipe3_io_vliw_in_46),
    .io_vliw_in_47(pipe3_io_vliw_in_47),
    .io_vliw_in_48(pipe3_io_vliw_in_48),
    .io_vliw_in_49(pipe3_io_vliw_in_49),
    .io_vliw_in_50(pipe3_io_vliw_in_50),
    .io_vliw_in_51(pipe3_io_vliw_in_51),
    .io_vliw_in_52(pipe3_io_vliw_in_52),
    .io_vliw_in_53(pipe3_io_vliw_in_53),
    .io_vliw_in_54(pipe3_io_vliw_in_54),
    .io_vliw_in_55(pipe3_io_vliw_in_55),
    .io_vliw_in_56(pipe3_io_vliw_in_56),
    .io_vliw_in_57(pipe3_io_vliw_in_57),
    .io_vliw_in_58(pipe3_io_vliw_in_58),
    .io_vliw_in_59(pipe3_io_vliw_in_59),
    .io_vliw_in_60(pipe3_io_vliw_in_60),
    .io_vliw_in_61(pipe3_io_vliw_in_61),
    .io_vliw_in_62(pipe3_io_vliw_in_62),
    .io_vliw_in_63(pipe3_io_vliw_in_63),
    .io_vliw_in_64(pipe3_io_vliw_in_64),
    .io_vliw_in_65(pipe3_io_vliw_in_65),
    .io_vliw_in_66(pipe3_io_vliw_in_66),
    .io_vliw_in_67(pipe3_io_vliw_in_67),
    .io_vliw_in_68(pipe3_io_vliw_in_68),
    .io_vliw_in_69(pipe3_io_vliw_in_69),
    .io_nid_in(pipe3_io_nid_in),
    .io_nid_out(pipe3_io_nid_out),
    .io_tag_out_0(pipe3_io_tag_out_0),
    .io_tag_out_1(pipe3_io_tag_out_1),
    .io_tag_out_2(pipe3_io_tag_out_2),
    .io_tag_out_3(pipe3_io_tag_out_3),
    .io_tag_out_4(pipe3_io_tag_out_4),
    .io_tag_out_5(pipe3_io_tag_out_5),
    .io_tag_out_6(pipe3_io_tag_out_6),
    .io_tag_out_7(pipe3_io_tag_out_7),
    .io_tag_out_8(pipe3_io_tag_out_8),
    .io_tag_out_9(pipe3_io_tag_out_9),
    .io_tag_out_10(pipe3_io_tag_out_10),
    .io_tag_out_11(pipe3_io_tag_out_11),
    .io_tag_out_12(pipe3_io_tag_out_12),
    .io_tag_out_13(pipe3_io_tag_out_13),
    .io_tag_out_14(pipe3_io_tag_out_14),
    .io_tag_out_15(pipe3_io_tag_out_15),
    .io_tag_out_16(pipe3_io_tag_out_16),
    .io_tag_out_17(pipe3_io_tag_out_17),
    .io_tag_out_18(pipe3_io_tag_out_18),
    .io_tag_out_19(pipe3_io_tag_out_19),
    .io_tag_out_20(pipe3_io_tag_out_20),
    .io_tag_out_21(pipe3_io_tag_out_21),
    .io_tag_out_22(pipe3_io_tag_out_22),
    .io_tag_out_23(pipe3_io_tag_out_23),
    .io_tag_out_24(pipe3_io_tag_out_24),
    .io_tag_out_25(pipe3_io_tag_out_25),
    .io_tag_out_26(pipe3_io_tag_out_26),
    .io_tag_out_27(pipe3_io_tag_out_27),
    .io_tag_out_28(pipe3_io_tag_out_28),
    .io_tag_out_29(pipe3_io_tag_out_29),
    .io_tag_out_30(pipe3_io_tag_out_30),
    .io_tag_out_31(pipe3_io_tag_out_31),
    .io_tag_out_32(pipe3_io_tag_out_32),
    .io_tag_out_33(pipe3_io_tag_out_33),
    .io_tag_out_34(pipe3_io_tag_out_34),
    .io_tag_out_35(pipe3_io_tag_out_35),
    .io_tag_out_36(pipe3_io_tag_out_36),
    .io_tag_out_37(pipe3_io_tag_out_37),
    .io_tag_out_38(pipe3_io_tag_out_38),
    .io_tag_out_39(pipe3_io_tag_out_39),
    .io_tag_out_40(pipe3_io_tag_out_40),
    .io_tag_out_41(pipe3_io_tag_out_41),
    .io_tag_out_42(pipe3_io_tag_out_42),
    .io_tag_out_43(pipe3_io_tag_out_43),
    .io_tag_out_44(pipe3_io_tag_out_44),
    .io_tag_out_45(pipe3_io_tag_out_45),
    .io_tag_out_46(pipe3_io_tag_out_46),
    .io_tag_out_47(pipe3_io_tag_out_47),
    .io_tag_out_48(pipe3_io_tag_out_48),
    .io_tag_out_49(pipe3_io_tag_out_49),
    .io_tag_out_50(pipe3_io_tag_out_50),
    .io_tag_out_51(pipe3_io_tag_out_51),
    .io_tag_out_52(pipe3_io_tag_out_52),
    .io_tag_out_53(pipe3_io_tag_out_53),
    .io_tag_out_54(pipe3_io_tag_out_54),
    .io_tag_out_55(pipe3_io_tag_out_55),
    .io_tag_out_56(pipe3_io_tag_out_56),
    .io_tag_out_57(pipe3_io_tag_out_57),
    .io_tag_out_58(pipe3_io_tag_out_58),
    .io_tag_out_59(pipe3_io_tag_out_59),
    .io_tag_out_60(pipe3_io_tag_out_60),
    .io_tag_out_61(pipe3_io_tag_out_61),
    .io_tag_out_62(pipe3_io_tag_out_62),
    .io_tag_out_63(pipe3_io_tag_out_63),
    .io_tag_out_64(pipe3_io_tag_out_64),
    .io_tag_out_65(pipe3_io_tag_out_65),
    .io_tag_out_66(pipe3_io_tag_out_66),
    .io_tag_out_67(pipe3_io_tag_out_67),
    .io_tag_out_68(pipe3_io_tag_out_68),
    .io_tag_out_69(pipe3_io_tag_out_69),
    .io_field_set_field8_0(pipe3_io_field_set_field8_0),
    .io_field_set_field8_1(pipe3_io_field_set_field8_1),
    .io_field_set_field8_2(pipe3_io_field_set_field8_2),
    .io_field_set_field8_3(pipe3_io_field_set_field8_3),
    .io_field_set_field8_4(pipe3_io_field_set_field8_4),
    .io_field_set_field8_5(pipe3_io_field_set_field8_5),
    .io_field_set_field8_6(pipe3_io_field_set_field8_6),
    .io_field_set_field8_7(pipe3_io_field_set_field8_7),
    .io_field_set_field8_8(pipe3_io_field_set_field8_8),
    .io_field_set_field8_9(pipe3_io_field_set_field8_9),
    .io_field_set_field8_10(pipe3_io_field_set_field8_10),
    .io_field_set_field8_11(pipe3_io_field_set_field8_11),
    .io_field_set_field8_12(pipe3_io_field_set_field8_12),
    .io_field_set_field8_13(pipe3_io_field_set_field8_13),
    .io_field_set_field8_14(pipe3_io_field_set_field8_14),
    .io_field_set_field8_15(pipe3_io_field_set_field8_15),
    .io_field_set_field8_16(pipe3_io_field_set_field8_16),
    .io_field_set_field8_17(pipe3_io_field_set_field8_17),
    .io_field_set_field8_18(pipe3_io_field_set_field8_18),
    .io_field_set_field8_19(pipe3_io_field_set_field8_19),
    .io_field_set_field16_0(pipe3_io_field_set_field16_0),
    .io_field_set_field16_1(pipe3_io_field_set_field16_1),
    .io_field_set_field16_2(pipe3_io_field_set_field16_2),
    .io_field_set_field16_3(pipe3_io_field_set_field16_3),
    .io_field_set_field16_4(pipe3_io_field_set_field16_4),
    .io_field_set_field16_5(pipe3_io_field_set_field16_5),
    .io_field_set_field16_6(pipe3_io_field_set_field16_6),
    .io_field_set_field16_7(pipe3_io_field_set_field16_7),
    .io_field_set_field16_8(pipe3_io_field_set_field16_8),
    .io_field_set_field16_9(pipe3_io_field_set_field16_9),
    .io_field_set_field16_10(pipe3_io_field_set_field16_10),
    .io_field_set_field16_11(pipe3_io_field_set_field16_11),
    .io_field_set_field16_12(pipe3_io_field_set_field16_12),
    .io_field_set_field16_13(pipe3_io_field_set_field16_13),
    .io_field_set_field16_14(pipe3_io_field_set_field16_14),
    .io_field_set_field16_15(pipe3_io_field_set_field16_15),
    .io_field_set_field16_16(pipe3_io_field_set_field16_16),
    .io_field_set_field16_17(pipe3_io_field_set_field16_17),
    .io_field_set_field16_18(pipe3_io_field_set_field16_18),
    .io_field_set_field16_19(pipe3_io_field_set_field16_19),
    .io_field_set_field16_20(pipe3_io_field_set_field16_20),
    .io_field_set_field16_21(pipe3_io_field_set_field16_21),
    .io_field_set_field16_22(pipe3_io_field_set_field16_22),
    .io_field_set_field16_23(pipe3_io_field_set_field16_23),
    .io_field_set_field16_24(pipe3_io_field_set_field16_24),
    .io_field_set_field16_25(pipe3_io_field_set_field16_25),
    .io_field_set_field16_26(pipe3_io_field_set_field16_26),
    .io_field_set_field16_27(pipe3_io_field_set_field16_27),
    .io_field_set_field16_28(pipe3_io_field_set_field16_28),
    .io_field_set_field16_29(pipe3_io_field_set_field16_29),
    .io_field_set_field32_0(pipe3_io_field_set_field32_0),
    .io_field_set_field32_1(pipe3_io_field_set_field32_1),
    .io_field_set_field32_2(pipe3_io_field_set_field32_2),
    .io_field_set_field32_3(pipe3_io_field_set_field32_3),
    .io_field_set_field32_4(pipe3_io_field_set_field32_4),
    .io_field_set_field32_5(pipe3_io_field_set_field32_5),
    .io_field_set_field32_6(pipe3_io_field_set_field32_6),
    .io_field_set_field32_7(pipe3_io_field_set_field32_7),
    .io_field_set_field32_8(pipe3_io_field_set_field32_8),
    .io_field_set_field32_9(pipe3_io_field_set_field32_9),
    .io_field_set_field32_10(pipe3_io_field_set_field32_10),
    .io_field_set_field32_11(pipe3_io_field_set_field32_11),
    .io_field_set_field32_12(pipe3_io_field_set_field32_12),
    .io_field_set_field32_13(pipe3_io_field_set_field32_13),
    .io_field_set_field32_14(pipe3_io_field_set_field32_14),
    .io_field_set_field32_15(pipe3_io_field_set_field32_15),
    .io_field_set_field32_16(pipe3_io_field_set_field32_16),
    .io_field_set_field32_17(pipe3_io_field_set_field32_17),
    .io_field_set_field32_18(pipe3_io_field_set_field32_18),
    .io_field_set_field32_19(pipe3_io_field_set_field32_19)
  );
  PrimitiveWriteBackPISA pipe4 ( // @[executor_pisa.scala 289:23]
    .clock(pipe4_clock),
    .io_pipe_phv_in_data_0(pipe4_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe4_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe4_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe4_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe4_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe4_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe4_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe4_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe4_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe4_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe4_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe4_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe4_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe4_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe4_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe4_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe4_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe4_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe4_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe4_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe4_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe4_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe4_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe4_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe4_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe4_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe4_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe4_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe4_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe4_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe4_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe4_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe4_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe4_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe4_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe4_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe4_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe4_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe4_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe4_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe4_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe4_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe4_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe4_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe4_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe4_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe4_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe4_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe4_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe4_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe4_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe4_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe4_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe4_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe4_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe4_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe4_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe4_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe4_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe4_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe4_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe4_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe4_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe4_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe4_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe4_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe4_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe4_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe4_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe4_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe4_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe4_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe4_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe4_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe4_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe4_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe4_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe4_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe4_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe4_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe4_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe4_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe4_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe4_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe4_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe4_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe4_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe4_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe4_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe4_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe4_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe4_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe4_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe4_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe4_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe4_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe4_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe4_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe4_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe4_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe4_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe4_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe4_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe4_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe4_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe4_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe4_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe4_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe4_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe4_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe4_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe4_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe4_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe4_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe4_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe4_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe4_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe4_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe4_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe4_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe4_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe4_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe4_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe4_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe4_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe4_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe4_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe4_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe4_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe4_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe4_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe4_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe4_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe4_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe4_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe4_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe4_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe4_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe4_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe4_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe4_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe4_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe4_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe4_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe4_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe4_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe4_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe4_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe4_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe4_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe4_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe4_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe4_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe4_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe4_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe4_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe4_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe4_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe4_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe4_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_next_config_id(pipe4_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe4_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe4_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe4_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe4_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe4_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe4_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe4_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe4_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe4_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe4_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe4_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe4_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe4_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe4_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe4_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe4_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe4_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe4_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe4_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe4_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe4_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe4_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe4_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe4_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe4_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe4_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe4_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe4_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe4_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe4_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe4_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe4_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe4_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe4_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe4_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe4_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe4_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe4_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe4_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe4_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe4_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe4_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe4_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe4_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe4_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe4_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe4_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe4_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe4_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe4_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe4_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe4_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe4_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe4_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe4_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe4_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe4_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe4_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe4_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe4_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe4_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe4_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe4_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe4_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe4_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe4_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe4_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe4_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe4_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe4_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe4_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe4_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe4_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe4_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe4_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe4_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe4_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe4_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe4_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe4_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe4_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe4_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe4_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe4_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe4_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe4_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe4_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe4_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe4_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe4_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe4_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe4_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe4_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe4_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe4_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe4_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe4_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe4_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe4_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe4_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe4_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe4_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe4_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe4_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe4_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe4_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe4_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe4_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe4_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe4_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe4_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe4_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe4_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe4_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe4_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe4_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe4_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe4_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe4_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe4_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe4_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe4_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe4_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe4_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe4_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe4_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe4_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe4_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe4_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe4_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe4_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe4_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe4_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe4_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe4_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe4_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe4_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe4_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe4_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe4_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe4_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe4_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe4_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe4_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe4_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe4_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe4_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe4_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe4_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe4_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe4_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe4_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe4_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe4_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe4_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe4_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe4_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe4_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe4_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe4_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe4_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_next_config_id(pipe4_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe4_io_pipe_phv_out_is_valid_processor),
    .io_nid_in(pipe4_io_nid_in),
    .io_tag_in_0(pipe4_io_tag_in_0),
    .io_tag_in_1(pipe4_io_tag_in_1),
    .io_tag_in_2(pipe4_io_tag_in_2),
    .io_tag_in_3(pipe4_io_tag_in_3),
    .io_tag_in_4(pipe4_io_tag_in_4),
    .io_tag_in_5(pipe4_io_tag_in_5),
    .io_tag_in_6(pipe4_io_tag_in_6),
    .io_tag_in_7(pipe4_io_tag_in_7),
    .io_tag_in_8(pipe4_io_tag_in_8),
    .io_tag_in_9(pipe4_io_tag_in_9),
    .io_tag_in_10(pipe4_io_tag_in_10),
    .io_tag_in_11(pipe4_io_tag_in_11),
    .io_tag_in_12(pipe4_io_tag_in_12),
    .io_tag_in_13(pipe4_io_tag_in_13),
    .io_tag_in_14(pipe4_io_tag_in_14),
    .io_tag_in_15(pipe4_io_tag_in_15),
    .io_tag_in_16(pipe4_io_tag_in_16),
    .io_tag_in_17(pipe4_io_tag_in_17),
    .io_tag_in_18(pipe4_io_tag_in_18),
    .io_tag_in_19(pipe4_io_tag_in_19),
    .io_tag_in_20(pipe4_io_tag_in_20),
    .io_tag_in_21(pipe4_io_tag_in_21),
    .io_tag_in_22(pipe4_io_tag_in_22),
    .io_tag_in_23(pipe4_io_tag_in_23),
    .io_tag_in_24(pipe4_io_tag_in_24),
    .io_tag_in_25(pipe4_io_tag_in_25),
    .io_tag_in_26(pipe4_io_tag_in_26),
    .io_tag_in_27(pipe4_io_tag_in_27),
    .io_tag_in_28(pipe4_io_tag_in_28),
    .io_tag_in_29(pipe4_io_tag_in_29),
    .io_tag_in_30(pipe4_io_tag_in_30),
    .io_tag_in_31(pipe4_io_tag_in_31),
    .io_tag_in_32(pipe4_io_tag_in_32),
    .io_tag_in_33(pipe4_io_tag_in_33),
    .io_tag_in_34(pipe4_io_tag_in_34),
    .io_tag_in_35(pipe4_io_tag_in_35),
    .io_tag_in_36(pipe4_io_tag_in_36),
    .io_tag_in_37(pipe4_io_tag_in_37),
    .io_tag_in_38(pipe4_io_tag_in_38),
    .io_tag_in_39(pipe4_io_tag_in_39),
    .io_tag_in_40(pipe4_io_tag_in_40),
    .io_tag_in_41(pipe4_io_tag_in_41),
    .io_tag_in_42(pipe4_io_tag_in_42),
    .io_tag_in_43(pipe4_io_tag_in_43),
    .io_tag_in_44(pipe4_io_tag_in_44),
    .io_tag_in_45(pipe4_io_tag_in_45),
    .io_tag_in_46(pipe4_io_tag_in_46),
    .io_tag_in_47(pipe4_io_tag_in_47),
    .io_tag_in_48(pipe4_io_tag_in_48),
    .io_tag_in_49(pipe4_io_tag_in_49),
    .io_tag_in_50(pipe4_io_tag_in_50),
    .io_tag_in_51(pipe4_io_tag_in_51),
    .io_tag_in_52(pipe4_io_tag_in_52),
    .io_tag_in_53(pipe4_io_tag_in_53),
    .io_tag_in_54(pipe4_io_tag_in_54),
    .io_tag_in_55(pipe4_io_tag_in_55),
    .io_tag_in_56(pipe4_io_tag_in_56),
    .io_tag_in_57(pipe4_io_tag_in_57),
    .io_tag_in_58(pipe4_io_tag_in_58),
    .io_tag_in_59(pipe4_io_tag_in_59),
    .io_tag_in_60(pipe4_io_tag_in_60),
    .io_tag_in_61(pipe4_io_tag_in_61),
    .io_tag_in_62(pipe4_io_tag_in_62),
    .io_tag_in_63(pipe4_io_tag_in_63),
    .io_tag_in_64(pipe4_io_tag_in_64),
    .io_tag_in_65(pipe4_io_tag_in_65),
    .io_tag_in_66(pipe4_io_tag_in_66),
    .io_tag_in_67(pipe4_io_tag_in_67),
    .io_tag_in_68(pipe4_io_tag_in_68),
    .io_tag_in_69(pipe4_io_tag_in_69),
    .io_field_set_field8_0(pipe4_io_field_set_field8_0),
    .io_field_set_field8_1(pipe4_io_field_set_field8_1),
    .io_field_set_field8_2(pipe4_io_field_set_field8_2),
    .io_field_set_field8_3(pipe4_io_field_set_field8_3),
    .io_field_set_field8_4(pipe4_io_field_set_field8_4),
    .io_field_set_field8_5(pipe4_io_field_set_field8_5),
    .io_field_set_field8_6(pipe4_io_field_set_field8_6),
    .io_field_set_field8_7(pipe4_io_field_set_field8_7),
    .io_field_set_field8_8(pipe4_io_field_set_field8_8),
    .io_field_set_field8_9(pipe4_io_field_set_field8_9),
    .io_field_set_field8_10(pipe4_io_field_set_field8_10),
    .io_field_set_field8_11(pipe4_io_field_set_field8_11),
    .io_field_set_field8_12(pipe4_io_field_set_field8_12),
    .io_field_set_field8_13(pipe4_io_field_set_field8_13),
    .io_field_set_field8_14(pipe4_io_field_set_field8_14),
    .io_field_set_field8_15(pipe4_io_field_set_field8_15),
    .io_field_set_field8_16(pipe4_io_field_set_field8_16),
    .io_field_set_field8_17(pipe4_io_field_set_field8_17),
    .io_field_set_field8_18(pipe4_io_field_set_field8_18),
    .io_field_set_field8_19(pipe4_io_field_set_field8_19),
    .io_field_set_field16_0(pipe4_io_field_set_field16_0),
    .io_field_set_field16_1(pipe4_io_field_set_field16_1),
    .io_field_set_field16_2(pipe4_io_field_set_field16_2),
    .io_field_set_field16_3(pipe4_io_field_set_field16_3),
    .io_field_set_field16_4(pipe4_io_field_set_field16_4),
    .io_field_set_field16_5(pipe4_io_field_set_field16_5),
    .io_field_set_field16_6(pipe4_io_field_set_field16_6),
    .io_field_set_field16_7(pipe4_io_field_set_field16_7),
    .io_field_set_field16_8(pipe4_io_field_set_field16_8),
    .io_field_set_field16_9(pipe4_io_field_set_field16_9),
    .io_field_set_field16_10(pipe4_io_field_set_field16_10),
    .io_field_set_field16_11(pipe4_io_field_set_field16_11),
    .io_field_set_field16_12(pipe4_io_field_set_field16_12),
    .io_field_set_field16_13(pipe4_io_field_set_field16_13),
    .io_field_set_field16_14(pipe4_io_field_set_field16_14),
    .io_field_set_field16_15(pipe4_io_field_set_field16_15),
    .io_field_set_field16_16(pipe4_io_field_set_field16_16),
    .io_field_set_field16_17(pipe4_io_field_set_field16_17),
    .io_field_set_field16_18(pipe4_io_field_set_field16_18),
    .io_field_set_field16_19(pipe4_io_field_set_field16_19),
    .io_field_set_field16_20(pipe4_io_field_set_field16_20),
    .io_field_set_field16_21(pipe4_io_field_set_field16_21),
    .io_field_set_field16_22(pipe4_io_field_set_field16_22),
    .io_field_set_field16_23(pipe4_io_field_set_field16_23),
    .io_field_set_field16_24(pipe4_io_field_set_field16_24),
    .io_field_set_field16_25(pipe4_io_field_set_field16_25),
    .io_field_set_field16_26(pipe4_io_field_set_field16_26),
    .io_field_set_field16_27(pipe4_io_field_set_field16_27),
    .io_field_set_field16_28(pipe4_io_field_set_field16_28),
    .io_field_set_field16_29(pipe4_io_field_set_field16_29),
    .io_field_set_field32_0(pipe4_io_field_set_field32_0),
    .io_field_set_field32_1(pipe4_io_field_set_field32_1),
    .io_field_set_field32_2(pipe4_io_field_set_field32_2),
    .io_field_set_field32_3(pipe4_io_field_set_field32_3),
    .io_field_set_field32_4(pipe4_io_field_set_field32_4),
    .io_field_set_field32_5(pipe4_io_field_set_field32_5),
    .io_field_set_field32_6(pipe4_io_field_set_field32_6),
    .io_field_set_field32_7(pipe4_io_field_set_field32_7),
    .io_field_set_field32_8(pipe4_io_field_set_field32_8),
    .io_field_set_field32_9(pipe4_io_field_set_field32_9),
    .io_field_set_field32_10(pipe4_io_field_set_field32_10),
    .io_field_set_field32_11(pipe4_io_field_set_field32_11),
    .io_field_set_field32_12(pipe4_io_field_set_field32_12),
    .io_field_set_field32_13(pipe4_io_field_set_field32_13),
    .io_field_set_field32_14(pipe4_io_field_set_field32_14),
    .io_field_set_field32_15(pipe4_io_field_set_field32_15),
    .io_field_set_field32_16(pipe4_io_field_set_field32_16),
    .io_field_set_field32_17(pipe4_io_field_set_field32_17),
    .io_field_set_field32_18(pipe4_io_field_set_field32_18),
    .io_field_set_field32_19(pipe4_io_field_set_field32_19)
  );
  assign io_pipe_phv_out_data_0 = pipe4_io_pipe_phv_out_data_0; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_1 = pipe4_io_pipe_phv_out_data_1; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_2 = pipe4_io_pipe_phv_out_data_2; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_3 = pipe4_io_pipe_phv_out_data_3; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_4 = pipe4_io_pipe_phv_out_data_4; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_5 = pipe4_io_pipe_phv_out_data_5; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_6 = pipe4_io_pipe_phv_out_data_6; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_7 = pipe4_io_pipe_phv_out_data_7; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_8 = pipe4_io_pipe_phv_out_data_8; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_9 = pipe4_io_pipe_phv_out_data_9; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_10 = pipe4_io_pipe_phv_out_data_10; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_11 = pipe4_io_pipe_phv_out_data_11; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_12 = pipe4_io_pipe_phv_out_data_12; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_13 = pipe4_io_pipe_phv_out_data_13; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_14 = pipe4_io_pipe_phv_out_data_14; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_15 = pipe4_io_pipe_phv_out_data_15; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_16 = pipe4_io_pipe_phv_out_data_16; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_17 = pipe4_io_pipe_phv_out_data_17; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_18 = pipe4_io_pipe_phv_out_data_18; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_19 = pipe4_io_pipe_phv_out_data_19; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_20 = pipe4_io_pipe_phv_out_data_20; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_21 = pipe4_io_pipe_phv_out_data_21; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_22 = pipe4_io_pipe_phv_out_data_22; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_23 = pipe4_io_pipe_phv_out_data_23; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_24 = pipe4_io_pipe_phv_out_data_24; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_25 = pipe4_io_pipe_phv_out_data_25; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_26 = pipe4_io_pipe_phv_out_data_26; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_27 = pipe4_io_pipe_phv_out_data_27; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_28 = pipe4_io_pipe_phv_out_data_28; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_29 = pipe4_io_pipe_phv_out_data_29; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_30 = pipe4_io_pipe_phv_out_data_30; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_31 = pipe4_io_pipe_phv_out_data_31; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_32 = pipe4_io_pipe_phv_out_data_32; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_33 = pipe4_io_pipe_phv_out_data_33; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_34 = pipe4_io_pipe_phv_out_data_34; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_35 = pipe4_io_pipe_phv_out_data_35; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_36 = pipe4_io_pipe_phv_out_data_36; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_37 = pipe4_io_pipe_phv_out_data_37; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_38 = pipe4_io_pipe_phv_out_data_38; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_39 = pipe4_io_pipe_phv_out_data_39; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_40 = pipe4_io_pipe_phv_out_data_40; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_41 = pipe4_io_pipe_phv_out_data_41; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_42 = pipe4_io_pipe_phv_out_data_42; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_43 = pipe4_io_pipe_phv_out_data_43; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_44 = pipe4_io_pipe_phv_out_data_44; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_45 = pipe4_io_pipe_phv_out_data_45; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_46 = pipe4_io_pipe_phv_out_data_46; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_47 = pipe4_io_pipe_phv_out_data_47; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_48 = pipe4_io_pipe_phv_out_data_48; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_49 = pipe4_io_pipe_phv_out_data_49; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_50 = pipe4_io_pipe_phv_out_data_50; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_51 = pipe4_io_pipe_phv_out_data_51; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_52 = pipe4_io_pipe_phv_out_data_52; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_53 = pipe4_io_pipe_phv_out_data_53; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_54 = pipe4_io_pipe_phv_out_data_54; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_55 = pipe4_io_pipe_phv_out_data_55; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_56 = pipe4_io_pipe_phv_out_data_56; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_57 = pipe4_io_pipe_phv_out_data_57; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_58 = pipe4_io_pipe_phv_out_data_58; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_59 = pipe4_io_pipe_phv_out_data_59; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_60 = pipe4_io_pipe_phv_out_data_60; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_61 = pipe4_io_pipe_phv_out_data_61; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_62 = pipe4_io_pipe_phv_out_data_62; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_63 = pipe4_io_pipe_phv_out_data_63; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_64 = pipe4_io_pipe_phv_out_data_64; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_65 = pipe4_io_pipe_phv_out_data_65; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_66 = pipe4_io_pipe_phv_out_data_66; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_67 = pipe4_io_pipe_phv_out_data_67; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_68 = pipe4_io_pipe_phv_out_data_68; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_69 = pipe4_io_pipe_phv_out_data_69; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_70 = pipe4_io_pipe_phv_out_data_70; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_71 = pipe4_io_pipe_phv_out_data_71; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_72 = pipe4_io_pipe_phv_out_data_72; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_73 = pipe4_io_pipe_phv_out_data_73; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_74 = pipe4_io_pipe_phv_out_data_74; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_75 = pipe4_io_pipe_phv_out_data_75; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_76 = pipe4_io_pipe_phv_out_data_76; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_77 = pipe4_io_pipe_phv_out_data_77; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_78 = pipe4_io_pipe_phv_out_data_78; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_79 = pipe4_io_pipe_phv_out_data_79; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_80 = pipe4_io_pipe_phv_out_data_80; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_81 = pipe4_io_pipe_phv_out_data_81; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_82 = pipe4_io_pipe_phv_out_data_82; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_83 = pipe4_io_pipe_phv_out_data_83; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_84 = pipe4_io_pipe_phv_out_data_84; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_85 = pipe4_io_pipe_phv_out_data_85; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_86 = pipe4_io_pipe_phv_out_data_86; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_87 = pipe4_io_pipe_phv_out_data_87; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_88 = pipe4_io_pipe_phv_out_data_88; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_89 = pipe4_io_pipe_phv_out_data_89; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_90 = pipe4_io_pipe_phv_out_data_90; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_91 = pipe4_io_pipe_phv_out_data_91; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_92 = pipe4_io_pipe_phv_out_data_92; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_93 = pipe4_io_pipe_phv_out_data_93; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_94 = pipe4_io_pipe_phv_out_data_94; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_95 = pipe4_io_pipe_phv_out_data_95; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_96 = pipe4_io_pipe_phv_out_data_96; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_97 = pipe4_io_pipe_phv_out_data_97; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_98 = pipe4_io_pipe_phv_out_data_98; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_99 = pipe4_io_pipe_phv_out_data_99; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_100 = pipe4_io_pipe_phv_out_data_100; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_101 = pipe4_io_pipe_phv_out_data_101; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_102 = pipe4_io_pipe_phv_out_data_102; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_103 = pipe4_io_pipe_phv_out_data_103; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_104 = pipe4_io_pipe_phv_out_data_104; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_105 = pipe4_io_pipe_phv_out_data_105; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_106 = pipe4_io_pipe_phv_out_data_106; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_107 = pipe4_io_pipe_phv_out_data_107; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_108 = pipe4_io_pipe_phv_out_data_108; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_109 = pipe4_io_pipe_phv_out_data_109; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_110 = pipe4_io_pipe_phv_out_data_110; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_111 = pipe4_io_pipe_phv_out_data_111; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_112 = pipe4_io_pipe_phv_out_data_112; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_113 = pipe4_io_pipe_phv_out_data_113; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_114 = pipe4_io_pipe_phv_out_data_114; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_115 = pipe4_io_pipe_phv_out_data_115; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_116 = pipe4_io_pipe_phv_out_data_116; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_117 = pipe4_io_pipe_phv_out_data_117; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_118 = pipe4_io_pipe_phv_out_data_118; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_119 = pipe4_io_pipe_phv_out_data_119; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_120 = pipe4_io_pipe_phv_out_data_120; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_121 = pipe4_io_pipe_phv_out_data_121; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_122 = pipe4_io_pipe_phv_out_data_122; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_123 = pipe4_io_pipe_phv_out_data_123; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_124 = pipe4_io_pipe_phv_out_data_124; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_125 = pipe4_io_pipe_phv_out_data_125; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_126 = pipe4_io_pipe_phv_out_data_126; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_127 = pipe4_io_pipe_phv_out_data_127; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_128 = pipe4_io_pipe_phv_out_data_128; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_129 = pipe4_io_pipe_phv_out_data_129; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_130 = pipe4_io_pipe_phv_out_data_130; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_131 = pipe4_io_pipe_phv_out_data_131; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_132 = pipe4_io_pipe_phv_out_data_132; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_133 = pipe4_io_pipe_phv_out_data_133; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_134 = pipe4_io_pipe_phv_out_data_134; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_135 = pipe4_io_pipe_phv_out_data_135; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_136 = pipe4_io_pipe_phv_out_data_136; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_137 = pipe4_io_pipe_phv_out_data_137; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_138 = pipe4_io_pipe_phv_out_data_138; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_139 = pipe4_io_pipe_phv_out_data_139; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_140 = pipe4_io_pipe_phv_out_data_140; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_141 = pipe4_io_pipe_phv_out_data_141; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_142 = pipe4_io_pipe_phv_out_data_142; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_143 = pipe4_io_pipe_phv_out_data_143; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_144 = pipe4_io_pipe_phv_out_data_144; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_145 = pipe4_io_pipe_phv_out_data_145; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_146 = pipe4_io_pipe_phv_out_data_146; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_147 = pipe4_io_pipe_phv_out_data_147; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_148 = pipe4_io_pipe_phv_out_data_148; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_149 = pipe4_io_pipe_phv_out_data_149; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_150 = pipe4_io_pipe_phv_out_data_150; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_151 = pipe4_io_pipe_phv_out_data_151; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_152 = pipe4_io_pipe_phv_out_data_152; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_153 = pipe4_io_pipe_phv_out_data_153; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_154 = pipe4_io_pipe_phv_out_data_154; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_155 = pipe4_io_pipe_phv_out_data_155; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_156 = pipe4_io_pipe_phv_out_data_156; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_157 = pipe4_io_pipe_phv_out_data_157; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_158 = pipe4_io_pipe_phv_out_data_158; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_data_159 = pipe4_io_pipe_phv_out_data_159; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_next_config_id = pipe4_io_pipe_phv_out_next_config_id; // @[executor_pisa.scala 310:27]
  assign io_pipe_phv_out_is_valid_processor = pipe4_io_pipe_phv_out_is_valid_processor; // @[executor_pisa.scala 310:27]
  assign pipe1_clock = clock;
  assign pipe1_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_96 = io_pipe_phv_in_data_96; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_97 = io_pipe_phv_in_data_97; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_98 = io_pipe_phv_in_data_98; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_99 = io_pipe_phv_in_data_99; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_100 = io_pipe_phv_in_data_100; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_101 = io_pipe_phv_in_data_101; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_102 = io_pipe_phv_in_data_102; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_103 = io_pipe_phv_in_data_103; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_104 = io_pipe_phv_in_data_104; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_105 = io_pipe_phv_in_data_105; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_106 = io_pipe_phv_in_data_106; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_107 = io_pipe_phv_in_data_107; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_108 = io_pipe_phv_in_data_108; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_109 = io_pipe_phv_in_data_109; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_110 = io_pipe_phv_in_data_110; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_111 = io_pipe_phv_in_data_111; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_112 = io_pipe_phv_in_data_112; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_113 = io_pipe_phv_in_data_113; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_114 = io_pipe_phv_in_data_114; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_115 = io_pipe_phv_in_data_115; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_116 = io_pipe_phv_in_data_116; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_117 = io_pipe_phv_in_data_117; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_118 = io_pipe_phv_in_data_118; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_119 = io_pipe_phv_in_data_119; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_120 = io_pipe_phv_in_data_120; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_121 = io_pipe_phv_in_data_121; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_122 = io_pipe_phv_in_data_122; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_123 = io_pipe_phv_in_data_123; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_124 = io_pipe_phv_in_data_124; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_125 = io_pipe_phv_in_data_125; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_126 = io_pipe_phv_in_data_126; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_127 = io_pipe_phv_in_data_127; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_128 = io_pipe_phv_in_data_128; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_129 = io_pipe_phv_in_data_129; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_130 = io_pipe_phv_in_data_130; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_131 = io_pipe_phv_in_data_131; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_132 = io_pipe_phv_in_data_132; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_133 = io_pipe_phv_in_data_133; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_134 = io_pipe_phv_in_data_134; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_135 = io_pipe_phv_in_data_135; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_136 = io_pipe_phv_in_data_136; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_137 = io_pipe_phv_in_data_137; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_138 = io_pipe_phv_in_data_138; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_139 = io_pipe_phv_in_data_139; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_140 = io_pipe_phv_in_data_140; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_141 = io_pipe_phv_in_data_141; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_142 = io_pipe_phv_in_data_142; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_143 = io_pipe_phv_in_data_143; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_144 = io_pipe_phv_in_data_144; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_145 = io_pipe_phv_in_data_145; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_146 = io_pipe_phv_in_data_146; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_147 = io_pipe_phv_in_data_147; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_148 = io_pipe_phv_in_data_148; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_149 = io_pipe_phv_in_data_149; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_150 = io_pipe_phv_in_data_150; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_151 = io_pipe_phv_in_data_151; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_152 = io_pipe_phv_in_data_152; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_153 = io_pipe_phv_in_data_153; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_154 = io_pipe_phv_in_data_154; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_155 = io_pipe_phv_in_data_155; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_156 = io_pipe_phv_in_data_156; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_157 = io_pipe_phv_in_data_157; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_158 = io_pipe_phv_in_data_158; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_data_159 = io_pipe_phv_in_data_159; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_next_config_id = io_pipe_phv_in_next_config_id; // @[executor_pisa.scala 291:26]
  assign pipe1_io_pipe_phv_in_is_valid_processor = io_pipe_phv_in_is_valid_processor; // @[executor_pisa.scala 291:26]
  assign pipe1_io_hit = io_hit; // @[executor_pisa.scala 292:26]
  assign pipe1_io_match_value = io_match_value; // @[executor_pisa.scala 293:26]
  assign pipe1_io_action_mod_en_0 = io_action_mod_en_0; // @[executor_pisa.scala 294:26]
  assign pipe1_io_action_mod_en_1 = io_action_mod_en_1; // @[executor_pisa.scala 294:26]
  assign pipe1_io_action_mod_addr = io_action_mod_addr; // @[executor_pisa.scala 294:26]
  assign pipe1_io_action_mod_data_0 = io_action_mod_data_0; // @[executor_pisa.scala 294:26]
  assign pipe1_io_action_mod_data_1 = io_action_mod_data_1; // @[executor_pisa.scala 294:26]
  assign pipe2_clock = clock;
  assign pipe2_io_pipe_phv_in_data_0 = pipe1_io_pipe_phv_out_data_0; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_1 = pipe1_io_pipe_phv_out_data_1; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_2 = pipe1_io_pipe_phv_out_data_2; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_3 = pipe1_io_pipe_phv_out_data_3; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_4 = pipe1_io_pipe_phv_out_data_4; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_5 = pipe1_io_pipe_phv_out_data_5; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_6 = pipe1_io_pipe_phv_out_data_6; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_7 = pipe1_io_pipe_phv_out_data_7; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_8 = pipe1_io_pipe_phv_out_data_8; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_9 = pipe1_io_pipe_phv_out_data_9; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_10 = pipe1_io_pipe_phv_out_data_10; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_11 = pipe1_io_pipe_phv_out_data_11; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_12 = pipe1_io_pipe_phv_out_data_12; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_13 = pipe1_io_pipe_phv_out_data_13; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_14 = pipe1_io_pipe_phv_out_data_14; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_15 = pipe1_io_pipe_phv_out_data_15; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_16 = pipe1_io_pipe_phv_out_data_16; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_17 = pipe1_io_pipe_phv_out_data_17; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_18 = pipe1_io_pipe_phv_out_data_18; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_19 = pipe1_io_pipe_phv_out_data_19; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_20 = pipe1_io_pipe_phv_out_data_20; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_21 = pipe1_io_pipe_phv_out_data_21; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_22 = pipe1_io_pipe_phv_out_data_22; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_23 = pipe1_io_pipe_phv_out_data_23; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_24 = pipe1_io_pipe_phv_out_data_24; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_25 = pipe1_io_pipe_phv_out_data_25; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_26 = pipe1_io_pipe_phv_out_data_26; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_27 = pipe1_io_pipe_phv_out_data_27; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_28 = pipe1_io_pipe_phv_out_data_28; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_29 = pipe1_io_pipe_phv_out_data_29; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_30 = pipe1_io_pipe_phv_out_data_30; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_31 = pipe1_io_pipe_phv_out_data_31; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_32 = pipe1_io_pipe_phv_out_data_32; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_33 = pipe1_io_pipe_phv_out_data_33; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_34 = pipe1_io_pipe_phv_out_data_34; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_35 = pipe1_io_pipe_phv_out_data_35; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_36 = pipe1_io_pipe_phv_out_data_36; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_37 = pipe1_io_pipe_phv_out_data_37; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_38 = pipe1_io_pipe_phv_out_data_38; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_39 = pipe1_io_pipe_phv_out_data_39; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_40 = pipe1_io_pipe_phv_out_data_40; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_41 = pipe1_io_pipe_phv_out_data_41; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_42 = pipe1_io_pipe_phv_out_data_42; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_43 = pipe1_io_pipe_phv_out_data_43; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_44 = pipe1_io_pipe_phv_out_data_44; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_45 = pipe1_io_pipe_phv_out_data_45; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_46 = pipe1_io_pipe_phv_out_data_46; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_47 = pipe1_io_pipe_phv_out_data_47; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_48 = pipe1_io_pipe_phv_out_data_48; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_49 = pipe1_io_pipe_phv_out_data_49; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_50 = pipe1_io_pipe_phv_out_data_50; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_51 = pipe1_io_pipe_phv_out_data_51; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_52 = pipe1_io_pipe_phv_out_data_52; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_53 = pipe1_io_pipe_phv_out_data_53; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_54 = pipe1_io_pipe_phv_out_data_54; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_55 = pipe1_io_pipe_phv_out_data_55; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_56 = pipe1_io_pipe_phv_out_data_56; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_57 = pipe1_io_pipe_phv_out_data_57; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_58 = pipe1_io_pipe_phv_out_data_58; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_59 = pipe1_io_pipe_phv_out_data_59; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_60 = pipe1_io_pipe_phv_out_data_60; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_61 = pipe1_io_pipe_phv_out_data_61; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_62 = pipe1_io_pipe_phv_out_data_62; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_63 = pipe1_io_pipe_phv_out_data_63; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_64 = pipe1_io_pipe_phv_out_data_64; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_65 = pipe1_io_pipe_phv_out_data_65; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_66 = pipe1_io_pipe_phv_out_data_66; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_67 = pipe1_io_pipe_phv_out_data_67; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_68 = pipe1_io_pipe_phv_out_data_68; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_69 = pipe1_io_pipe_phv_out_data_69; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_70 = pipe1_io_pipe_phv_out_data_70; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_71 = pipe1_io_pipe_phv_out_data_71; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_72 = pipe1_io_pipe_phv_out_data_72; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_73 = pipe1_io_pipe_phv_out_data_73; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_74 = pipe1_io_pipe_phv_out_data_74; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_75 = pipe1_io_pipe_phv_out_data_75; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_76 = pipe1_io_pipe_phv_out_data_76; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_77 = pipe1_io_pipe_phv_out_data_77; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_78 = pipe1_io_pipe_phv_out_data_78; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_79 = pipe1_io_pipe_phv_out_data_79; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_80 = pipe1_io_pipe_phv_out_data_80; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_81 = pipe1_io_pipe_phv_out_data_81; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_82 = pipe1_io_pipe_phv_out_data_82; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_83 = pipe1_io_pipe_phv_out_data_83; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_84 = pipe1_io_pipe_phv_out_data_84; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_85 = pipe1_io_pipe_phv_out_data_85; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_86 = pipe1_io_pipe_phv_out_data_86; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_87 = pipe1_io_pipe_phv_out_data_87; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_88 = pipe1_io_pipe_phv_out_data_88; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_89 = pipe1_io_pipe_phv_out_data_89; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_90 = pipe1_io_pipe_phv_out_data_90; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_91 = pipe1_io_pipe_phv_out_data_91; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_92 = pipe1_io_pipe_phv_out_data_92; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_93 = pipe1_io_pipe_phv_out_data_93; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_94 = pipe1_io_pipe_phv_out_data_94; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_95 = pipe1_io_pipe_phv_out_data_95; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_96 = pipe1_io_pipe_phv_out_data_96; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_97 = pipe1_io_pipe_phv_out_data_97; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_98 = pipe1_io_pipe_phv_out_data_98; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_99 = pipe1_io_pipe_phv_out_data_99; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_100 = pipe1_io_pipe_phv_out_data_100; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_101 = pipe1_io_pipe_phv_out_data_101; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_102 = pipe1_io_pipe_phv_out_data_102; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_103 = pipe1_io_pipe_phv_out_data_103; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_104 = pipe1_io_pipe_phv_out_data_104; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_105 = pipe1_io_pipe_phv_out_data_105; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_106 = pipe1_io_pipe_phv_out_data_106; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_107 = pipe1_io_pipe_phv_out_data_107; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_108 = pipe1_io_pipe_phv_out_data_108; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_109 = pipe1_io_pipe_phv_out_data_109; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_110 = pipe1_io_pipe_phv_out_data_110; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_111 = pipe1_io_pipe_phv_out_data_111; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_112 = pipe1_io_pipe_phv_out_data_112; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_113 = pipe1_io_pipe_phv_out_data_113; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_114 = pipe1_io_pipe_phv_out_data_114; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_115 = pipe1_io_pipe_phv_out_data_115; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_116 = pipe1_io_pipe_phv_out_data_116; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_117 = pipe1_io_pipe_phv_out_data_117; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_118 = pipe1_io_pipe_phv_out_data_118; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_119 = pipe1_io_pipe_phv_out_data_119; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_120 = pipe1_io_pipe_phv_out_data_120; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_121 = pipe1_io_pipe_phv_out_data_121; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_122 = pipe1_io_pipe_phv_out_data_122; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_123 = pipe1_io_pipe_phv_out_data_123; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_124 = pipe1_io_pipe_phv_out_data_124; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_125 = pipe1_io_pipe_phv_out_data_125; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_126 = pipe1_io_pipe_phv_out_data_126; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_127 = pipe1_io_pipe_phv_out_data_127; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_128 = pipe1_io_pipe_phv_out_data_128; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_129 = pipe1_io_pipe_phv_out_data_129; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_130 = pipe1_io_pipe_phv_out_data_130; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_131 = pipe1_io_pipe_phv_out_data_131; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_132 = pipe1_io_pipe_phv_out_data_132; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_133 = pipe1_io_pipe_phv_out_data_133; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_134 = pipe1_io_pipe_phv_out_data_134; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_135 = pipe1_io_pipe_phv_out_data_135; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_136 = pipe1_io_pipe_phv_out_data_136; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_137 = pipe1_io_pipe_phv_out_data_137; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_138 = pipe1_io_pipe_phv_out_data_138; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_139 = pipe1_io_pipe_phv_out_data_139; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_140 = pipe1_io_pipe_phv_out_data_140; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_141 = pipe1_io_pipe_phv_out_data_141; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_142 = pipe1_io_pipe_phv_out_data_142; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_143 = pipe1_io_pipe_phv_out_data_143; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_144 = pipe1_io_pipe_phv_out_data_144; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_145 = pipe1_io_pipe_phv_out_data_145; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_146 = pipe1_io_pipe_phv_out_data_146; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_147 = pipe1_io_pipe_phv_out_data_147; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_148 = pipe1_io_pipe_phv_out_data_148; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_149 = pipe1_io_pipe_phv_out_data_149; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_150 = pipe1_io_pipe_phv_out_data_150; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_151 = pipe1_io_pipe_phv_out_data_151; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_152 = pipe1_io_pipe_phv_out_data_152; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_153 = pipe1_io_pipe_phv_out_data_153; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_154 = pipe1_io_pipe_phv_out_data_154; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_155 = pipe1_io_pipe_phv_out_data_155; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_156 = pipe1_io_pipe_phv_out_data_156; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_157 = pipe1_io_pipe_phv_out_data_157; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_158 = pipe1_io_pipe_phv_out_data_158; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_data_159 = pipe1_io_pipe_phv_out_data_159; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_next_config_id = pipe1_io_pipe_phv_out_next_config_id; // @[executor_pisa.scala 296:26]
  assign pipe2_io_pipe_phv_in_is_valid_processor = pipe1_io_pipe_phv_out_is_valid_processor; // @[executor_pisa.scala 296:26]
  assign pipe2_io_args_in_0 = pipe1_io_args_out_0; // @[executor_pisa.scala 297:26]
  assign pipe2_io_args_in_1 = pipe1_io_args_out_1; // @[executor_pisa.scala 297:26]
  assign pipe2_io_args_in_2 = pipe1_io_args_out_2; // @[executor_pisa.scala 297:26]
  assign pipe2_io_args_in_3 = pipe1_io_args_out_3; // @[executor_pisa.scala 297:26]
  assign pipe2_io_args_in_4 = pipe1_io_args_out_4; // @[executor_pisa.scala 297:26]
  assign pipe2_io_args_in_5 = pipe1_io_args_out_5; // @[executor_pisa.scala 297:26]
  assign pipe2_io_args_in_6 = pipe1_io_args_out_6; // @[executor_pisa.scala 297:26]
  assign pipe2_io_vliw_in_0 = pipe1_io_vliw_out_0; // @[executor_pisa.scala 298:26]
  assign pipe2_io_vliw_in_1 = pipe1_io_vliw_out_1; // @[executor_pisa.scala 298:26]
  assign pipe2_io_vliw_in_2 = pipe1_io_vliw_out_2; // @[executor_pisa.scala 298:26]
  assign pipe2_io_vliw_in_3 = pipe1_io_vliw_out_3; // @[executor_pisa.scala 298:26]
  assign pipe3_clock = clock;
  assign pipe3_io_pipe_phv_in_data_0 = pipe2_io_pipe_phv_out_data_0; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_1 = pipe2_io_pipe_phv_out_data_1; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_2 = pipe2_io_pipe_phv_out_data_2; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_3 = pipe2_io_pipe_phv_out_data_3; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_4 = pipe2_io_pipe_phv_out_data_4; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_5 = pipe2_io_pipe_phv_out_data_5; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_6 = pipe2_io_pipe_phv_out_data_6; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_7 = pipe2_io_pipe_phv_out_data_7; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_8 = pipe2_io_pipe_phv_out_data_8; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_9 = pipe2_io_pipe_phv_out_data_9; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_10 = pipe2_io_pipe_phv_out_data_10; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_11 = pipe2_io_pipe_phv_out_data_11; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_12 = pipe2_io_pipe_phv_out_data_12; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_13 = pipe2_io_pipe_phv_out_data_13; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_14 = pipe2_io_pipe_phv_out_data_14; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_15 = pipe2_io_pipe_phv_out_data_15; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_16 = pipe2_io_pipe_phv_out_data_16; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_17 = pipe2_io_pipe_phv_out_data_17; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_18 = pipe2_io_pipe_phv_out_data_18; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_19 = pipe2_io_pipe_phv_out_data_19; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_20 = pipe2_io_pipe_phv_out_data_20; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_21 = pipe2_io_pipe_phv_out_data_21; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_22 = pipe2_io_pipe_phv_out_data_22; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_23 = pipe2_io_pipe_phv_out_data_23; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_24 = pipe2_io_pipe_phv_out_data_24; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_25 = pipe2_io_pipe_phv_out_data_25; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_26 = pipe2_io_pipe_phv_out_data_26; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_27 = pipe2_io_pipe_phv_out_data_27; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_28 = pipe2_io_pipe_phv_out_data_28; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_29 = pipe2_io_pipe_phv_out_data_29; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_30 = pipe2_io_pipe_phv_out_data_30; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_31 = pipe2_io_pipe_phv_out_data_31; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_32 = pipe2_io_pipe_phv_out_data_32; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_33 = pipe2_io_pipe_phv_out_data_33; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_34 = pipe2_io_pipe_phv_out_data_34; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_35 = pipe2_io_pipe_phv_out_data_35; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_36 = pipe2_io_pipe_phv_out_data_36; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_37 = pipe2_io_pipe_phv_out_data_37; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_38 = pipe2_io_pipe_phv_out_data_38; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_39 = pipe2_io_pipe_phv_out_data_39; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_40 = pipe2_io_pipe_phv_out_data_40; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_41 = pipe2_io_pipe_phv_out_data_41; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_42 = pipe2_io_pipe_phv_out_data_42; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_43 = pipe2_io_pipe_phv_out_data_43; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_44 = pipe2_io_pipe_phv_out_data_44; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_45 = pipe2_io_pipe_phv_out_data_45; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_46 = pipe2_io_pipe_phv_out_data_46; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_47 = pipe2_io_pipe_phv_out_data_47; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_48 = pipe2_io_pipe_phv_out_data_48; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_49 = pipe2_io_pipe_phv_out_data_49; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_50 = pipe2_io_pipe_phv_out_data_50; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_51 = pipe2_io_pipe_phv_out_data_51; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_52 = pipe2_io_pipe_phv_out_data_52; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_53 = pipe2_io_pipe_phv_out_data_53; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_54 = pipe2_io_pipe_phv_out_data_54; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_55 = pipe2_io_pipe_phv_out_data_55; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_56 = pipe2_io_pipe_phv_out_data_56; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_57 = pipe2_io_pipe_phv_out_data_57; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_58 = pipe2_io_pipe_phv_out_data_58; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_59 = pipe2_io_pipe_phv_out_data_59; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_60 = pipe2_io_pipe_phv_out_data_60; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_61 = pipe2_io_pipe_phv_out_data_61; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_62 = pipe2_io_pipe_phv_out_data_62; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_63 = pipe2_io_pipe_phv_out_data_63; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_64 = pipe2_io_pipe_phv_out_data_64; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_65 = pipe2_io_pipe_phv_out_data_65; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_66 = pipe2_io_pipe_phv_out_data_66; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_67 = pipe2_io_pipe_phv_out_data_67; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_68 = pipe2_io_pipe_phv_out_data_68; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_69 = pipe2_io_pipe_phv_out_data_69; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_70 = pipe2_io_pipe_phv_out_data_70; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_71 = pipe2_io_pipe_phv_out_data_71; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_72 = pipe2_io_pipe_phv_out_data_72; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_73 = pipe2_io_pipe_phv_out_data_73; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_74 = pipe2_io_pipe_phv_out_data_74; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_75 = pipe2_io_pipe_phv_out_data_75; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_76 = pipe2_io_pipe_phv_out_data_76; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_77 = pipe2_io_pipe_phv_out_data_77; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_78 = pipe2_io_pipe_phv_out_data_78; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_79 = pipe2_io_pipe_phv_out_data_79; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_80 = pipe2_io_pipe_phv_out_data_80; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_81 = pipe2_io_pipe_phv_out_data_81; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_82 = pipe2_io_pipe_phv_out_data_82; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_83 = pipe2_io_pipe_phv_out_data_83; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_84 = pipe2_io_pipe_phv_out_data_84; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_85 = pipe2_io_pipe_phv_out_data_85; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_86 = pipe2_io_pipe_phv_out_data_86; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_87 = pipe2_io_pipe_phv_out_data_87; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_88 = pipe2_io_pipe_phv_out_data_88; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_89 = pipe2_io_pipe_phv_out_data_89; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_90 = pipe2_io_pipe_phv_out_data_90; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_91 = pipe2_io_pipe_phv_out_data_91; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_92 = pipe2_io_pipe_phv_out_data_92; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_93 = pipe2_io_pipe_phv_out_data_93; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_94 = pipe2_io_pipe_phv_out_data_94; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_95 = pipe2_io_pipe_phv_out_data_95; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_96 = pipe2_io_pipe_phv_out_data_96; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_97 = pipe2_io_pipe_phv_out_data_97; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_98 = pipe2_io_pipe_phv_out_data_98; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_99 = pipe2_io_pipe_phv_out_data_99; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_100 = pipe2_io_pipe_phv_out_data_100; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_101 = pipe2_io_pipe_phv_out_data_101; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_102 = pipe2_io_pipe_phv_out_data_102; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_103 = pipe2_io_pipe_phv_out_data_103; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_104 = pipe2_io_pipe_phv_out_data_104; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_105 = pipe2_io_pipe_phv_out_data_105; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_106 = pipe2_io_pipe_phv_out_data_106; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_107 = pipe2_io_pipe_phv_out_data_107; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_108 = pipe2_io_pipe_phv_out_data_108; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_109 = pipe2_io_pipe_phv_out_data_109; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_110 = pipe2_io_pipe_phv_out_data_110; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_111 = pipe2_io_pipe_phv_out_data_111; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_112 = pipe2_io_pipe_phv_out_data_112; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_113 = pipe2_io_pipe_phv_out_data_113; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_114 = pipe2_io_pipe_phv_out_data_114; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_115 = pipe2_io_pipe_phv_out_data_115; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_116 = pipe2_io_pipe_phv_out_data_116; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_117 = pipe2_io_pipe_phv_out_data_117; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_118 = pipe2_io_pipe_phv_out_data_118; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_119 = pipe2_io_pipe_phv_out_data_119; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_120 = pipe2_io_pipe_phv_out_data_120; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_121 = pipe2_io_pipe_phv_out_data_121; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_122 = pipe2_io_pipe_phv_out_data_122; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_123 = pipe2_io_pipe_phv_out_data_123; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_124 = pipe2_io_pipe_phv_out_data_124; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_125 = pipe2_io_pipe_phv_out_data_125; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_126 = pipe2_io_pipe_phv_out_data_126; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_127 = pipe2_io_pipe_phv_out_data_127; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_128 = pipe2_io_pipe_phv_out_data_128; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_129 = pipe2_io_pipe_phv_out_data_129; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_130 = pipe2_io_pipe_phv_out_data_130; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_131 = pipe2_io_pipe_phv_out_data_131; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_132 = pipe2_io_pipe_phv_out_data_132; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_133 = pipe2_io_pipe_phv_out_data_133; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_134 = pipe2_io_pipe_phv_out_data_134; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_135 = pipe2_io_pipe_phv_out_data_135; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_136 = pipe2_io_pipe_phv_out_data_136; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_137 = pipe2_io_pipe_phv_out_data_137; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_138 = pipe2_io_pipe_phv_out_data_138; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_139 = pipe2_io_pipe_phv_out_data_139; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_140 = pipe2_io_pipe_phv_out_data_140; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_141 = pipe2_io_pipe_phv_out_data_141; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_142 = pipe2_io_pipe_phv_out_data_142; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_143 = pipe2_io_pipe_phv_out_data_143; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_144 = pipe2_io_pipe_phv_out_data_144; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_145 = pipe2_io_pipe_phv_out_data_145; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_146 = pipe2_io_pipe_phv_out_data_146; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_147 = pipe2_io_pipe_phv_out_data_147; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_148 = pipe2_io_pipe_phv_out_data_148; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_149 = pipe2_io_pipe_phv_out_data_149; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_150 = pipe2_io_pipe_phv_out_data_150; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_151 = pipe2_io_pipe_phv_out_data_151; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_152 = pipe2_io_pipe_phv_out_data_152; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_153 = pipe2_io_pipe_phv_out_data_153; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_154 = pipe2_io_pipe_phv_out_data_154; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_155 = pipe2_io_pipe_phv_out_data_155; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_156 = pipe2_io_pipe_phv_out_data_156; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_157 = pipe2_io_pipe_phv_out_data_157; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_158 = pipe2_io_pipe_phv_out_data_158; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_data_159 = pipe2_io_pipe_phv_out_data_159; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_next_config_id = pipe2_io_pipe_phv_out_next_config_id; // @[executor_pisa.scala 300:26]
  assign pipe3_io_pipe_phv_in_is_valid_processor = pipe2_io_pipe_phv_out_is_valid_processor; // @[executor_pisa.scala 300:26]
  assign pipe3_io_args_in_0 = pipe2_io_args_out_0; // @[executor_pisa.scala 301:26]
  assign pipe3_io_args_in_1 = pipe2_io_args_out_1; // @[executor_pisa.scala 301:26]
  assign pipe3_io_args_in_2 = pipe2_io_args_out_2; // @[executor_pisa.scala 301:26]
  assign pipe3_io_args_in_3 = pipe2_io_args_out_3; // @[executor_pisa.scala 301:26]
  assign pipe3_io_args_in_4 = pipe2_io_args_out_4; // @[executor_pisa.scala 301:26]
  assign pipe3_io_args_in_5 = pipe2_io_args_out_5; // @[executor_pisa.scala 301:26]
  assign pipe3_io_args_in_6 = pipe2_io_args_out_6; // @[executor_pisa.scala 301:26]
  assign pipe3_io_vliw_in_0 = pipe2_io_vliw_out_0; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_1 = pipe2_io_vliw_out_1; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_2 = pipe2_io_vliw_out_2; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_3 = pipe2_io_vliw_out_3; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_4 = pipe2_io_vliw_out_4; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_5 = pipe2_io_vliw_out_5; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_6 = pipe2_io_vliw_out_6; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_7 = pipe2_io_vliw_out_7; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_8 = pipe2_io_vliw_out_8; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_9 = pipe2_io_vliw_out_9; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_10 = pipe2_io_vliw_out_10; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_11 = pipe2_io_vliw_out_11; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_12 = pipe2_io_vliw_out_12; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_13 = pipe2_io_vliw_out_13; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_14 = pipe2_io_vliw_out_14; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_15 = pipe2_io_vliw_out_15; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_16 = pipe2_io_vliw_out_16; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_17 = pipe2_io_vliw_out_17; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_18 = pipe2_io_vliw_out_18; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_19 = pipe2_io_vliw_out_19; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_20 = pipe2_io_vliw_out_20; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_21 = pipe2_io_vliw_out_21; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_22 = pipe2_io_vliw_out_22; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_23 = pipe2_io_vliw_out_23; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_24 = pipe2_io_vliw_out_24; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_25 = pipe2_io_vliw_out_25; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_26 = pipe2_io_vliw_out_26; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_27 = pipe2_io_vliw_out_27; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_28 = pipe2_io_vliw_out_28; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_29 = pipe2_io_vliw_out_29; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_30 = pipe2_io_vliw_out_30; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_31 = pipe2_io_vliw_out_31; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_32 = pipe2_io_vliw_out_32; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_33 = pipe2_io_vliw_out_33; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_34 = pipe2_io_vliw_out_34; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_35 = pipe2_io_vliw_out_35; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_36 = pipe2_io_vliw_out_36; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_37 = pipe2_io_vliw_out_37; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_38 = pipe2_io_vliw_out_38; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_39 = pipe2_io_vliw_out_39; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_40 = pipe2_io_vliw_out_40; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_41 = pipe2_io_vliw_out_41; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_42 = pipe2_io_vliw_out_42; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_43 = pipe2_io_vliw_out_43; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_44 = pipe2_io_vliw_out_44; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_45 = pipe2_io_vliw_out_45; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_46 = pipe2_io_vliw_out_46; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_47 = pipe2_io_vliw_out_47; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_48 = pipe2_io_vliw_out_48; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_49 = pipe2_io_vliw_out_49; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_50 = pipe2_io_vliw_out_50; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_51 = pipe2_io_vliw_out_51; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_52 = pipe2_io_vliw_out_52; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_53 = pipe2_io_vliw_out_53; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_54 = pipe2_io_vliw_out_54; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_55 = pipe2_io_vliw_out_55; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_56 = pipe2_io_vliw_out_56; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_57 = pipe2_io_vliw_out_57; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_58 = pipe2_io_vliw_out_58; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_59 = pipe2_io_vliw_out_59; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_60 = pipe2_io_vliw_out_60; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_61 = pipe2_io_vliw_out_61; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_62 = pipe2_io_vliw_out_62; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_63 = pipe2_io_vliw_out_63; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_64 = pipe2_io_vliw_out_64; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_65 = pipe2_io_vliw_out_65; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_66 = pipe2_io_vliw_out_66; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_67 = pipe2_io_vliw_out_67; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_68 = pipe2_io_vliw_out_68; // @[executor_pisa.scala 302:26]
  assign pipe3_io_vliw_in_69 = pipe2_io_vliw_out_69; // @[executor_pisa.scala 302:26]
  assign pipe3_io_nid_in = pipe2_io_nid_out; // @[executor_pisa.scala 303:26]
  assign pipe4_clock = clock;
  assign pipe4_io_pipe_phv_in_data_0 = pipe3_io_pipe_phv_out_data_0; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_1 = pipe3_io_pipe_phv_out_data_1; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_2 = pipe3_io_pipe_phv_out_data_2; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_3 = pipe3_io_pipe_phv_out_data_3; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_4 = pipe3_io_pipe_phv_out_data_4; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_5 = pipe3_io_pipe_phv_out_data_5; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_6 = pipe3_io_pipe_phv_out_data_6; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_7 = pipe3_io_pipe_phv_out_data_7; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_8 = pipe3_io_pipe_phv_out_data_8; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_9 = pipe3_io_pipe_phv_out_data_9; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_10 = pipe3_io_pipe_phv_out_data_10; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_11 = pipe3_io_pipe_phv_out_data_11; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_12 = pipe3_io_pipe_phv_out_data_12; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_13 = pipe3_io_pipe_phv_out_data_13; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_14 = pipe3_io_pipe_phv_out_data_14; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_15 = pipe3_io_pipe_phv_out_data_15; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_16 = pipe3_io_pipe_phv_out_data_16; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_17 = pipe3_io_pipe_phv_out_data_17; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_18 = pipe3_io_pipe_phv_out_data_18; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_19 = pipe3_io_pipe_phv_out_data_19; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_20 = pipe3_io_pipe_phv_out_data_20; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_21 = pipe3_io_pipe_phv_out_data_21; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_22 = pipe3_io_pipe_phv_out_data_22; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_23 = pipe3_io_pipe_phv_out_data_23; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_24 = pipe3_io_pipe_phv_out_data_24; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_25 = pipe3_io_pipe_phv_out_data_25; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_26 = pipe3_io_pipe_phv_out_data_26; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_27 = pipe3_io_pipe_phv_out_data_27; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_28 = pipe3_io_pipe_phv_out_data_28; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_29 = pipe3_io_pipe_phv_out_data_29; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_30 = pipe3_io_pipe_phv_out_data_30; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_31 = pipe3_io_pipe_phv_out_data_31; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_32 = pipe3_io_pipe_phv_out_data_32; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_33 = pipe3_io_pipe_phv_out_data_33; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_34 = pipe3_io_pipe_phv_out_data_34; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_35 = pipe3_io_pipe_phv_out_data_35; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_36 = pipe3_io_pipe_phv_out_data_36; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_37 = pipe3_io_pipe_phv_out_data_37; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_38 = pipe3_io_pipe_phv_out_data_38; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_39 = pipe3_io_pipe_phv_out_data_39; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_40 = pipe3_io_pipe_phv_out_data_40; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_41 = pipe3_io_pipe_phv_out_data_41; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_42 = pipe3_io_pipe_phv_out_data_42; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_43 = pipe3_io_pipe_phv_out_data_43; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_44 = pipe3_io_pipe_phv_out_data_44; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_45 = pipe3_io_pipe_phv_out_data_45; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_46 = pipe3_io_pipe_phv_out_data_46; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_47 = pipe3_io_pipe_phv_out_data_47; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_48 = pipe3_io_pipe_phv_out_data_48; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_49 = pipe3_io_pipe_phv_out_data_49; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_50 = pipe3_io_pipe_phv_out_data_50; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_51 = pipe3_io_pipe_phv_out_data_51; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_52 = pipe3_io_pipe_phv_out_data_52; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_53 = pipe3_io_pipe_phv_out_data_53; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_54 = pipe3_io_pipe_phv_out_data_54; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_55 = pipe3_io_pipe_phv_out_data_55; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_56 = pipe3_io_pipe_phv_out_data_56; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_57 = pipe3_io_pipe_phv_out_data_57; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_58 = pipe3_io_pipe_phv_out_data_58; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_59 = pipe3_io_pipe_phv_out_data_59; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_60 = pipe3_io_pipe_phv_out_data_60; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_61 = pipe3_io_pipe_phv_out_data_61; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_62 = pipe3_io_pipe_phv_out_data_62; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_63 = pipe3_io_pipe_phv_out_data_63; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_64 = pipe3_io_pipe_phv_out_data_64; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_65 = pipe3_io_pipe_phv_out_data_65; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_66 = pipe3_io_pipe_phv_out_data_66; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_67 = pipe3_io_pipe_phv_out_data_67; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_68 = pipe3_io_pipe_phv_out_data_68; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_69 = pipe3_io_pipe_phv_out_data_69; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_70 = pipe3_io_pipe_phv_out_data_70; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_71 = pipe3_io_pipe_phv_out_data_71; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_72 = pipe3_io_pipe_phv_out_data_72; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_73 = pipe3_io_pipe_phv_out_data_73; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_74 = pipe3_io_pipe_phv_out_data_74; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_75 = pipe3_io_pipe_phv_out_data_75; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_76 = pipe3_io_pipe_phv_out_data_76; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_77 = pipe3_io_pipe_phv_out_data_77; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_78 = pipe3_io_pipe_phv_out_data_78; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_79 = pipe3_io_pipe_phv_out_data_79; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_80 = pipe3_io_pipe_phv_out_data_80; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_81 = pipe3_io_pipe_phv_out_data_81; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_82 = pipe3_io_pipe_phv_out_data_82; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_83 = pipe3_io_pipe_phv_out_data_83; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_84 = pipe3_io_pipe_phv_out_data_84; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_85 = pipe3_io_pipe_phv_out_data_85; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_86 = pipe3_io_pipe_phv_out_data_86; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_87 = pipe3_io_pipe_phv_out_data_87; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_88 = pipe3_io_pipe_phv_out_data_88; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_89 = pipe3_io_pipe_phv_out_data_89; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_90 = pipe3_io_pipe_phv_out_data_90; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_91 = pipe3_io_pipe_phv_out_data_91; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_92 = pipe3_io_pipe_phv_out_data_92; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_93 = pipe3_io_pipe_phv_out_data_93; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_94 = pipe3_io_pipe_phv_out_data_94; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_95 = pipe3_io_pipe_phv_out_data_95; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_96 = pipe3_io_pipe_phv_out_data_96; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_97 = pipe3_io_pipe_phv_out_data_97; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_98 = pipe3_io_pipe_phv_out_data_98; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_99 = pipe3_io_pipe_phv_out_data_99; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_100 = pipe3_io_pipe_phv_out_data_100; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_101 = pipe3_io_pipe_phv_out_data_101; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_102 = pipe3_io_pipe_phv_out_data_102; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_103 = pipe3_io_pipe_phv_out_data_103; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_104 = pipe3_io_pipe_phv_out_data_104; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_105 = pipe3_io_pipe_phv_out_data_105; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_106 = pipe3_io_pipe_phv_out_data_106; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_107 = pipe3_io_pipe_phv_out_data_107; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_108 = pipe3_io_pipe_phv_out_data_108; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_109 = pipe3_io_pipe_phv_out_data_109; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_110 = pipe3_io_pipe_phv_out_data_110; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_111 = pipe3_io_pipe_phv_out_data_111; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_112 = pipe3_io_pipe_phv_out_data_112; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_113 = pipe3_io_pipe_phv_out_data_113; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_114 = pipe3_io_pipe_phv_out_data_114; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_115 = pipe3_io_pipe_phv_out_data_115; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_116 = pipe3_io_pipe_phv_out_data_116; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_117 = pipe3_io_pipe_phv_out_data_117; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_118 = pipe3_io_pipe_phv_out_data_118; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_119 = pipe3_io_pipe_phv_out_data_119; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_120 = pipe3_io_pipe_phv_out_data_120; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_121 = pipe3_io_pipe_phv_out_data_121; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_122 = pipe3_io_pipe_phv_out_data_122; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_123 = pipe3_io_pipe_phv_out_data_123; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_124 = pipe3_io_pipe_phv_out_data_124; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_125 = pipe3_io_pipe_phv_out_data_125; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_126 = pipe3_io_pipe_phv_out_data_126; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_127 = pipe3_io_pipe_phv_out_data_127; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_128 = pipe3_io_pipe_phv_out_data_128; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_129 = pipe3_io_pipe_phv_out_data_129; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_130 = pipe3_io_pipe_phv_out_data_130; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_131 = pipe3_io_pipe_phv_out_data_131; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_132 = pipe3_io_pipe_phv_out_data_132; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_133 = pipe3_io_pipe_phv_out_data_133; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_134 = pipe3_io_pipe_phv_out_data_134; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_135 = pipe3_io_pipe_phv_out_data_135; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_136 = pipe3_io_pipe_phv_out_data_136; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_137 = pipe3_io_pipe_phv_out_data_137; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_138 = pipe3_io_pipe_phv_out_data_138; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_139 = pipe3_io_pipe_phv_out_data_139; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_140 = pipe3_io_pipe_phv_out_data_140; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_141 = pipe3_io_pipe_phv_out_data_141; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_142 = pipe3_io_pipe_phv_out_data_142; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_143 = pipe3_io_pipe_phv_out_data_143; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_144 = pipe3_io_pipe_phv_out_data_144; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_145 = pipe3_io_pipe_phv_out_data_145; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_146 = pipe3_io_pipe_phv_out_data_146; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_147 = pipe3_io_pipe_phv_out_data_147; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_148 = pipe3_io_pipe_phv_out_data_148; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_149 = pipe3_io_pipe_phv_out_data_149; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_150 = pipe3_io_pipe_phv_out_data_150; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_151 = pipe3_io_pipe_phv_out_data_151; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_152 = pipe3_io_pipe_phv_out_data_152; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_153 = pipe3_io_pipe_phv_out_data_153; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_154 = pipe3_io_pipe_phv_out_data_154; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_155 = pipe3_io_pipe_phv_out_data_155; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_156 = pipe3_io_pipe_phv_out_data_156; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_157 = pipe3_io_pipe_phv_out_data_157; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_158 = pipe3_io_pipe_phv_out_data_158; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_data_159 = pipe3_io_pipe_phv_out_data_159; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_next_config_id = pipe3_io_pipe_phv_out_next_config_id; // @[executor_pisa.scala 305:26]
  assign pipe4_io_pipe_phv_in_is_valid_processor = pipe3_io_pipe_phv_out_is_valid_processor; // @[executor_pisa.scala 305:26]
  assign pipe4_io_nid_in = pipe3_io_nid_out; // @[executor_pisa.scala 306:26]
  assign pipe4_io_tag_in_0 = pipe3_io_tag_out_0; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_1 = pipe3_io_tag_out_1; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_2 = pipe3_io_tag_out_2; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_3 = pipe3_io_tag_out_3; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_4 = pipe3_io_tag_out_4; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_5 = pipe3_io_tag_out_5; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_6 = pipe3_io_tag_out_6; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_7 = pipe3_io_tag_out_7; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_8 = pipe3_io_tag_out_8; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_9 = pipe3_io_tag_out_9; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_10 = pipe3_io_tag_out_10; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_11 = pipe3_io_tag_out_11; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_12 = pipe3_io_tag_out_12; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_13 = pipe3_io_tag_out_13; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_14 = pipe3_io_tag_out_14; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_15 = pipe3_io_tag_out_15; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_16 = pipe3_io_tag_out_16; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_17 = pipe3_io_tag_out_17; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_18 = pipe3_io_tag_out_18; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_19 = pipe3_io_tag_out_19; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_20 = pipe3_io_tag_out_20; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_21 = pipe3_io_tag_out_21; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_22 = pipe3_io_tag_out_22; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_23 = pipe3_io_tag_out_23; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_24 = pipe3_io_tag_out_24; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_25 = pipe3_io_tag_out_25; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_26 = pipe3_io_tag_out_26; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_27 = pipe3_io_tag_out_27; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_28 = pipe3_io_tag_out_28; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_29 = pipe3_io_tag_out_29; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_30 = pipe3_io_tag_out_30; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_31 = pipe3_io_tag_out_31; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_32 = pipe3_io_tag_out_32; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_33 = pipe3_io_tag_out_33; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_34 = pipe3_io_tag_out_34; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_35 = pipe3_io_tag_out_35; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_36 = pipe3_io_tag_out_36; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_37 = pipe3_io_tag_out_37; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_38 = pipe3_io_tag_out_38; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_39 = pipe3_io_tag_out_39; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_40 = pipe3_io_tag_out_40; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_41 = pipe3_io_tag_out_41; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_42 = pipe3_io_tag_out_42; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_43 = pipe3_io_tag_out_43; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_44 = pipe3_io_tag_out_44; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_45 = pipe3_io_tag_out_45; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_46 = pipe3_io_tag_out_46; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_47 = pipe3_io_tag_out_47; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_48 = pipe3_io_tag_out_48; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_49 = pipe3_io_tag_out_49; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_50 = pipe3_io_tag_out_50; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_51 = pipe3_io_tag_out_51; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_52 = pipe3_io_tag_out_52; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_53 = pipe3_io_tag_out_53; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_54 = pipe3_io_tag_out_54; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_55 = pipe3_io_tag_out_55; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_56 = pipe3_io_tag_out_56; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_57 = pipe3_io_tag_out_57; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_58 = pipe3_io_tag_out_58; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_59 = pipe3_io_tag_out_59; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_60 = pipe3_io_tag_out_60; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_61 = pipe3_io_tag_out_61; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_62 = pipe3_io_tag_out_62; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_63 = pipe3_io_tag_out_63; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_64 = pipe3_io_tag_out_64; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_65 = pipe3_io_tag_out_65; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_66 = pipe3_io_tag_out_66; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_67 = pipe3_io_tag_out_67; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_68 = pipe3_io_tag_out_68; // @[executor_pisa.scala 307:26]
  assign pipe4_io_tag_in_69 = pipe3_io_tag_out_69; // @[executor_pisa.scala 307:26]
  assign pipe4_io_field_set_field8_0 = pipe3_io_field_set_field8_0; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field8_1 = pipe3_io_field_set_field8_1; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field8_2 = pipe3_io_field_set_field8_2; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field8_3 = pipe3_io_field_set_field8_3; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field8_4 = pipe3_io_field_set_field8_4; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field8_5 = pipe3_io_field_set_field8_5; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field8_6 = pipe3_io_field_set_field8_6; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field8_7 = pipe3_io_field_set_field8_7; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field8_8 = pipe3_io_field_set_field8_8; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field8_9 = pipe3_io_field_set_field8_9; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field8_10 = pipe3_io_field_set_field8_10; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field8_11 = pipe3_io_field_set_field8_11; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field8_12 = pipe3_io_field_set_field8_12; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field8_13 = pipe3_io_field_set_field8_13; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field8_14 = pipe3_io_field_set_field8_14; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field8_15 = pipe3_io_field_set_field8_15; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field8_16 = pipe3_io_field_set_field8_16; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field8_17 = pipe3_io_field_set_field8_17; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field8_18 = pipe3_io_field_set_field8_18; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field8_19 = pipe3_io_field_set_field8_19; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_0 = pipe3_io_field_set_field16_0; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_1 = pipe3_io_field_set_field16_1; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_2 = pipe3_io_field_set_field16_2; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_3 = pipe3_io_field_set_field16_3; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_4 = pipe3_io_field_set_field16_4; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_5 = pipe3_io_field_set_field16_5; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_6 = pipe3_io_field_set_field16_6; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_7 = pipe3_io_field_set_field16_7; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_8 = pipe3_io_field_set_field16_8; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_9 = pipe3_io_field_set_field16_9; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_10 = pipe3_io_field_set_field16_10; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_11 = pipe3_io_field_set_field16_11; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_12 = pipe3_io_field_set_field16_12; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_13 = pipe3_io_field_set_field16_13; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_14 = pipe3_io_field_set_field16_14; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_15 = pipe3_io_field_set_field16_15; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_16 = pipe3_io_field_set_field16_16; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_17 = pipe3_io_field_set_field16_17; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_18 = pipe3_io_field_set_field16_18; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_19 = pipe3_io_field_set_field16_19; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_20 = pipe3_io_field_set_field16_20; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_21 = pipe3_io_field_set_field16_21; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_22 = pipe3_io_field_set_field16_22; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_23 = pipe3_io_field_set_field16_23; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_24 = pipe3_io_field_set_field16_24; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_25 = pipe3_io_field_set_field16_25; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_26 = pipe3_io_field_set_field16_26; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_27 = pipe3_io_field_set_field16_27; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_28 = pipe3_io_field_set_field16_28; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field16_29 = pipe3_io_field_set_field16_29; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field32_0 = pipe3_io_field_set_field32_0; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field32_1 = pipe3_io_field_set_field32_1; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field32_2 = pipe3_io_field_set_field32_2; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field32_3 = pipe3_io_field_set_field32_3; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field32_4 = pipe3_io_field_set_field32_4; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field32_5 = pipe3_io_field_set_field32_5; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field32_6 = pipe3_io_field_set_field32_6; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field32_7 = pipe3_io_field_set_field32_7; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field32_8 = pipe3_io_field_set_field32_8; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field32_9 = pipe3_io_field_set_field32_9; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field32_10 = pipe3_io_field_set_field32_10; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field32_11 = pipe3_io_field_set_field32_11; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field32_12 = pipe3_io_field_set_field32_12; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field32_13 = pipe3_io_field_set_field32_13; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field32_14 = pipe3_io_field_set_field32_14; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field32_15 = pipe3_io_field_set_field32_15; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field32_16 = pipe3_io_field_set_field32_16; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field32_17 = pipe3_io_field_set_field32_17; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field32_18 = pipe3_io_field_set_field32_18; // @[executor_pisa.scala 308:26]
  assign pipe4_io_field_set_field32_19 = pipe3_io_field_set_field32_19; // @[executor_pisa.scala 308:26]
endmodule
