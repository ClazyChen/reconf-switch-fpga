module InPort(
  input           io_en,
  input  [1023:0] io_data,
  output [7:0]    io_phv_out_data_0,
  output [7:0]    io_phv_out_data_1,
  output [7:0]    io_phv_out_data_2,
  output [7:0]    io_phv_out_data_3,
  output [7:0]    io_phv_out_data_4,
  output [7:0]    io_phv_out_data_5,
  output [7:0]    io_phv_out_data_6,
  output [7:0]    io_phv_out_data_7,
  output [7:0]    io_phv_out_data_8,
  output [7:0]    io_phv_out_data_9,
  output [7:0]    io_phv_out_data_10,
  output [7:0]    io_phv_out_data_11,
  output [7:0]    io_phv_out_data_12,
  output [7:0]    io_phv_out_data_13,
  output [7:0]    io_phv_out_data_14,
  output [7:0]    io_phv_out_data_15,
  output [7:0]    io_phv_out_data_16,
  output [7:0]    io_phv_out_data_17,
  output [7:0]    io_phv_out_data_18,
  output [7:0]    io_phv_out_data_19,
  output [7:0]    io_phv_out_data_20,
  output [7:0]    io_phv_out_data_21,
  output [7:0]    io_phv_out_data_22,
  output [7:0]    io_phv_out_data_23,
  output [7:0]    io_phv_out_data_24,
  output [7:0]    io_phv_out_data_25,
  output [7:0]    io_phv_out_data_26,
  output [7:0]    io_phv_out_data_27,
  output [7:0]    io_phv_out_data_28,
  output [7:0]    io_phv_out_data_29,
  output [7:0]    io_phv_out_data_30,
  output [7:0]    io_phv_out_data_31,
  output [7:0]    io_phv_out_data_32,
  output [7:0]    io_phv_out_data_33,
  output [7:0]    io_phv_out_data_34,
  output [7:0]    io_phv_out_data_35,
  output [7:0]    io_phv_out_data_36,
  output [7:0]    io_phv_out_data_37,
  output [7:0]    io_phv_out_data_38,
  output [7:0]    io_phv_out_data_39,
  output [7:0]    io_phv_out_data_40,
  output [7:0]    io_phv_out_data_41,
  output [7:0]    io_phv_out_data_42,
  output [7:0]    io_phv_out_data_43,
  output [7:0]    io_phv_out_data_44,
  output [7:0]    io_phv_out_data_45,
  output [7:0]    io_phv_out_data_46,
  output [7:0]    io_phv_out_data_47,
  output [7:0]    io_phv_out_data_48,
  output [7:0]    io_phv_out_data_49,
  output [7:0]    io_phv_out_data_50,
  output [7:0]    io_phv_out_data_51,
  output [7:0]    io_phv_out_data_52,
  output [7:0]    io_phv_out_data_53,
  output [7:0]    io_phv_out_data_54,
  output [7:0]    io_phv_out_data_55,
  output [7:0]    io_phv_out_data_56,
  output [7:0]    io_phv_out_data_57,
  output [7:0]    io_phv_out_data_58,
  output [7:0]    io_phv_out_data_59,
  output [7:0]    io_phv_out_data_60,
  output [7:0]    io_phv_out_data_61,
  output [7:0]    io_phv_out_data_62,
  output [7:0]    io_phv_out_data_63,
  output [7:0]    io_phv_out_data_64,
  output [7:0]    io_phv_out_data_65,
  output [7:0]    io_phv_out_data_66,
  output [7:0]    io_phv_out_data_67,
  output [7:0]    io_phv_out_data_68,
  output [7:0]    io_phv_out_data_69,
  output [7:0]    io_phv_out_data_70,
  output [7:0]    io_phv_out_data_71,
  output [7:0]    io_phv_out_data_72,
  output [7:0]    io_phv_out_data_73,
  output [7:0]    io_phv_out_data_74,
  output [7:0]    io_phv_out_data_75,
  output [7:0]    io_phv_out_data_76,
  output [7:0]    io_phv_out_data_77,
  output [7:0]    io_phv_out_data_78,
  output [7:0]    io_phv_out_data_79,
  output [7:0]    io_phv_out_data_80,
  output [7:0]    io_phv_out_data_81,
  output [7:0]    io_phv_out_data_82,
  output [7:0]    io_phv_out_data_83,
  output [7:0]    io_phv_out_data_84,
  output [7:0]    io_phv_out_data_85,
  output [7:0]    io_phv_out_data_86,
  output [7:0]    io_phv_out_data_87,
  output [7:0]    io_phv_out_data_88,
  output [7:0]    io_phv_out_data_89,
  output [7:0]    io_phv_out_data_90,
  output [7:0]    io_phv_out_data_91,
  output [7:0]    io_phv_out_data_92,
  output [7:0]    io_phv_out_data_93,
  output [7:0]    io_phv_out_data_94,
  output [7:0]    io_phv_out_data_95,
  output [7:0]    io_phv_out_data_96,
  output [7:0]    io_phv_out_data_97,
  output [7:0]    io_phv_out_data_98,
  output [7:0]    io_phv_out_data_99,
  output [7:0]    io_phv_out_data_100,
  output [7:0]    io_phv_out_data_101,
  output [7:0]    io_phv_out_data_102,
  output [7:0]    io_phv_out_data_103,
  output [7:0]    io_phv_out_data_104,
  output [7:0]    io_phv_out_data_105,
  output [7:0]    io_phv_out_data_106,
  output [7:0]    io_phv_out_data_107,
  output [7:0]    io_phv_out_data_108,
  output [7:0]    io_phv_out_data_109,
  output [7:0]    io_phv_out_data_110,
  output [7:0]    io_phv_out_data_111,
  output [7:0]    io_phv_out_data_112,
  output [7:0]    io_phv_out_data_113,
  output [7:0]    io_phv_out_data_114,
  output [7:0]    io_phv_out_data_115,
  output [7:0]    io_phv_out_data_116,
  output [7:0]    io_phv_out_data_117,
  output [7:0]    io_phv_out_data_118,
  output [7:0]    io_phv_out_data_119,
  output [7:0]    io_phv_out_data_120,
  output [7:0]    io_phv_out_data_121,
  output [7:0]    io_phv_out_data_122,
  output [7:0]    io_phv_out_data_123,
  output [7:0]    io_phv_out_data_124,
  output [7:0]    io_phv_out_data_125,
  output [7:0]    io_phv_out_data_126,
  output [7:0]    io_phv_out_data_127,
  output          io_phv_out_valid
);
  assign io_phv_out_data_0 = io_data[1023:1016]; // @[inport.scala 14:38]
  assign io_phv_out_data_1 = io_data[1015:1008]; // @[inport.scala 14:38]
  assign io_phv_out_data_2 = io_data[1007:1000]; // @[inport.scala 14:38]
  assign io_phv_out_data_3 = io_data[999:992]; // @[inport.scala 14:38]
  assign io_phv_out_data_4 = io_data[991:984]; // @[inport.scala 14:38]
  assign io_phv_out_data_5 = io_data[983:976]; // @[inport.scala 14:38]
  assign io_phv_out_data_6 = io_data[975:968]; // @[inport.scala 14:38]
  assign io_phv_out_data_7 = io_data[967:960]; // @[inport.scala 14:38]
  assign io_phv_out_data_8 = io_data[959:952]; // @[inport.scala 14:38]
  assign io_phv_out_data_9 = io_data[951:944]; // @[inport.scala 14:38]
  assign io_phv_out_data_10 = io_data[943:936]; // @[inport.scala 14:38]
  assign io_phv_out_data_11 = io_data[935:928]; // @[inport.scala 14:38]
  assign io_phv_out_data_12 = io_data[927:920]; // @[inport.scala 14:38]
  assign io_phv_out_data_13 = io_data[919:912]; // @[inport.scala 14:38]
  assign io_phv_out_data_14 = io_data[911:904]; // @[inport.scala 14:38]
  assign io_phv_out_data_15 = io_data[903:896]; // @[inport.scala 14:38]
  assign io_phv_out_data_16 = io_data[895:888]; // @[inport.scala 14:38]
  assign io_phv_out_data_17 = io_data[887:880]; // @[inport.scala 14:38]
  assign io_phv_out_data_18 = io_data[879:872]; // @[inport.scala 14:38]
  assign io_phv_out_data_19 = io_data[871:864]; // @[inport.scala 14:38]
  assign io_phv_out_data_20 = io_data[863:856]; // @[inport.scala 14:38]
  assign io_phv_out_data_21 = io_data[855:848]; // @[inport.scala 14:38]
  assign io_phv_out_data_22 = io_data[847:840]; // @[inport.scala 14:38]
  assign io_phv_out_data_23 = io_data[839:832]; // @[inport.scala 14:38]
  assign io_phv_out_data_24 = io_data[831:824]; // @[inport.scala 14:38]
  assign io_phv_out_data_25 = io_data[823:816]; // @[inport.scala 14:38]
  assign io_phv_out_data_26 = io_data[815:808]; // @[inport.scala 14:38]
  assign io_phv_out_data_27 = io_data[807:800]; // @[inport.scala 14:38]
  assign io_phv_out_data_28 = io_data[799:792]; // @[inport.scala 14:38]
  assign io_phv_out_data_29 = io_data[791:784]; // @[inport.scala 14:38]
  assign io_phv_out_data_30 = io_data[783:776]; // @[inport.scala 14:38]
  assign io_phv_out_data_31 = io_data[775:768]; // @[inport.scala 14:38]
  assign io_phv_out_data_32 = io_data[767:760]; // @[inport.scala 14:38]
  assign io_phv_out_data_33 = io_data[759:752]; // @[inport.scala 14:38]
  assign io_phv_out_data_34 = io_data[751:744]; // @[inport.scala 14:38]
  assign io_phv_out_data_35 = io_data[743:736]; // @[inport.scala 14:38]
  assign io_phv_out_data_36 = io_data[735:728]; // @[inport.scala 14:38]
  assign io_phv_out_data_37 = io_data[727:720]; // @[inport.scala 14:38]
  assign io_phv_out_data_38 = io_data[719:712]; // @[inport.scala 14:38]
  assign io_phv_out_data_39 = io_data[711:704]; // @[inport.scala 14:38]
  assign io_phv_out_data_40 = io_data[703:696]; // @[inport.scala 14:38]
  assign io_phv_out_data_41 = io_data[695:688]; // @[inport.scala 14:38]
  assign io_phv_out_data_42 = io_data[687:680]; // @[inport.scala 14:38]
  assign io_phv_out_data_43 = io_data[679:672]; // @[inport.scala 14:38]
  assign io_phv_out_data_44 = io_data[671:664]; // @[inport.scala 14:38]
  assign io_phv_out_data_45 = io_data[663:656]; // @[inport.scala 14:38]
  assign io_phv_out_data_46 = io_data[655:648]; // @[inport.scala 14:38]
  assign io_phv_out_data_47 = io_data[647:640]; // @[inport.scala 14:38]
  assign io_phv_out_data_48 = io_data[639:632]; // @[inport.scala 14:38]
  assign io_phv_out_data_49 = io_data[631:624]; // @[inport.scala 14:38]
  assign io_phv_out_data_50 = io_data[623:616]; // @[inport.scala 14:38]
  assign io_phv_out_data_51 = io_data[615:608]; // @[inport.scala 14:38]
  assign io_phv_out_data_52 = io_data[607:600]; // @[inport.scala 14:38]
  assign io_phv_out_data_53 = io_data[599:592]; // @[inport.scala 14:38]
  assign io_phv_out_data_54 = io_data[591:584]; // @[inport.scala 14:38]
  assign io_phv_out_data_55 = io_data[583:576]; // @[inport.scala 14:38]
  assign io_phv_out_data_56 = io_data[575:568]; // @[inport.scala 14:38]
  assign io_phv_out_data_57 = io_data[567:560]; // @[inport.scala 14:38]
  assign io_phv_out_data_58 = io_data[559:552]; // @[inport.scala 14:38]
  assign io_phv_out_data_59 = io_data[551:544]; // @[inport.scala 14:38]
  assign io_phv_out_data_60 = io_data[543:536]; // @[inport.scala 14:38]
  assign io_phv_out_data_61 = io_data[535:528]; // @[inport.scala 14:38]
  assign io_phv_out_data_62 = io_data[527:520]; // @[inport.scala 14:38]
  assign io_phv_out_data_63 = io_data[519:512]; // @[inport.scala 14:38]
  assign io_phv_out_data_64 = io_data[511:504]; // @[inport.scala 14:38]
  assign io_phv_out_data_65 = io_data[503:496]; // @[inport.scala 14:38]
  assign io_phv_out_data_66 = io_data[495:488]; // @[inport.scala 14:38]
  assign io_phv_out_data_67 = io_data[487:480]; // @[inport.scala 14:38]
  assign io_phv_out_data_68 = io_data[479:472]; // @[inport.scala 14:38]
  assign io_phv_out_data_69 = io_data[471:464]; // @[inport.scala 14:38]
  assign io_phv_out_data_70 = io_data[463:456]; // @[inport.scala 14:38]
  assign io_phv_out_data_71 = io_data[455:448]; // @[inport.scala 14:38]
  assign io_phv_out_data_72 = io_data[447:440]; // @[inport.scala 14:38]
  assign io_phv_out_data_73 = io_data[439:432]; // @[inport.scala 14:38]
  assign io_phv_out_data_74 = io_data[431:424]; // @[inport.scala 14:38]
  assign io_phv_out_data_75 = io_data[423:416]; // @[inport.scala 14:38]
  assign io_phv_out_data_76 = io_data[415:408]; // @[inport.scala 14:38]
  assign io_phv_out_data_77 = io_data[407:400]; // @[inport.scala 14:38]
  assign io_phv_out_data_78 = io_data[399:392]; // @[inport.scala 14:38]
  assign io_phv_out_data_79 = io_data[391:384]; // @[inport.scala 14:38]
  assign io_phv_out_data_80 = io_data[383:376]; // @[inport.scala 14:38]
  assign io_phv_out_data_81 = io_data[375:368]; // @[inport.scala 14:38]
  assign io_phv_out_data_82 = io_data[367:360]; // @[inport.scala 14:38]
  assign io_phv_out_data_83 = io_data[359:352]; // @[inport.scala 14:38]
  assign io_phv_out_data_84 = io_data[351:344]; // @[inport.scala 14:38]
  assign io_phv_out_data_85 = io_data[343:336]; // @[inport.scala 14:38]
  assign io_phv_out_data_86 = io_data[335:328]; // @[inport.scala 14:38]
  assign io_phv_out_data_87 = io_data[327:320]; // @[inport.scala 14:38]
  assign io_phv_out_data_88 = io_data[319:312]; // @[inport.scala 14:38]
  assign io_phv_out_data_89 = io_data[311:304]; // @[inport.scala 14:38]
  assign io_phv_out_data_90 = io_data[303:296]; // @[inport.scala 14:38]
  assign io_phv_out_data_91 = io_data[295:288]; // @[inport.scala 14:38]
  assign io_phv_out_data_92 = io_data[287:280]; // @[inport.scala 14:38]
  assign io_phv_out_data_93 = io_data[279:272]; // @[inport.scala 14:38]
  assign io_phv_out_data_94 = io_data[271:264]; // @[inport.scala 14:38]
  assign io_phv_out_data_95 = io_data[263:256]; // @[inport.scala 14:38]
  assign io_phv_out_data_96 = io_data[255:248]; // @[inport.scala 14:38]
  assign io_phv_out_data_97 = io_data[247:240]; // @[inport.scala 14:38]
  assign io_phv_out_data_98 = io_data[239:232]; // @[inport.scala 14:38]
  assign io_phv_out_data_99 = io_data[231:224]; // @[inport.scala 14:38]
  assign io_phv_out_data_100 = io_data[223:216]; // @[inport.scala 14:38]
  assign io_phv_out_data_101 = io_data[215:208]; // @[inport.scala 14:38]
  assign io_phv_out_data_102 = io_data[207:200]; // @[inport.scala 14:38]
  assign io_phv_out_data_103 = io_data[199:192]; // @[inport.scala 14:38]
  assign io_phv_out_data_104 = io_data[191:184]; // @[inport.scala 14:38]
  assign io_phv_out_data_105 = io_data[183:176]; // @[inport.scala 14:38]
  assign io_phv_out_data_106 = io_data[175:168]; // @[inport.scala 14:38]
  assign io_phv_out_data_107 = io_data[167:160]; // @[inport.scala 14:38]
  assign io_phv_out_data_108 = io_data[159:152]; // @[inport.scala 14:38]
  assign io_phv_out_data_109 = io_data[151:144]; // @[inport.scala 14:38]
  assign io_phv_out_data_110 = io_data[143:136]; // @[inport.scala 14:38]
  assign io_phv_out_data_111 = io_data[135:128]; // @[inport.scala 14:38]
  assign io_phv_out_data_112 = io_data[127:120]; // @[inport.scala 14:38]
  assign io_phv_out_data_113 = io_data[119:112]; // @[inport.scala 14:38]
  assign io_phv_out_data_114 = io_data[111:104]; // @[inport.scala 14:38]
  assign io_phv_out_data_115 = io_data[103:96]; // @[inport.scala 14:38]
  assign io_phv_out_data_116 = io_data[95:88]; // @[inport.scala 14:38]
  assign io_phv_out_data_117 = io_data[87:80]; // @[inport.scala 14:38]
  assign io_phv_out_data_118 = io_data[79:72]; // @[inport.scala 14:38]
  assign io_phv_out_data_119 = io_data[71:64]; // @[inport.scala 14:38]
  assign io_phv_out_data_120 = io_data[63:56]; // @[inport.scala 14:38]
  assign io_phv_out_data_121 = io_data[55:48]; // @[inport.scala 14:38]
  assign io_phv_out_data_122 = io_data[47:40]; // @[inport.scala 14:38]
  assign io_phv_out_data_123 = io_data[39:32]; // @[inport.scala 14:38]
  assign io_phv_out_data_124 = io_data[31:24]; // @[inport.scala 14:38]
  assign io_phv_out_data_125 = io_data[23:16]; // @[inport.scala 14:38]
  assign io_phv_out_data_126 = io_data[15:8]; // @[inport.scala 14:38]
  assign io_phv_out_data_127 = io_data[7:0]; // @[inport.scala 14:38]
  assign io_phv_out_valid = io_en; // @[inport.scala 31:39]
endmodule
