module OutPort(
  input         clock,
  input  [7:0]  io_phv_in_data_0,
  input  [7:0]  io_phv_in_data_1,
  input  [7:0]  io_phv_in_data_2,
  input  [7:0]  io_phv_in_data_3,
  input  [7:0]  io_phv_in_data_4,
  input  [7:0]  io_phv_in_data_5,
  input  [7:0]  io_phv_in_data_6,
  input  [7:0]  io_phv_in_data_7,
  input  [7:0]  io_phv_in_data_8,
  input  [7:0]  io_phv_in_data_9,
  input  [7:0]  io_phv_in_data_10,
  input  [7:0]  io_phv_in_data_11,
  input  [7:0]  io_phv_in_data_12,
  input  [7:0]  io_phv_in_data_13,
  input  [7:0]  io_phv_in_data_14,
  input  [7:0]  io_phv_in_data_15,
  input  [7:0]  io_phv_in_data_16,
  input  [7:0]  io_phv_in_data_17,
  input  [7:0]  io_phv_in_data_18,
  input  [7:0]  io_phv_in_data_19,
  input  [7:0]  io_phv_in_data_20,
  input  [7:0]  io_phv_in_data_21,
  input  [7:0]  io_phv_in_data_22,
  input  [7:0]  io_phv_in_data_23,
  input  [7:0]  io_phv_in_data_24,
  input  [7:0]  io_phv_in_data_25,
  input  [7:0]  io_phv_in_data_26,
  input  [7:0]  io_phv_in_data_27,
  input  [7:0]  io_phv_in_data_28,
  input  [7:0]  io_phv_in_data_29,
  input  [7:0]  io_phv_in_data_30,
  input  [7:0]  io_phv_in_data_31,
  input  [7:0]  io_phv_in_data_32,
  input  [7:0]  io_phv_in_data_33,
  input  [7:0]  io_phv_in_data_34,
  input  [7:0]  io_phv_in_data_35,
  input  [7:0]  io_phv_in_data_36,
  input  [7:0]  io_phv_in_data_37,
  input  [7:0]  io_phv_in_data_38,
  input  [7:0]  io_phv_in_data_39,
  input  [7:0]  io_phv_in_data_40,
  input  [7:0]  io_phv_in_data_41,
  input  [7:0]  io_phv_in_data_42,
  input  [7:0]  io_phv_in_data_43,
  input  [7:0]  io_phv_in_data_44,
  input  [7:0]  io_phv_in_data_45,
  input  [7:0]  io_phv_in_data_46,
  input  [7:0]  io_phv_in_data_47,
  input  [7:0]  io_phv_in_data_48,
  input  [7:0]  io_phv_in_data_49,
  input  [7:0]  io_phv_in_data_50,
  input  [7:0]  io_phv_in_data_51,
  input  [7:0]  io_phv_in_data_52,
  input  [7:0]  io_phv_in_data_53,
  input  [7:0]  io_phv_in_data_54,
  input  [7:0]  io_phv_in_data_55,
  input  [7:0]  io_phv_in_data_56,
  input  [7:0]  io_phv_in_data_57,
  input  [7:0]  io_phv_in_data_58,
  input  [7:0]  io_phv_in_data_59,
  input  [7:0]  io_phv_in_data_60,
  input  [7:0]  io_phv_in_data_61,
  input  [7:0]  io_phv_in_data_62,
  input  [7:0]  io_phv_in_data_63,
  input  [7:0]  io_phv_in_data_64,
  input  [7:0]  io_phv_in_data_65,
  input  [7:0]  io_phv_in_data_66,
  input  [7:0]  io_phv_in_data_67,
  input  [7:0]  io_phv_in_data_68,
  input  [7:0]  io_phv_in_data_69,
  input  [7:0]  io_phv_in_data_70,
  input  [7:0]  io_phv_in_data_71,
  input  [7:0]  io_phv_in_data_72,
  input  [7:0]  io_phv_in_data_73,
  input  [7:0]  io_phv_in_data_74,
  input  [7:0]  io_phv_in_data_75,
  input  [7:0]  io_phv_in_data_76,
  input  [7:0]  io_phv_in_data_77,
  input  [7:0]  io_phv_in_data_78,
  input  [7:0]  io_phv_in_data_79,
  input  [7:0]  io_phv_in_data_80,
  input  [7:0]  io_phv_in_data_81,
  input  [7:0]  io_phv_in_data_82,
  input  [7:0]  io_phv_in_data_83,
  input  [7:0]  io_phv_in_data_84,
  input  [7:0]  io_phv_in_data_85,
  input  [7:0]  io_phv_in_data_86,
  input  [7:0]  io_phv_in_data_87,
  input  [7:0]  io_phv_in_data_88,
  input  [7:0]  io_phv_in_data_89,
  input  [7:0]  io_phv_in_data_90,
  input  [7:0]  io_phv_in_data_91,
  input  [7:0]  io_phv_in_data_92,
  input  [7:0]  io_phv_in_data_93,
  input  [7:0]  io_phv_in_data_94,
  input  [7:0]  io_phv_in_data_95,
  input  [7:0]  io_phv_in_data_96,
  input  [7:0]  io_phv_in_data_97,
  input  [7:0]  io_phv_in_data_98,
  input  [7:0]  io_phv_in_data_99,
  input  [7:0]  io_phv_in_data_100,
  input  [7:0]  io_phv_in_data_101,
  input  [7:0]  io_phv_in_data_102,
  input  [7:0]  io_phv_in_data_103,
  input  [7:0]  io_phv_in_data_104,
  input  [7:0]  io_phv_in_data_105,
  input  [7:0]  io_phv_in_data_106,
  input  [7:0]  io_phv_in_data_107,
  input  [7:0]  io_phv_in_data_108,
  input  [7:0]  io_phv_in_data_109,
  input  [7:0]  io_phv_in_data_110,
  input  [7:0]  io_phv_in_data_111,
  input  [7:0]  io_phv_in_data_112,
  input  [7:0]  io_phv_in_data_113,
  input  [7:0]  io_phv_in_data_114,
  input  [7:0]  io_phv_in_data_115,
  input  [7:0]  io_phv_in_data_116,
  input  [7:0]  io_phv_in_data_117,
  input  [7:0]  io_phv_in_data_118,
  input  [7:0]  io_phv_in_data_119,
  input  [7:0]  io_phv_in_data_120,
  input  [7:0]  io_phv_in_data_121,
  input  [7:0]  io_phv_in_data_122,
  input  [7:0]  io_phv_in_data_123,
  input  [7:0]  io_phv_in_data_124,
  input  [7:0]  io_phv_in_data_125,
  input  [7:0]  io_phv_in_data_126,
  input  [7:0]  io_phv_in_data_127,
  input  [7:0]  io_phv_in_data_128,
  input  [7:0]  io_phv_in_data_129,
  input  [7:0]  io_phv_in_data_130,
  input  [7:0]  io_phv_in_data_131,
  input  [7:0]  io_phv_in_data_132,
  input  [7:0]  io_phv_in_data_133,
  input  [7:0]  io_phv_in_data_134,
  input  [7:0]  io_phv_in_data_135,
  input  [7:0]  io_phv_in_data_136,
  input  [7:0]  io_phv_in_data_137,
  input  [7:0]  io_phv_in_data_138,
  input  [7:0]  io_phv_in_data_139,
  input  [7:0]  io_phv_in_data_140,
  input  [7:0]  io_phv_in_data_141,
  input  [7:0]  io_phv_in_data_142,
  input  [7:0]  io_phv_in_data_143,
  input  [7:0]  io_phv_in_data_144,
  input  [7:0]  io_phv_in_data_145,
  input  [7:0]  io_phv_in_data_146,
  input  [7:0]  io_phv_in_data_147,
  input  [7:0]  io_phv_in_data_148,
  input  [7:0]  io_phv_in_data_149,
  input  [7:0]  io_phv_in_data_150,
  input  [7:0]  io_phv_in_data_151,
  input  [7:0]  io_phv_in_data_152,
  input  [7:0]  io_phv_in_data_153,
  input  [7:0]  io_phv_in_data_154,
  input  [7:0]  io_phv_in_data_155,
  input  [7:0]  io_phv_in_data_156,
  input  [7:0]  io_phv_in_data_157,
  input  [7:0]  io_phv_in_data_158,
  input  [7:0]  io_phv_in_data_159,
  input  [7:0]  io_phv_in_data_160,
  input  [7:0]  io_phv_in_data_161,
  input  [7:0]  io_phv_in_data_162,
  input  [7:0]  io_phv_in_data_163,
  input  [7:0]  io_phv_in_data_164,
  input  [7:0]  io_phv_in_data_165,
  input  [7:0]  io_phv_in_data_166,
  input  [7:0]  io_phv_in_data_167,
  input  [7:0]  io_phv_in_data_168,
  input  [7:0]  io_phv_in_data_169,
  input  [7:0]  io_phv_in_data_170,
  input  [7:0]  io_phv_in_data_171,
  input  [7:0]  io_phv_in_data_172,
  input  [7:0]  io_phv_in_data_173,
  input  [7:0]  io_phv_in_data_174,
  input  [7:0]  io_phv_in_data_175,
  input  [7:0]  io_phv_in_data_176,
  input  [7:0]  io_phv_in_data_177,
  input  [7:0]  io_phv_in_data_178,
  input  [7:0]  io_phv_in_data_179,
  input  [7:0]  io_phv_in_data_180,
  input  [7:0]  io_phv_in_data_181,
  input  [7:0]  io_phv_in_data_182,
  input  [7:0]  io_phv_in_data_183,
  input  [7:0]  io_phv_in_data_184,
  input  [7:0]  io_phv_in_data_185,
  input  [7:0]  io_phv_in_data_186,
  input  [7:0]  io_phv_in_data_187,
  input  [7:0]  io_phv_in_data_188,
  input  [7:0]  io_phv_in_data_189,
  input  [7:0]  io_phv_in_data_190,
  input  [7:0]  io_phv_in_data_191,
  input  [7:0]  io_phv_in_data_192,
  input  [7:0]  io_phv_in_data_193,
  input  [7:0]  io_phv_in_data_194,
  input  [7:0]  io_phv_in_data_195,
  input  [7:0]  io_phv_in_data_196,
  input  [7:0]  io_phv_in_data_197,
  input  [7:0]  io_phv_in_data_198,
  input  [7:0]  io_phv_in_data_199,
  input  [7:0]  io_phv_in_data_200,
  input  [7:0]  io_phv_in_data_201,
  input  [7:0]  io_phv_in_data_202,
  input  [7:0]  io_phv_in_data_203,
  input  [7:0]  io_phv_in_data_204,
  input  [7:0]  io_phv_in_data_205,
  input  [7:0]  io_phv_in_data_206,
  input  [7:0]  io_phv_in_data_207,
  input  [7:0]  io_phv_in_data_208,
  input  [7:0]  io_phv_in_data_209,
  input  [7:0]  io_phv_in_data_210,
  input  [7:0]  io_phv_in_data_211,
  input  [7:0]  io_phv_in_data_212,
  input  [7:0]  io_phv_in_data_213,
  input  [7:0]  io_phv_in_data_214,
  input  [7:0]  io_phv_in_data_215,
  input  [7:0]  io_phv_in_data_216,
  input  [7:0]  io_phv_in_data_217,
  input  [7:0]  io_phv_in_data_218,
  input  [7:0]  io_phv_in_data_219,
  input  [7:0]  io_phv_in_data_220,
  input  [7:0]  io_phv_in_data_221,
  input  [7:0]  io_phv_in_data_222,
  input  [7:0]  io_phv_in_data_223,
  input  [7:0]  io_phv_in_data_224,
  input  [7:0]  io_phv_in_data_225,
  input  [7:0]  io_phv_in_data_226,
  input  [7:0]  io_phv_in_data_227,
  input  [7:0]  io_phv_in_data_228,
  input  [7:0]  io_phv_in_data_229,
  input  [7:0]  io_phv_in_data_230,
  input  [7:0]  io_phv_in_data_231,
  input  [7:0]  io_phv_in_data_232,
  input  [7:0]  io_phv_in_data_233,
  input  [7:0]  io_phv_in_data_234,
  input  [7:0]  io_phv_in_data_235,
  input  [7:0]  io_phv_in_data_236,
  input  [7:0]  io_phv_in_data_237,
  input  [7:0]  io_phv_in_data_238,
  input  [7:0]  io_phv_in_data_239,
  input  [7:0]  io_phv_in_data_240,
  input  [7:0]  io_phv_in_data_241,
  input  [7:0]  io_phv_in_data_242,
  input  [7:0]  io_phv_in_data_243,
  input  [7:0]  io_phv_in_data_244,
  input  [7:0]  io_phv_in_data_245,
  input  [7:0]  io_phv_in_data_246,
  input  [7:0]  io_phv_in_data_247,
  input  [7:0]  io_phv_in_data_248,
  input  [7:0]  io_phv_in_data_249,
  input  [7:0]  io_phv_in_data_250,
  input  [7:0]  io_phv_in_data_251,
  input  [7:0]  io_phv_in_data_252,
  input  [7:0]  io_phv_in_data_253,
  input  [7:0]  io_phv_in_data_254,
  input  [7:0]  io_phv_in_data_255,
  input  [4:0]  io_pcie_o_cs,
  input         io_pcie_o_r_en,
  input  [7:0]  io_pcie_o_r_addr,
  output [63:0] io_pcie_o_r_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  sram_0_clock; // @[outport.scala 23:25]
  wire  sram_0_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_0_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_0_io_w_data; // @[outport.scala 23:25]
  wire  sram_0_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_0_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_0_io_r_data; // @[outport.scala 23:25]
  wire  sram_1_clock; // @[outport.scala 23:25]
  wire  sram_1_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_1_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_1_io_w_data; // @[outport.scala 23:25]
  wire  sram_1_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_1_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_1_io_r_data; // @[outport.scala 23:25]
  wire  sram_2_clock; // @[outport.scala 23:25]
  wire  sram_2_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_2_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_2_io_w_data; // @[outport.scala 23:25]
  wire  sram_2_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_2_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_2_io_r_data; // @[outport.scala 23:25]
  wire  sram_3_clock; // @[outport.scala 23:25]
  wire  sram_3_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_3_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_3_io_w_data; // @[outport.scala 23:25]
  wire  sram_3_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_3_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_3_io_r_data; // @[outport.scala 23:25]
  wire  sram_4_clock; // @[outport.scala 23:25]
  wire  sram_4_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_4_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_4_io_w_data; // @[outport.scala 23:25]
  wire  sram_4_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_4_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_4_io_r_data; // @[outport.scala 23:25]
  wire  sram_5_clock; // @[outport.scala 23:25]
  wire  sram_5_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_5_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_5_io_w_data; // @[outport.scala 23:25]
  wire  sram_5_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_5_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_5_io_r_data; // @[outport.scala 23:25]
  wire  sram_6_clock; // @[outport.scala 23:25]
  wire  sram_6_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_6_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_6_io_w_data; // @[outport.scala 23:25]
  wire  sram_6_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_6_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_6_io_r_data; // @[outport.scala 23:25]
  wire  sram_7_clock; // @[outport.scala 23:25]
  wire  sram_7_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_7_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_7_io_w_data; // @[outport.scala 23:25]
  wire  sram_7_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_7_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_7_io_r_data; // @[outport.scala 23:25]
  wire  sram_8_clock; // @[outport.scala 23:25]
  wire  sram_8_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_8_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_8_io_w_data; // @[outport.scala 23:25]
  wire  sram_8_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_8_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_8_io_r_data; // @[outport.scala 23:25]
  wire  sram_9_clock; // @[outport.scala 23:25]
  wire  sram_9_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_9_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_9_io_w_data; // @[outport.scala 23:25]
  wire  sram_9_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_9_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_9_io_r_data; // @[outport.scala 23:25]
  wire  sram_10_clock; // @[outport.scala 23:25]
  wire  sram_10_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_10_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_10_io_w_data; // @[outport.scala 23:25]
  wire  sram_10_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_10_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_10_io_r_data; // @[outport.scala 23:25]
  wire  sram_11_clock; // @[outport.scala 23:25]
  wire  sram_11_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_11_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_11_io_w_data; // @[outport.scala 23:25]
  wire  sram_11_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_11_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_11_io_r_data; // @[outport.scala 23:25]
  wire  sram_12_clock; // @[outport.scala 23:25]
  wire  sram_12_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_12_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_12_io_w_data; // @[outport.scala 23:25]
  wire  sram_12_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_12_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_12_io_r_data; // @[outport.scala 23:25]
  wire  sram_13_clock; // @[outport.scala 23:25]
  wire  sram_13_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_13_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_13_io_w_data; // @[outport.scala 23:25]
  wire  sram_13_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_13_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_13_io_r_data; // @[outport.scala 23:25]
  wire  sram_14_clock; // @[outport.scala 23:25]
  wire  sram_14_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_14_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_14_io_w_data; // @[outport.scala 23:25]
  wire  sram_14_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_14_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_14_io_r_data; // @[outport.scala 23:25]
  wire  sram_15_clock; // @[outport.scala 23:25]
  wire  sram_15_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_15_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_15_io_w_data; // @[outport.scala 23:25]
  wire  sram_15_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_15_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_15_io_r_data; // @[outport.scala 23:25]
  wire  sram_16_clock; // @[outport.scala 23:25]
  wire  sram_16_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_16_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_16_io_w_data; // @[outport.scala 23:25]
  wire  sram_16_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_16_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_16_io_r_data; // @[outport.scala 23:25]
  wire  sram_17_clock; // @[outport.scala 23:25]
  wire  sram_17_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_17_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_17_io_w_data; // @[outport.scala 23:25]
  wire  sram_17_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_17_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_17_io_r_data; // @[outport.scala 23:25]
  wire  sram_18_clock; // @[outport.scala 23:25]
  wire  sram_18_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_18_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_18_io_w_data; // @[outport.scala 23:25]
  wire  sram_18_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_18_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_18_io_r_data; // @[outport.scala 23:25]
  wire  sram_19_clock; // @[outport.scala 23:25]
  wire  sram_19_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_19_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_19_io_w_data; // @[outport.scala 23:25]
  wire  sram_19_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_19_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_19_io_r_data; // @[outport.scala 23:25]
  wire  sram_20_clock; // @[outport.scala 23:25]
  wire  sram_20_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_20_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_20_io_w_data; // @[outport.scala 23:25]
  wire  sram_20_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_20_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_20_io_r_data; // @[outport.scala 23:25]
  wire  sram_21_clock; // @[outport.scala 23:25]
  wire  sram_21_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_21_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_21_io_w_data; // @[outport.scala 23:25]
  wire  sram_21_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_21_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_21_io_r_data; // @[outport.scala 23:25]
  wire  sram_22_clock; // @[outport.scala 23:25]
  wire  sram_22_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_22_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_22_io_w_data; // @[outport.scala 23:25]
  wire  sram_22_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_22_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_22_io_r_data; // @[outport.scala 23:25]
  wire  sram_23_clock; // @[outport.scala 23:25]
  wire  sram_23_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_23_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_23_io_w_data; // @[outport.scala 23:25]
  wire  sram_23_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_23_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_23_io_r_data; // @[outport.scala 23:25]
  wire  sram_24_clock; // @[outport.scala 23:25]
  wire  sram_24_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_24_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_24_io_w_data; // @[outport.scala 23:25]
  wire  sram_24_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_24_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_24_io_r_data; // @[outport.scala 23:25]
  wire  sram_25_clock; // @[outport.scala 23:25]
  wire  sram_25_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_25_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_25_io_w_data; // @[outport.scala 23:25]
  wire  sram_25_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_25_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_25_io_r_data; // @[outport.scala 23:25]
  wire  sram_26_clock; // @[outport.scala 23:25]
  wire  sram_26_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_26_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_26_io_w_data; // @[outport.scala 23:25]
  wire  sram_26_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_26_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_26_io_r_data; // @[outport.scala 23:25]
  wire  sram_27_clock; // @[outport.scala 23:25]
  wire  sram_27_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_27_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_27_io_w_data; // @[outport.scala 23:25]
  wire  sram_27_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_27_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_27_io_r_data; // @[outport.scala 23:25]
  wire  sram_28_clock; // @[outport.scala 23:25]
  wire  sram_28_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_28_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_28_io_w_data; // @[outport.scala 23:25]
  wire  sram_28_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_28_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_28_io_r_data; // @[outport.scala 23:25]
  wire  sram_29_clock; // @[outport.scala 23:25]
  wire  sram_29_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_29_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_29_io_w_data; // @[outport.scala 23:25]
  wire  sram_29_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_29_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_29_io_r_data; // @[outport.scala 23:25]
  wire  sram_30_clock; // @[outport.scala 23:25]
  wire  sram_30_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_30_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_30_io_w_data; // @[outport.scala 23:25]
  wire  sram_30_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_30_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_30_io_r_data; // @[outport.scala 23:25]
  wire  sram_31_clock; // @[outport.scala 23:25]
  wire  sram_31_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_31_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_31_io_w_data; // @[outport.scala 23:25]
  wire  sram_31_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_31_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_31_io_r_data; // @[outport.scala 23:25]
  reg [7:0] addr; // @[outport.scala 17:19]
  wire [55:0] exe_io_w_data_hi_5 = {io_phv_in_data_0,io_phv_in_data_1,io_phv_in_data_2,io_phv_in_data_3,io_phv_in_data_4
    ,io_phv_in_data_5,io_phv_in_data_6}; // @[Cat.scala 30:58]
  wire  cs_hit = io_pcie_o_cs == 5'h0; // @[outport.scala 31:35]
  wire [63:0] _GEN_0 = cs_hit ? sram_0_io_r_data : 64'h0; // @[outport.scala 34:23 outport.scala 35:31 outport.scala 20:22]
  wire [55:0] exe_io_w_data_hi_11 = {io_phv_in_data_8,io_phv_in_data_9,io_phv_in_data_10,io_phv_in_data_11,
    io_phv_in_data_12,io_phv_in_data_13,io_phv_in_data_14}; // @[Cat.scala 30:58]
  wire  cs_hit_1 = io_pcie_o_cs == 5'h1; // @[outport.scala 31:35]
  wire [63:0] _GEN_1 = cs_hit_1 ? sram_1_io_r_data : _GEN_0; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_17 = {io_phv_in_data_16,io_phv_in_data_17,io_phv_in_data_18,io_phv_in_data_19,
    io_phv_in_data_20,io_phv_in_data_21,io_phv_in_data_22}; // @[Cat.scala 30:58]
  wire  cs_hit_2 = io_pcie_o_cs == 5'h2; // @[outport.scala 31:35]
  wire [63:0] _GEN_2 = cs_hit_2 ? sram_2_io_r_data : _GEN_1; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_23 = {io_phv_in_data_24,io_phv_in_data_25,io_phv_in_data_26,io_phv_in_data_27,
    io_phv_in_data_28,io_phv_in_data_29,io_phv_in_data_30}; // @[Cat.scala 30:58]
  wire  cs_hit_3 = io_pcie_o_cs == 5'h3; // @[outport.scala 31:35]
  wire [63:0] _GEN_3 = cs_hit_3 ? sram_3_io_r_data : _GEN_2; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_29 = {io_phv_in_data_32,io_phv_in_data_33,io_phv_in_data_34,io_phv_in_data_35,
    io_phv_in_data_36,io_phv_in_data_37,io_phv_in_data_38}; // @[Cat.scala 30:58]
  wire  cs_hit_4 = io_pcie_o_cs == 5'h4; // @[outport.scala 31:35]
  wire [63:0] _GEN_4 = cs_hit_4 ? sram_4_io_r_data : _GEN_3; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_35 = {io_phv_in_data_40,io_phv_in_data_41,io_phv_in_data_42,io_phv_in_data_43,
    io_phv_in_data_44,io_phv_in_data_45,io_phv_in_data_46}; // @[Cat.scala 30:58]
  wire  cs_hit_5 = io_pcie_o_cs == 5'h5; // @[outport.scala 31:35]
  wire [63:0] _GEN_5 = cs_hit_5 ? sram_5_io_r_data : _GEN_4; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_41 = {io_phv_in_data_48,io_phv_in_data_49,io_phv_in_data_50,io_phv_in_data_51,
    io_phv_in_data_52,io_phv_in_data_53,io_phv_in_data_54}; // @[Cat.scala 30:58]
  wire  cs_hit_6 = io_pcie_o_cs == 5'h6; // @[outport.scala 31:35]
  wire [63:0] _GEN_6 = cs_hit_6 ? sram_6_io_r_data : _GEN_5; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_47 = {io_phv_in_data_56,io_phv_in_data_57,io_phv_in_data_58,io_phv_in_data_59,
    io_phv_in_data_60,io_phv_in_data_61,io_phv_in_data_62}; // @[Cat.scala 30:58]
  wire  cs_hit_7 = io_pcie_o_cs == 5'h7; // @[outport.scala 31:35]
  wire [63:0] _GEN_7 = cs_hit_7 ? sram_7_io_r_data : _GEN_6; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_53 = {io_phv_in_data_64,io_phv_in_data_65,io_phv_in_data_66,io_phv_in_data_67,
    io_phv_in_data_68,io_phv_in_data_69,io_phv_in_data_70}; // @[Cat.scala 30:58]
  wire  cs_hit_8 = io_pcie_o_cs == 5'h8; // @[outport.scala 31:35]
  wire [63:0] _GEN_8 = cs_hit_8 ? sram_8_io_r_data : _GEN_7; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_59 = {io_phv_in_data_72,io_phv_in_data_73,io_phv_in_data_74,io_phv_in_data_75,
    io_phv_in_data_76,io_phv_in_data_77,io_phv_in_data_78}; // @[Cat.scala 30:58]
  wire  cs_hit_9 = io_pcie_o_cs == 5'h9; // @[outport.scala 31:35]
  wire [63:0] _GEN_9 = cs_hit_9 ? sram_9_io_r_data : _GEN_8; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_65 = {io_phv_in_data_80,io_phv_in_data_81,io_phv_in_data_82,io_phv_in_data_83,
    io_phv_in_data_84,io_phv_in_data_85,io_phv_in_data_86}; // @[Cat.scala 30:58]
  wire  cs_hit_10 = io_pcie_o_cs == 5'ha; // @[outport.scala 31:35]
  wire [63:0] _GEN_10 = cs_hit_10 ? sram_10_io_r_data : _GEN_9; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_71 = {io_phv_in_data_88,io_phv_in_data_89,io_phv_in_data_90,io_phv_in_data_91,
    io_phv_in_data_92,io_phv_in_data_93,io_phv_in_data_94}; // @[Cat.scala 30:58]
  wire  cs_hit_11 = io_pcie_o_cs == 5'hb; // @[outport.scala 31:35]
  wire [63:0] _GEN_11 = cs_hit_11 ? sram_11_io_r_data : _GEN_10; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_77 = {io_phv_in_data_96,io_phv_in_data_97,io_phv_in_data_98,io_phv_in_data_99,
    io_phv_in_data_100,io_phv_in_data_101,io_phv_in_data_102}; // @[Cat.scala 30:58]
  wire  cs_hit_12 = io_pcie_o_cs == 5'hc; // @[outport.scala 31:35]
  wire [63:0] _GEN_12 = cs_hit_12 ? sram_12_io_r_data : _GEN_11; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_83 = {io_phv_in_data_104,io_phv_in_data_105,io_phv_in_data_106,io_phv_in_data_107,
    io_phv_in_data_108,io_phv_in_data_109,io_phv_in_data_110}; // @[Cat.scala 30:58]
  wire  cs_hit_13 = io_pcie_o_cs == 5'hd; // @[outport.scala 31:35]
  wire [63:0] _GEN_13 = cs_hit_13 ? sram_13_io_r_data : _GEN_12; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_89 = {io_phv_in_data_112,io_phv_in_data_113,io_phv_in_data_114,io_phv_in_data_115,
    io_phv_in_data_116,io_phv_in_data_117,io_phv_in_data_118}; // @[Cat.scala 30:58]
  wire  cs_hit_14 = io_pcie_o_cs == 5'he; // @[outport.scala 31:35]
  wire [63:0] _GEN_14 = cs_hit_14 ? sram_14_io_r_data : _GEN_13; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_95 = {io_phv_in_data_120,io_phv_in_data_121,io_phv_in_data_122,io_phv_in_data_123,
    io_phv_in_data_124,io_phv_in_data_125,io_phv_in_data_126}; // @[Cat.scala 30:58]
  wire  cs_hit_15 = io_pcie_o_cs == 5'hf; // @[outport.scala 31:35]
  wire [63:0] _GEN_15 = cs_hit_15 ? sram_15_io_r_data : _GEN_14; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_101 = {io_phv_in_data_128,io_phv_in_data_129,io_phv_in_data_130,io_phv_in_data_131,
    io_phv_in_data_132,io_phv_in_data_133,io_phv_in_data_134}; // @[Cat.scala 30:58]
  wire  cs_hit_16 = io_pcie_o_cs == 5'h10; // @[outport.scala 31:35]
  wire [63:0] _GEN_16 = cs_hit_16 ? sram_16_io_r_data : _GEN_15; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_107 = {io_phv_in_data_136,io_phv_in_data_137,io_phv_in_data_138,io_phv_in_data_139,
    io_phv_in_data_140,io_phv_in_data_141,io_phv_in_data_142}; // @[Cat.scala 30:58]
  wire  cs_hit_17 = io_pcie_o_cs == 5'h11; // @[outport.scala 31:35]
  wire [63:0] _GEN_17 = cs_hit_17 ? sram_17_io_r_data : _GEN_16; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_113 = {io_phv_in_data_144,io_phv_in_data_145,io_phv_in_data_146,io_phv_in_data_147,
    io_phv_in_data_148,io_phv_in_data_149,io_phv_in_data_150}; // @[Cat.scala 30:58]
  wire  cs_hit_18 = io_pcie_o_cs == 5'h12; // @[outport.scala 31:35]
  wire [63:0] _GEN_18 = cs_hit_18 ? sram_18_io_r_data : _GEN_17; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_119 = {io_phv_in_data_152,io_phv_in_data_153,io_phv_in_data_154,io_phv_in_data_155,
    io_phv_in_data_156,io_phv_in_data_157,io_phv_in_data_158}; // @[Cat.scala 30:58]
  wire  cs_hit_19 = io_pcie_o_cs == 5'h13; // @[outport.scala 31:35]
  wire [63:0] _GEN_19 = cs_hit_19 ? sram_19_io_r_data : _GEN_18; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_125 = {io_phv_in_data_160,io_phv_in_data_161,io_phv_in_data_162,io_phv_in_data_163,
    io_phv_in_data_164,io_phv_in_data_165,io_phv_in_data_166}; // @[Cat.scala 30:58]
  wire  cs_hit_20 = io_pcie_o_cs == 5'h14; // @[outport.scala 31:35]
  wire [63:0] _GEN_20 = cs_hit_20 ? sram_20_io_r_data : _GEN_19; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_131 = {io_phv_in_data_168,io_phv_in_data_169,io_phv_in_data_170,io_phv_in_data_171,
    io_phv_in_data_172,io_phv_in_data_173,io_phv_in_data_174}; // @[Cat.scala 30:58]
  wire  cs_hit_21 = io_pcie_o_cs == 5'h15; // @[outport.scala 31:35]
  wire [63:0] _GEN_21 = cs_hit_21 ? sram_21_io_r_data : _GEN_20; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_137 = {io_phv_in_data_176,io_phv_in_data_177,io_phv_in_data_178,io_phv_in_data_179,
    io_phv_in_data_180,io_phv_in_data_181,io_phv_in_data_182}; // @[Cat.scala 30:58]
  wire  cs_hit_22 = io_pcie_o_cs == 5'h16; // @[outport.scala 31:35]
  wire [63:0] _GEN_22 = cs_hit_22 ? sram_22_io_r_data : _GEN_21; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_143 = {io_phv_in_data_184,io_phv_in_data_185,io_phv_in_data_186,io_phv_in_data_187,
    io_phv_in_data_188,io_phv_in_data_189,io_phv_in_data_190}; // @[Cat.scala 30:58]
  wire  cs_hit_23 = io_pcie_o_cs == 5'h17; // @[outport.scala 31:35]
  wire [63:0] _GEN_23 = cs_hit_23 ? sram_23_io_r_data : _GEN_22; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_149 = {io_phv_in_data_192,io_phv_in_data_193,io_phv_in_data_194,io_phv_in_data_195,
    io_phv_in_data_196,io_phv_in_data_197,io_phv_in_data_198}; // @[Cat.scala 30:58]
  wire  cs_hit_24 = io_pcie_o_cs == 5'h18; // @[outport.scala 31:35]
  wire [63:0] _GEN_24 = cs_hit_24 ? sram_24_io_r_data : _GEN_23; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_155 = {io_phv_in_data_200,io_phv_in_data_201,io_phv_in_data_202,io_phv_in_data_203,
    io_phv_in_data_204,io_phv_in_data_205,io_phv_in_data_206}; // @[Cat.scala 30:58]
  wire  cs_hit_25 = io_pcie_o_cs == 5'h19; // @[outport.scala 31:35]
  wire [63:0] _GEN_25 = cs_hit_25 ? sram_25_io_r_data : _GEN_24; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_161 = {io_phv_in_data_208,io_phv_in_data_209,io_phv_in_data_210,io_phv_in_data_211,
    io_phv_in_data_212,io_phv_in_data_213,io_phv_in_data_214}; // @[Cat.scala 30:58]
  wire  cs_hit_26 = io_pcie_o_cs == 5'h1a; // @[outport.scala 31:35]
  wire [63:0] _GEN_26 = cs_hit_26 ? sram_26_io_r_data : _GEN_25; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_167 = {io_phv_in_data_216,io_phv_in_data_217,io_phv_in_data_218,io_phv_in_data_219,
    io_phv_in_data_220,io_phv_in_data_221,io_phv_in_data_222}; // @[Cat.scala 30:58]
  wire  cs_hit_27 = io_pcie_o_cs == 5'h1b; // @[outport.scala 31:35]
  wire [63:0] _GEN_27 = cs_hit_27 ? sram_27_io_r_data : _GEN_26; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_173 = {io_phv_in_data_224,io_phv_in_data_225,io_phv_in_data_226,io_phv_in_data_227,
    io_phv_in_data_228,io_phv_in_data_229,io_phv_in_data_230}; // @[Cat.scala 30:58]
  wire  cs_hit_28 = io_pcie_o_cs == 5'h1c; // @[outport.scala 31:35]
  wire [63:0] _GEN_28 = cs_hit_28 ? sram_28_io_r_data : _GEN_27; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_179 = {io_phv_in_data_232,io_phv_in_data_233,io_phv_in_data_234,io_phv_in_data_235,
    io_phv_in_data_236,io_phv_in_data_237,io_phv_in_data_238}; // @[Cat.scala 30:58]
  wire  cs_hit_29 = io_pcie_o_cs == 5'h1d; // @[outport.scala 31:35]
  wire [63:0] _GEN_29 = cs_hit_29 ? sram_29_io_r_data : _GEN_28; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_185 = {io_phv_in_data_240,io_phv_in_data_241,io_phv_in_data_242,io_phv_in_data_243,
    io_phv_in_data_244,io_phv_in_data_245,io_phv_in_data_246}; // @[Cat.scala 30:58]
  wire  cs_hit_30 = io_pcie_o_cs == 5'h1e; // @[outport.scala 31:35]
  wire [63:0] _GEN_30 = cs_hit_30 ? sram_30_io_r_data : _GEN_29; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_191 = {io_phv_in_data_248,io_phv_in_data_249,io_phv_in_data_250,io_phv_in_data_251,
    io_phv_in_data_252,io_phv_in_data_253,io_phv_in_data_254}; // @[Cat.scala 30:58]
  wire  cs_hit_31 = io_pcie_o_cs == 5'h1f; // @[outport.scala 31:35]
  SRAM sram_0 ( // @[outport.scala 23:25]
    .clock(sram_0_clock),
    .io_w_en(sram_0_io_w_en),
    .io_w_addr(sram_0_io_w_addr),
    .io_w_data(sram_0_io_w_data),
    .io_r_en(sram_0_io_r_en),
    .io_r_addr(sram_0_io_r_addr),
    .io_r_data(sram_0_io_r_data)
  );
  SRAM sram_1 ( // @[outport.scala 23:25]
    .clock(sram_1_clock),
    .io_w_en(sram_1_io_w_en),
    .io_w_addr(sram_1_io_w_addr),
    .io_w_data(sram_1_io_w_data),
    .io_r_en(sram_1_io_r_en),
    .io_r_addr(sram_1_io_r_addr),
    .io_r_data(sram_1_io_r_data)
  );
  SRAM sram_2 ( // @[outport.scala 23:25]
    .clock(sram_2_clock),
    .io_w_en(sram_2_io_w_en),
    .io_w_addr(sram_2_io_w_addr),
    .io_w_data(sram_2_io_w_data),
    .io_r_en(sram_2_io_r_en),
    .io_r_addr(sram_2_io_r_addr),
    .io_r_data(sram_2_io_r_data)
  );
  SRAM sram_3 ( // @[outport.scala 23:25]
    .clock(sram_3_clock),
    .io_w_en(sram_3_io_w_en),
    .io_w_addr(sram_3_io_w_addr),
    .io_w_data(sram_3_io_w_data),
    .io_r_en(sram_3_io_r_en),
    .io_r_addr(sram_3_io_r_addr),
    .io_r_data(sram_3_io_r_data)
  );
  SRAM sram_4 ( // @[outport.scala 23:25]
    .clock(sram_4_clock),
    .io_w_en(sram_4_io_w_en),
    .io_w_addr(sram_4_io_w_addr),
    .io_w_data(sram_4_io_w_data),
    .io_r_en(sram_4_io_r_en),
    .io_r_addr(sram_4_io_r_addr),
    .io_r_data(sram_4_io_r_data)
  );
  SRAM sram_5 ( // @[outport.scala 23:25]
    .clock(sram_5_clock),
    .io_w_en(sram_5_io_w_en),
    .io_w_addr(sram_5_io_w_addr),
    .io_w_data(sram_5_io_w_data),
    .io_r_en(sram_5_io_r_en),
    .io_r_addr(sram_5_io_r_addr),
    .io_r_data(sram_5_io_r_data)
  );
  SRAM sram_6 ( // @[outport.scala 23:25]
    .clock(sram_6_clock),
    .io_w_en(sram_6_io_w_en),
    .io_w_addr(sram_6_io_w_addr),
    .io_w_data(sram_6_io_w_data),
    .io_r_en(sram_6_io_r_en),
    .io_r_addr(sram_6_io_r_addr),
    .io_r_data(sram_6_io_r_data)
  );
  SRAM sram_7 ( // @[outport.scala 23:25]
    .clock(sram_7_clock),
    .io_w_en(sram_7_io_w_en),
    .io_w_addr(sram_7_io_w_addr),
    .io_w_data(sram_7_io_w_data),
    .io_r_en(sram_7_io_r_en),
    .io_r_addr(sram_7_io_r_addr),
    .io_r_data(sram_7_io_r_data)
  );
  SRAM sram_8 ( // @[outport.scala 23:25]
    .clock(sram_8_clock),
    .io_w_en(sram_8_io_w_en),
    .io_w_addr(sram_8_io_w_addr),
    .io_w_data(sram_8_io_w_data),
    .io_r_en(sram_8_io_r_en),
    .io_r_addr(sram_8_io_r_addr),
    .io_r_data(sram_8_io_r_data)
  );
  SRAM sram_9 ( // @[outport.scala 23:25]
    .clock(sram_9_clock),
    .io_w_en(sram_9_io_w_en),
    .io_w_addr(sram_9_io_w_addr),
    .io_w_data(sram_9_io_w_data),
    .io_r_en(sram_9_io_r_en),
    .io_r_addr(sram_9_io_r_addr),
    .io_r_data(sram_9_io_r_data)
  );
  SRAM sram_10 ( // @[outport.scala 23:25]
    .clock(sram_10_clock),
    .io_w_en(sram_10_io_w_en),
    .io_w_addr(sram_10_io_w_addr),
    .io_w_data(sram_10_io_w_data),
    .io_r_en(sram_10_io_r_en),
    .io_r_addr(sram_10_io_r_addr),
    .io_r_data(sram_10_io_r_data)
  );
  SRAM sram_11 ( // @[outport.scala 23:25]
    .clock(sram_11_clock),
    .io_w_en(sram_11_io_w_en),
    .io_w_addr(sram_11_io_w_addr),
    .io_w_data(sram_11_io_w_data),
    .io_r_en(sram_11_io_r_en),
    .io_r_addr(sram_11_io_r_addr),
    .io_r_data(sram_11_io_r_data)
  );
  SRAM sram_12 ( // @[outport.scala 23:25]
    .clock(sram_12_clock),
    .io_w_en(sram_12_io_w_en),
    .io_w_addr(sram_12_io_w_addr),
    .io_w_data(sram_12_io_w_data),
    .io_r_en(sram_12_io_r_en),
    .io_r_addr(sram_12_io_r_addr),
    .io_r_data(sram_12_io_r_data)
  );
  SRAM sram_13 ( // @[outport.scala 23:25]
    .clock(sram_13_clock),
    .io_w_en(sram_13_io_w_en),
    .io_w_addr(sram_13_io_w_addr),
    .io_w_data(sram_13_io_w_data),
    .io_r_en(sram_13_io_r_en),
    .io_r_addr(sram_13_io_r_addr),
    .io_r_data(sram_13_io_r_data)
  );
  SRAM sram_14 ( // @[outport.scala 23:25]
    .clock(sram_14_clock),
    .io_w_en(sram_14_io_w_en),
    .io_w_addr(sram_14_io_w_addr),
    .io_w_data(sram_14_io_w_data),
    .io_r_en(sram_14_io_r_en),
    .io_r_addr(sram_14_io_r_addr),
    .io_r_data(sram_14_io_r_data)
  );
  SRAM sram_15 ( // @[outport.scala 23:25]
    .clock(sram_15_clock),
    .io_w_en(sram_15_io_w_en),
    .io_w_addr(sram_15_io_w_addr),
    .io_w_data(sram_15_io_w_data),
    .io_r_en(sram_15_io_r_en),
    .io_r_addr(sram_15_io_r_addr),
    .io_r_data(sram_15_io_r_data)
  );
  SRAM sram_16 ( // @[outport.scala 23:25]
    .clock(sram_16_clock),
    .io_w_en(sram_16_io_w_en),
    .io_w_addr(sram_16_io_w_addr),
    .io_w_data(sram_16_io_w_data),
    .io_r_en(sram_16_io_r_en),
    .io_r_addr(sram_16_io_r_addr),
    .io_r_data(sram_16_io_r_data)
  );
  SRAM sram_17 ( // @[outport.scala 23:25]
    .clock(sram_17_clock),
    .io_w_en(sram_17_io_w_en),
    .io_w_addr(sram_17_io_w_addr),
    .io_w_data(sram_17_io_w_data),
    .io_r_en(sram_17_io_r_en),
    .io_r_addr(sram_17_io_r_addr),
    .io_r_data(sram_17_io_r_data)
  );
  SRAM sram_18 ( // @[outport.scala 23:25]
    .clock(sram_18_clock),
    .io_w_en(sram_18_io_w_en),
    .io_w_addr(sram_18_io_w_addr),
    .io_w_data(sram_18_io_w_data),
    .io_r_en(sram_18_io_r_en),
    .io_r_addr(sram_18_io_r_addr),
    .io_r_data(sram_18_io_r_data)
  );
  SRAM sram_19 ( // @[outport.scala 23:25]
    .clock(sram_19_clock),
    .io_w_en(sram_19_io_w_en),
    .io_w_addr(sram_19_io_w_addr),
    .io_w_data(sram_19_io_w_data),
    .io_r_en(sram_19_io_r_en),
    .io_r_addr(sram_19_io_r_addr),
    .io_r_data(sram_19_io_r_data)
  );
  SRAM sram_20 ( // @[outport.scala 23:25]
    .clock(sram_20_clock),
    .io_w_en(sram_20_io_w_en),
    .io_w_addr(sram_20_io_w_addr),
    .io_w_data(sram_20_io_w_data),
    .io_r_en(sram_20_io_r_en),
    .io_r_addr(sram_20_io_r_addr),
    .io_r_data(sram_20_io_r_data)
  );
  SRAM sram_21 ( // @[outport.scala 23:25]
    .clock(sram_21_clock),
    .io_w_en(sram_21_io_w_en),
    .io_w_addr(sram_21_io_w_addr),
    .io_w_data(sram_21_io_w_data),
    .io_r_en(sram_21_io_r_en),
    .io_r_addr(sram_21_io_r_addr),
    .io_r_data(sram_21_io_r_data)
  );
  SRAM sram_22 ( // @[outport.scala 23:25]
    .clock(sram_22_clock),
    .io_w_en(sram_22_io_w_en),
    .io_w_addr(sram_22_io_w_addr),
    .io_w_data(sram_22_io_w_data),
    .io_r_en(sram_22_io_r_en),
    .io_r_addr(sram_22_io_r_addr),
    .io_r_data(sram_22_io_r_data)
  );
  SRAM sram_23 ( // @[outport.scala 23:25]
    .clock(sram_23_clock),
    .io_w_en(sram_23_io_w_en),
    .io_w_addr(sram_23_io_w_addr),
    .io_w_data(sram_23_io_w_data),
    .io_r_en(sram_23_io_r_en),
    .io_r_addr(sram_23_io_r_addr),
    .io_r_data(sram_23_io_r_data)
  );
  SRAM sram_24 ( // @[outport.scala 23:25]
    .clock(sram_24_clock),
    .io_w_en(sram_24_io_w_en),
    .io_w_addr(sram_24_io_w_addr),
    .io_w_data(sram_24_io_w_data),
    .io_r_en(sram_24_io_r_en),
    .io_r_addr(sram_24_io_r_addr),
    .io_r_data(sram_24_io_r_data)
  );
  SRAM sram_25 ( // @[outport.scala 23:25]
    .clock(sram_25_clock),
    .io_w_en(sram_25_io_w_en),
    .io_w_addr(sram_25_io_w_addr),
    .io_w_data(sram_25_io_w_data),
    .io_r_en(sram_25_io_r_en),
    .io_r_addr(sram_25_io_r_addr),
    .io_r_data(sram_25_io_r_data)
  );
  SRAM sram_26 ( // @[outport.scala 23:25]
    .clock(sram_26_clock),
    .io_w_en(sram_26_io_w_en),
    .io_w_addr(sram_26_io_w_addr),
    .io_w_data(sram_26_io_w_data),
    .io_r_en(sram_26_io_r_en),
    .io_r_addr(sram_26_io_r_addr),
    .io_r_data(sram_26_io_r_data)
  );
  SRAM sram_27 ( // @[outport.scala 23:25]
    .clock(sram_27_clock),
    .io_w_en(sram_27_io_w_en),
    .io_w_addr(sram_27_io_w_addr),
    .io_w_data(sram_27_io_w_data),
    .io_r_en(sram_27_io_r_en),
    .io_r_addr(sram_27_io_r_addr),
    .io_r_data(sram_27_io_r_data)
  );
  SRAM sram_28 ( // @[outport.scala 23:25]
    .clock(sram_28_clock),
    .io_w_en(sram_28_io_w_en),
    .io_w_addr(sram_28_io_w_addr),
    .io_w_data(sram_28_io_w_data),
    .io_r_en(sram_28_io_r_en),
    .io_r_addr(sram_28_io_r_addr),
    .io_r_data(sram_28_io_r_data)
  );
  SRAM sram_29 ( // @[outport.scala 23:25]
    .clock(sram_29_clock),
    .io_w_en(sram_29_io_w_en),
    .io_w_addr(sram_29_io_w_addr),
    .io_w_data(sram_29_io_w_data),
    .io_r_en(sram_29_io_r_en),
    .io_r_addr(sram_29_io_r_addr),
    .io_r_data(sram_29_io_r_data)
  );
  SRAM sram_30 ( // @[outport.scala 23:25]
    .clock(sram_30_clock),
    .io_w_en(sram_30_io_w_en),
    .io_w_addr(sram_30_io_w_addr),
    .io_w_data(sram_30_io_w_data),
    .io_r_en(sram_30_io_r_en),
    .io_r_addr(sram_30_io_r_addr),
    .io_r_data(sram_30_io_r_data)
  );
  SRAM sram_31 ( // @[outport.scala 23:25]
    .clock(sram_31_clock),
    .io_w_en(sram_31_io_w_en),
    .io_w_addr(sram_31_io_w_addr),
    .io_w_data(sram_31_io_w_data),
    .io_r_en(sram_31_io_r_en),
    .io_r_addr(sram_31_io_r_addr),
    .io_r_data(sram_31_io_r_data)
  );
  assign io_pcie_o_r_data = cs_hit_31 ? sram_31_io_r_data : _GEN_30; // @[outport.scala 34:23 outport.scala 35:31]
  assign sram_0_clock = clock;
  assign sram_0_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_0_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_0_io_w_data = {exe_io_w_data_hi_5,io_phv_in_data_7}; // @[Cat.scala 30:58]
  assign sram_0_io_r_en = io_pcie_o_r_en & cs_hit; // @[outport.scala 32:42]
  assign sram_0_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_1_clock = clock;
  assign sram_1_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_1_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_1_io_w_data = {exe_io_w_data_hi_11,io_phv_in_data_15}; // @[Cat.scala 30:58]
  assign sram_1_io_r_en = io_pcie_o_r_en & cs_hit_1; // @[outport.scala 32:42]
  assign sram_1_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_2_clock = clock;
  assign sram_2_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_2_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_2_io_w_data = {exe_io_w_data_hi_17,io_phv_in_data_23}; // @[Cat.scala 30:58]
  assign sram_2_io_r_en = io_pcie_o_r_en & cs_hit_2; // @[outport.scala 32:42]
  assign sram_2_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_3_clock = clock;
  assign sram_3_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_3_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_3_io_w_data = {exe_io_w_data_hi_23,io_phv_in_data_31}; // @[Cat.scala 30:58]
  assign sram_3_io_r_en = io_pcie_o_r_en & cs_hit_3; // @[outport.scala 32:42]
  assign sram_3_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_4_clock = clock;
  assign sram_4_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_4_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_4_io_w_data = {exe_io_w_data_hi_29,io_phv_in_data_39}; // @[Cat.scala 30:58]
  assign sram_4_io_r_en = io_pcie_o_r_en & cs_hit_4; // @[outport.scala 32:42]
  assign sram_4_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_5_clock = clock;
  assign sram_5_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_5_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_5_io_w_data = {exe_io_w_data_hi_35,io_phv_in_data_47}; // @[Cat.scala 30:58]
  assign sram_5_io_r_en = io_pcie_o_r_en & cs_hit_5; // @[outport.scala 32:42]
  assign sram_5_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_6_clock = clock;
  assign sram_6_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_6_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_6_io_w_data = {exe_io_w_data_hi_41,io_phv_in_data_55}; // @[Cat.scala 30:58]
  assign sram_6_io_r_en = io_pcie_o_r_en & cs_hit_6; // @[outport.scala 32:42]
  assign sram_6_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_7_clock = clock;
  assign sram_7_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_7_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_7_io_w_data = {exe_io_w_data_hi_47,io_phv_in_data_63}; // @[Cat.scala 30:58]
  assign sram_7_io_r_en = io_pcie_o_r_en & cs_hit_7; // @[outport.scala 32:42]
  assign sram_7_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_8_clock = clock;
  assign sram_8_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_8_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_8_io_w_data = {exe_io_w_data_hi_53,io_phv_in_data_71}; // @[Cat.scala 30:58]
  assign sram_8_io_r_en = io_pcie_o_r_en & cs_hit_8; // @[outport.scala 32:42]
  assign sram_8_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_9_clock = clock;
  assign sram_9_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_9_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_9_io_w_data = {exe_io_w_data_hi_59,io_phv_in_data_79}; // @[Cat.scala 30:58]
  assign sram_9_io_r_en = io_pcie_o_r_en & cs_hit_9; // @[outport.scala 32:42]
  assign sram_9_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_10_clock = clock;
  assign sram_10_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_10_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_10_io_w_data = {exe_io_w_data_hi_65,io_phv_in_data_87}; // @[Cat.scala 30:58]
  assign sram_10_io_r_en = io_pcie_o_r_en & cs_hit_10; // @[outport.scala 32:42]
  assign sram_10_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_11_clock = clock;
  assign sram_11_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_11_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_11_io_w_data = {exe_io_w_data_hi_71,io_phv_in_data_95}; // @[Cat.scala 30:58]
  assign sram_11_io_r_en = io_pcie_o_r_en & cs_hit_11; // @[outport.scala 32:42]
  assign sram_11_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_12_clock = clock;
  assign sram_12_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_12_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_12_io_w_data = {exe_io_w_data_hi_77,io_phv_in_data_103}; // @[Cat.scala 30:58]
  assign sram_12_io_r_en = io_pcie_o_r_en & cs_hit_12; // @[outport.scala 32:42]
  assign sram_12_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_13_clock = clock;
  assign sram_13_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_13_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_13_io_w_data = {exe_io_w_data_hi_83,io_phv_in_data_111}; // @[Cat.scala 30:58]
  assign sram_13_io_r_en = io_pcie_o_r_en & cs_hit_13; // @[outport.scala 32:42]
  assign sram_13_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_14_clock = clock;
  assign sram_14_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_14_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_14_io_w_data = {exe_io_w_data_hi_89,io_phv_in_data_119}; // @[Cat.scala 30:58]
  assign sram_14_io_r_en = io_pcie_o_r_en & cs_hit_14; // @[outport.scala 32:42]
  assign sram_14_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_15_clock = clock;
  assign sram_15_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_15_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_15_io_w_data = {exe_io_w_data_hi_95,io_phv_in_data_127}; // @[Cat.scala 30:58]
  assign sram_15_io_r_en = io_pcie_o_r_en & cs_hit_15; // @[outport.scala 32:42]
  assign sram_15_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_16_clock = clock;
  assign sram_16_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_16_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_16_io_w_data = {exe_io_w_data_hi_101,io_phv_in_data_135}; // @[Cat.scala 30:58]
  assign sram_16_io_r_en = io_pcie_o_r_en & cs_hit_16; // @[outport.scala 32:42]
  assign sram_16_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_17_clock = clock;
  assign sram_17_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_17_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_17_io_w_data = {exe_io_w_data_hi_107,io_phv_in_data_143}; // @[Cat.scala 30:58]
  assign sram_17_io_r_en = io_pcie_o_r_en & cs_hit_17; // @[outport.scala 32:42]
  assign sram_17_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_18_clock = clock;
  assign sram_18_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_18_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_18_io_w_data = {exe_io_w_data_hi_113,io_phv_in_data_151}; // @[Cat.scala 30:58]
  assign sram_18_io_r_en = io_pcie_o_r_en & cs_hit_18; // @[outport.scala 32:42]
  assign sram_18_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_19_clock = clock;
  assign sram_19_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_19_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_19_io_w_data = {exe_io_w_data_hi_119,io_phv_in_data_159}; // @[Cat.scala 30:58]
  assign sram_19_io_r_en = io_pcie_o_r_en & cs_hit_19; // @[outport.scala 32:42]
  assign sram_19_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_20_clock = clock;
  assign sram_20_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_20_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_20_io_w_data = {exe_io_w_data_hi_125,io_phv_in_data_167}; // @[Cat.scala 30:58]
  assign sram_20_io_r_en = io_pcie_o_r_en & cs_hit_20; // @[outport.scala 32:42]
  assign sram_20_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_21_clock = clock;
  assign sram_21_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_21_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_21_io_w_data = {exe_io_w_data_hi_131,io_phv_in_data_175}; // @[Cat.scala 30:58]
  assign sram_21_io_r_en = io_pcie_o_r_en & cs_hit_21; // @[outport.scala 32:42]
  assign sram_21_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_22_clock = clock;
  assign sram_22_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_22_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_22_io_w_data = {exe_io_w_data_hi_137,io_phv_in_data_183}; // @[Cat.scala 30:58]
  assign sram_22_io_r_en = io_pcie_o_r_en & cs_hit_22; // @[outport.scala 32:42]
  assign sram_22_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_23_clock = clock;
  assign sram_23_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_23_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_23_io_w_data = {exe_io_w_data_hi_143,io_phv_in_data_191}; // @[Cat.scala 30:58]
  assign sram_23_io_r_en = io_pcie_o_r_en & cs_hit_23; // @[outport.scala 32:42]
  assign sram_23_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_24_clock = clock;
  assign sram_24_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_24_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_24_io_w_data = {exe_io_w_data_hi_149,io_phv_in_data_199}; // @[Cat.scala 30:58]
  assign sram_24_io_r_en = io_pcie_o_r_en & cs_hit_24; // @[outport.scala 32:42]
  assign sram_24_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_25_clock = clock;
  assign sram_25_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_25_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_25_io_w_data = {exe_io_w_data_hi_155,io_phv_in_data_207}; // @[Cat.scala 30:58]
  assign sram_25_io_r_en = io_pcie_o_r_en & cs_hit_25; // @[outport.scala 32:42]
  assign sram_25_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_26_clock = clock;
  assign sram_26_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_26_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_26_io_w_data = {exe_io_w_data_hi_161,io_phv_in_data_215}; // @[Cat.scala 30:58]
  assign sram_26_io_r_en = io_pcie_o_r_en & cs_hit_26; // @[outport.scala 32:42]
  assign sram_26_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_27_clock = clock;
  assign sram_27_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_27_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_27_io_w_data = {exe_io_w_data_hi_167,io_phv_in_data_223}; // @[Cat.scala 30:58]
  assign sram_27_io_r_en = io_pcie_o_r_en & cs_hit_27; // @[outport.scala 32:42]
  assign sram_27_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_28_clock = clock;
  assign sram_28_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_28_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_28_io_w_data = {exe_io_w_data_hi_173,io_phv_in_data_231}; // @[Cat.scala 30:58]
  assign sram_28_io_r_en = io_pcie_o_r_en & cs_hit_28; // @[outport.scala 32:42]
  assign sram_28_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_29_clock = clock;
  assign sram_29_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_29_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_29_io_w_data = {exe_io_w_data_hi_179,io_phv_in_data_239}; // @[Cat.scala 30:58]
  assign sram_29_io_r_en = io_pcie_o_r_en & cs_hit_29; // @[outport.scala 32:42]
  assign sram_29_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_30_clock = clock;
  assign sram_30_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_30_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_30_io_w_data = {exe_io_w_data_hi_185,io_phv_in_data_247}; // @[Cat.scala 30:58]
  assign sram_30_io_r_en = io_pcie_o_r_en & cs_hit_30; // @[outport.scala 32:42]
  assign sram_30_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_31_clock = clock;
  assign sram_31_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_31_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_31_io_w_data = {exe_io_w_data_hi_191,io_phv_in_data_255}; // @[Cat.scala 30:58]
  assign sram_31_io_r_en = io_pcie_o_r_en & cs_hit_31; // @[outport.scala 32:42]
  assign sram_31_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  always @(posedge clock) begin
    addr <= addr + 8'h1; // @[outport.scala 18:18]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr = _RAND_0[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
