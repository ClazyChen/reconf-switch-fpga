module PISA(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [7:0]  io_pipe_phv_in_data_160,
  input  [7:0]  io_pipe_phv_in_data_161,
  input  [7:0]  io_pipe_phv_in_data_162,
  input  [7:0]  io_pipe_phv_in_data_163,
  input  [7:0]  io_pipe_phv_in_data_164,
  input  [7:0]  io_pipe_phv_in_data_165,
  input  [7:0]  io_pipe_phv_in_data_166,
  input  [7:0]  io_pipe_phv_in_data_167,
  input  [7:0]  io_pipe_phv_in_data_168,
  input  [7:0]  io_pipe_phv_in_data_169,
  input  [7:0]  io_pipe_phv_in_data_170,
  input  [7:0]  io_pipe_phv_in_data_171,
  input  [7:0]  io_pipe_phv_in_data_172,
  input  [7:0]  io_pipe_phv_in_data_173,
  input  [7:0]  io_pipe_phv_in_data_174,
  input  [7:0]  io_pipe_phv_in_data_175,
  input  [7:0]  io_pipe_phv_in_data_176,
  input  [7:0]  io_pipe_phv_in_data_177,
  input  [7:0]  io_pipe_phv_in_data_178,
  input  [7:0]  io_pipe_phv_in_data_179,
  input  [7:0]  io_pipe_phv_in_data_180,
  input  [7:0]  io_pipe_phv_in_data_181,
  input  [7:0]  io_pipe_phv_in_data_182,
  input  [7:0]  io_pipe_phv_in_data_183,
  input  [7:0]  io_pipe_phv_in_data_184,
  input  [7:0]  io_pipe_phv_in_data_185,
  input  [7:0]  io_pipe_phv_in_data_186,
  input  [7:0]  io_pipe_phv_in_data_187,
  input  [7:0]  io_pipe_phv_in_data_188,
  input  [7:0]  io_pipe_phv_in_data_189,
  input  [7:0]  io_pipe_phv_in_data_190,
  input  [7:0]  io_pipe_phv_in_data_191,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [7:0]  io_pipe_phv_out_data_160,
  output [7:0]  io_pipe_phv_out_data_161,
  output [7:0]  io_pipe_phv_out_data_162,
  output [7:0]  io_pipe_phv_out_data_163,
  output [7:0]  io_pipe_phv_out_data_164,
  output [7:0]  io_pipe_phv_out_data_165,
  output [7:0]  io_pipe_phv_out_data_166,
  output [7:0]  io_pipe_phv_out_data_167,
  output [7:0]  io_pipe_phv_out_data_168,
  output [7:0]  io_pipe_phv_out_data_169,
  output [7:0]  io_pipe_phv_out_data_170,
  output [7:0]  io_pipe_phv_out_data_171,
  output [7:0]  io_pipe_phv_out_data_172,
  output [7:0]  io_pipe_phv_out_data_173,
  output [7:0]  io_pipe_phv_out_data_174,
  output [7:0]  io_pipe_phv_out_data_175,
  output [7:0]  io_pipe_phv_out_data_176,
  output [7:0]  io_pipe_phv_out_data_177,
  output [7:0]  io_pipe_phv_out_data_178,
  output [7:0]  io_pipe_phv_out_data_179,
  output [7:0]  io_pipe_phv_out_data_180,
  output [7:0]  io_pipe_phv_out_data_181,
  output [7:0]  io_pipe_phv_out_data_182,
  output [7:0]  io_pipe_phv_out_data_183,
  output [7:0]  io_pipe_phv_out_data_184,
  output [7:0]  io_pipe_phv_out_data_185,
  output [7:0]  io_pipe_phv_out_data_186,
  output [7:0]  io_pipe_phv_out_data_187,
  output [7:0]  io_pipe_phv_out_data_188,
  output [7:0]  io_pipe_phv_out_data_189,
  output [7:0]  io_pipe_phv_out_data_190,
  output [7:0]  io_pipe_phv_out_data_191,
  output [7:0]  io_pipe_phv_out_data_192,
  output [7:0]  io_pipe_phv_out_data_193,
  output [7:0]  io_pipe_phv_out_data_194,
  output [7:0]  io_pipe_phv_out_data_195,
  output [7:0]  io_pipe_phv_out_data_196,
  output [7:0]  io_pipe_phv_out_data_197,
  output [7:0]  io_pipe_phv_out_data_198,
  output [7:0]  io_pipe_phv_out_data_199,
  output [7:0]  io_pipe_phv_out_data_200,
  output [7:0]  io_pipe_phv_out_data_201,
  output [7:0]  io_pipe_phv_out_data_202,
  output [7:0]  io_pipe_phv_out_data_203,
  output [7:0]  io_pipe_phv_out_data_204,
  output [7:0]  io_pipe_phv_out_data_205,
  output [7:0]  io_pipe_phv_out_data_206,
  output [7:0]  io_pipe_phv_out_data_207,
  output [7:0]  io_pipe_phv_out_data_208,
  output [7:0]  io_pipe_phv_out_data_209,
  output [7:0]  io_pipe_phv_out_data_210,
  output [7:0]  io_pipe_phv_out_data_211,
  output [7:0]  io_pipe_phv_out_data_212,
  output [7:0]  io_pipe_phv_out_data_213,
  output [7:0]  io_pipe_phv_out_data_214,
  output [7:0]  io_pipe_phv_out_data_215,
  output [7:0]  io_pipe_phv_out_data_216,
  output [7:0]  io_pipe_phv_out_data_217,
  output [7:0]  io_pipe_phv_out_data_218,
  output [7:0]  io_pipe_phv_out_data_219,
  output [7:0]  io_pipe_phv_out_data_220,
  output [7:0]  io_pipe_phv_out_data_221,
  output [7:0]  io_pipe_phv_out_data_222,
  output [7:0]  io_pipe_phv_out_data_223,
  output [7:0]  io_pipe_phv_out_data_224,
  output [7:0]  io_pipe_phv_out_data_225,
  output [7:0]  io_pipe_phv_out_data_226,
  output [7:0]  io_pipe_phv_out_data_227,
  output [7:0]  io_pipe_phv_out_data_228,
  output [7:0]  io_pipe_phv_out_data_229,
  output [7:0]  io_pipe_phv_out_data_230,
  output [7:0]  io_pipe_phv_out_data_231,
  output [7:0]  io_pipe_phv_out_data_232,
  output [7:0]  io_pipe_phv_out_data_233,
  output [7:0]  io_pipe_phv_out_data_234,
  output [7:0]  io_pipe_phv_out_data_235,
  output [7:0]  io_pipe_phv_out_data_236,
  output [7:0]  io_pipe_phv_out_data_237,
  output [7:0]  io_pipe_phv_out_data_238,
  output [7:0]  io_pipe_phv_out_data_239,
  output [7:0]  io_pipe_phv_out_data_240,
  output [7:0]  io_pipe_phv_out_data_241,
  output [7:0]  io_pipe_phv_out_data_242,
  output [7:0]  io_pipe_phv_out_data_243,
  output [7:0]  io_pipe_phv_out_data_244,
  output [7:0]  io_pipe_phv_out_data_245,
  output [7:0]  io_pipe_phv_out_data_246,
  output [7:0]  io_pipe_phv_out_data_247,
  output [7:0]  io_pipe_phv_out_data_248,
  output [7:0]  io_pipe_phv_out_data_249,
  output [7:0]  io_pipe_phv_out_data_250,
  output [7:0]  io_pipe_phv_out_data_251,
  output [7:0]  io_pipe_phv_out_data_252,
  output [7:0]  io_pipe_phv_out_data_253,
  output [7:0]  io_pipe_phv_out_data_254,
  output [7:0]  io_pipe_phv_out_data_255,
  input         io_mod_par_mod_en,
  input         io_mod_par_mod_last_mau_id_mod,
  input  [3:0]  io_mod_par_mod_last_mau_id,
  input  [2:0]  io_mod_par_mod_cs,
  input         io_mod_par_mod_module_mod_state_id_mod,
  input  [7:0]  io_mod_par_mod_module_mod_state_id,
  input         io_mod_par_mod_module_mod_sram_w_cs,
  input         io_mod_par_mod_module_mod_sram_w_en,
  input  [7:0]  io_mod_par_mod_module_mod_sram_w_addr,
  input  [63:0] io_mod_par_mod_module_mod_sram_w_data,
  input         io_mod_proc_mod_0_mat_mod_en,
  input         io_mod_proc_mod_0_mat_mod_config_id,
  input         io_mod_proc_mod_0_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_0_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_0_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_0_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_0_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_0_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_0_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_0_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_0_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_0_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_0_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_0_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_0_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_0_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_0_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_0_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_0_mat_mod_w_data,
  input         io_mod_proc_mod_0_exe_mod_en_0,
  input         io_mod_proc_mod_0_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_0_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_0_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_0_exe_mod_data_1,
  input         io_mod_proc_mod_1_mat_mod_en,
  input         io_mod_proc_mod_1_mat_mod_config_id,
  input         io_mod_proc_mod_1_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_1_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_1_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_1_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_1_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_1_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_1_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_1_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_1_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_1_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_1_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_1_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_1_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_1_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_1_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_1_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_1_mat_mod_w_data,
  input         io_mod_proc_mod_1_exe_mod_en_0,
  input         io_mod_proc_mod_1_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_1_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_1_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_1_exe_mod_data_1,
  input         io_mod_proc_mod_2_mat_mod_en,
  input         io_mod_proc_mod_2_mat_mod_config_id,
  input         io_mod_proc_mod_2_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_2_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_2_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_2_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_2_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_2_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_2_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_2_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_2_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_2_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_2_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_2_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_2_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_2_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_2_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_2_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_2_mat_mod_w_data,
  input         io_mod_proc_mod_2_exe_mod_en_0,
  input         io_mod_proc_mod_2_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_2_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_2_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_2_exe_mod_data_1,
  input         io_mod_proc_mod_3_mat_mod_en,
  input         io_mod_proc_mod_3_mat_mod_config_id,
  input         io_mod_proc_mod_3_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_3_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_3_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_3_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_3_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_3_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_3_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_3_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_3_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_3_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_3_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_3_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_3_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_3_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_3_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_3_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_3_mat_mod_w_data,
  input         io_mod_proc_mod_3_exe_mod_en_0,
  input         io_mod_proc_mod_3_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_3_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_3_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_3_exe_mod_data_1,
  input         io_mod_proc_mod_4_mat_mod_en,
  input         io_mod_proc_mod_4_mat_mod_config_id,
  input         io_mod_proc_mod_4_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_4_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_4_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_4_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_4_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_4_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_4_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_4_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_4_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_4_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_4_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_4_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_4_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_4_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_4_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_4_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_4_mat_mod_w_data,
  input         io_mod_proc_mod_4_exe_mod_en_0,
  input         io_mod_proc_mod_4_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_4_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_4_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_4_exe_mod_data_1,
  input         io_mod_proc_mod_5_mat_mod_en,
  input         io_mod_proc_mod_5_mat_mod_config_id,
  input         io_mod_proc_mod_5_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_5_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_5_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_5_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_5_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_5_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_5_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_5_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_5_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_5_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_5_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_5_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_5_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_5_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_5_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_5_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_5_mat_mod_w_data,
  input         io_mod_proc_mod_5_exe_mod_en_0,
  input         io_mod_proc_mod_5_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_5_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_5_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_5_exe_mod_data_1,
  input         io_mod_proc_mod_6_mat_mod_en,
  input         io_mod_proc_mod_6_mat_mod_config_id,
  input         io_mod_proc_mod_6_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_6_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_6_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_6_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_6_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_6_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_6_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_6_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_6_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_6_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_6_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_6_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_6_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_6_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_6_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_6_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_6_mat_mod_w_data,
  input         io_mod_proc_mod_6_exe_mod_en_0,
  input         io_mod_proc_mod_6_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_6_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_6_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_6_exe_mod_data_1,
  input         io_mod_proc_mod_7_mat_mod_en,
  input         io_mod_proc_mod_7_mat_mod_config_id,
  input         io_mod_proc_mod_7_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_7_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_7_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_7_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_7_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_7_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_7_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_7_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_7_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_7_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_7_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_7_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_7_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_7_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_7_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_7_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_7_mat_mod_w_data,
  input         io_mod_proc_mod_7_exe_mod_en_0,
  input         io_mod_proc_mod_7_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_7_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_7_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_7_exe_mod_data_1,
  input         io_mod_proc_mod_8_mat_mod_en,
  input         io_mod_proc_mod_8_mat_mod_config_id,
  input         io_mod_proc_mod_8_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_8_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_8_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_8_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_8_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_8_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_8_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_8_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_8_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_8_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_8_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_8_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_8_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_8_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_8_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_8_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_8_mat_mod_w_data,
  input         io_mod_proc_mod_8_exe_mod_en_0,
  input         io_mod_proc_mod_8_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_8_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_8_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_8_exe_mod_data_1,
  input         io_mod_proc_mod_9_mat_mod_en,
  input         io_mod_proc_mod_9_mat_mod_config_id,
  input         io_mod_proc_mod_9_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_9_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_9_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_9_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_9_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_9_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_9_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_9_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_9_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_9_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_9_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_9_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_9_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_9_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_9_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_9_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_9_mat_mod_w_data,
  input         io_mod_proc_mod_9_exe_mod_en_0,
  input         io_mod_proc_mod_9_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_9_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_9_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_9_exe_mod_data_1,
  input         io_mod_proc_mod_10_mat_mod_en,
  input         io_mod_proc_mod_10_mat_mod_config_id,
  input         io_mod_proc_mod_10_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_10_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_10_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_10_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_10_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_10_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_10_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_10_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_10_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_10_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_10_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_10_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_10_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_10_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_10_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_10_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_10_mat_mod_w_data,
  input         io_mod_proc_mod_10_exe_mod_en_0,
  input         io_mod_proc_mod_10_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_10_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_10_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_10_exe_mod_data_1,
  input         io_mod_proc_mod_11_mat_mod_en,
  input         io_mod_proc_mod_11_mat_mod_config_id,
  input         io_mod_proc_mod_11_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_11_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_11_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_11_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_11_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_11_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_11_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_11_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_11_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_11_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_11_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_11_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_11_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_11_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_11_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_11_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_11_mat_mod_w_data,
  input         io_mod_proc_mod_11_exe_mod_en_0,
  input         io_mod_proc_mod_11_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_11_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_11_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_11_exe_mod_data_1
);
  wire  init_clock; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_0; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_1; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_2; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_3; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_4; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_5; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_6; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_7; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_8; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_9; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_10; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_11; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_12; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_13; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_14; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_15; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_16; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_17; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_18; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_19; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_20; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_21; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_22; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_23; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_24; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_25; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_26; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_27; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_28; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_29; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_30; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_31; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_32; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_33; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_34; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_35; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_36; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_37; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_38; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_39; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_40; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_41; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_42; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_43; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_44; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_45; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_46; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_47; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_48; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_49; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_50; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_51; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_52; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_53; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_54; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_55; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_56; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_57; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_58; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_59; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_60; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_61; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_62; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_63; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_64; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_65; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_66; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_67; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_68; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_69; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_70; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_71; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_72; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_73; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_74; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_75; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_76; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_77; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_78; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_79; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_80; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_81; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_82; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_83; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_84; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_85; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_86; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_87; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_88; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_89; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_90; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_91; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_92; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_93; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_94; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_95; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_96; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_97; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_98; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_99; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_100; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_101; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_102; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_103; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_104; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_105; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_106; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_107; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_108; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_109; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_110; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_111; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_112; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_113; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_114; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_115; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_116; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_117; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_118; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_119; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_120; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_121; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_122; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_123; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_124; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_125; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_126; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_127; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_128; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_129; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_130; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_131; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_132; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_133; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_134; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_135; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_136; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_137; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_138; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_139; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_140; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_141; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_142; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_143; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_144; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_145; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_146; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_147; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_148; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_149; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_150; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_151; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_152; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_153; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_154; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_155; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_156; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_157; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_158; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_159; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_160; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_161; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_162; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_163; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_164; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_165; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_166; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_167; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_168; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_169; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_170; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_171; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_172; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_173; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_174; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_175; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_176; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_177; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_178; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_179; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_180; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_181; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_182; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_183; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_184; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_185; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_186; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_187; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_188; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_189; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_190; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_191; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_0; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_1; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_2; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_3; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_4; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_5; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_6; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_7; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_8; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_9; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_10; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_11; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_12; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_13; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_14; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_15; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_16; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_17; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_18; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_19; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_20; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_21; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_22; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_23; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_24; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_25; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_26; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_27; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_28; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_29; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_30; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_31; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_32; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_33; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_34; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_35; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_36; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_37; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_38; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_39; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_40; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_41; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_42; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_43; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_44; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_45; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_46; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_47; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_48; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_49; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_50; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_51; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_52; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_53; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_54; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_55; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_56; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_57; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_58; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_59; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_60; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_61; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_62; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_63; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_64; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_65; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_66; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_67; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_68; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_69; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_70; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_71; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_72; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_73; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_74; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_75; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_76; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_77; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_78; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_79; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_80; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_81; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_82; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_83; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_84; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_85; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_86; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_87; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_88; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_89; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_90; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_91; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_92; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_93; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_94; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_95; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_96; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_97; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_98; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_99; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_100; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_101; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_102; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_103; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_104; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_105; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_106; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_107; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_108; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_109; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_110; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_111; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_112; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_113; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_114; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_115; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_116; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_117; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_118; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_119; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_120; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_121; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_122; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_123; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_124; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_125; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_126; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_127; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_128; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_129; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_130; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_131; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_132; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_133; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_134; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_135; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_136; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_137; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_138; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_139; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_140; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_141; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_142; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_143; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_144; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_145; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_146; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_147; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_148; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_149; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_150; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_151; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_152; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_153; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_154; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_155; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_156; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_157; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_158; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_159; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_160; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_161; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_162; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_163; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_164; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_165; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_166; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_167; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_168; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_169; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_170; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_171; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_172; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_173; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_174; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_175; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_176; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_177; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_178; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_179; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_180; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_181; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_182; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_183; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_184; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_185; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_186; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_187; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_188; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_189; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_190; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_191; // @[pisa.scala 19:22]
  wire  PAR_clock; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_0; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_1; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_2; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_3; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_4; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_5; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_6; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_7; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_8; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_9; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_10; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_11; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_12; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_13; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_14; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_15; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_16; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_17; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_18; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_19; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_20; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_21; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_22; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_23; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_24; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_25; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_26; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_27; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_28; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_29; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_30; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_31; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_32; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_33; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_34; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_35; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_36; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_37; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_38; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_39; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_40; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_41; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_42; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_43; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_44; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_45; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_46; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_47; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_48; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_49; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_50; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_51; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_52; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_53; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_54; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_55; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_56; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_57; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_58; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_59; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_60; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_61; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_62; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_63; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_64; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_65; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_66; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_67; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_68; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_69; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_70; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_71; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_72; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_73; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_74; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_75; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_76; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_77; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_78; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_79; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_80; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_81; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_82; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_83; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_84; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_85; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_86; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_87; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_88; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_89; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_90; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_91; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_92; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_93; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_94; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_95; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_96; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_97; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_98; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_99; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_100; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_101; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_102; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_103; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_104; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_105; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_106; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_107; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_108; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_109; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_110; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_111; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_112; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_113; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_114; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_115; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_116; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_117; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_118; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_119; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_120; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_121; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_122; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_123; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_124; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_125; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_126; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_127; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_128; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_129; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_130; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_131; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_132; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_133; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_134; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_135; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_136; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_137; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_138; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_139; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_140; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_141; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_142; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_143; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_144; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_145; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_146; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_147; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_148; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_149; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_150; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_151; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_152; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_153; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_154; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_155; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_156; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_157; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_158; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_159; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_160; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_161; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_162; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_163; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_164; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_165; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_166; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_167; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_168; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_169; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_170; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_171; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_172; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_173; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_174; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_175; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_176; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_177; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_178; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_179; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_180; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_181; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_182; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_183; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_184; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_185; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_186; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_187; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_188; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_189; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_190; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_191; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_0; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_1; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_2; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_3; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_4; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_5; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_6; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_7; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_8; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_9; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_10; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_11; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_12; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_13; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_14; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_15; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_16; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_17; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_18; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_19; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_20; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_21; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_22; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_23; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_24; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_25; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_26; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_27; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_28; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_29; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_30; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_31; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_32; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_33; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_34; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_35; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_36; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_37; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_38; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_39; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_40; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_41; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_42; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_43; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_44; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_45; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_46; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_47; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_48; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_49; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_50; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_51; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_52; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_53; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_54; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_55; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_56; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_57; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_58; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_59; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_60; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_61; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_62; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_63; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_64; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_65; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_66; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_67; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_68; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_69; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_70; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_71; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_72; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_73; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_74; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_75; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_76; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_77; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_78; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_79; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_80; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_81; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_82; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_83; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_84; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_85; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_86; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_87; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_88; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_89; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_90; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_91; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_92; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_93; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_94; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_95; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_96; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_97; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_98; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_99; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_100; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_101; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_102; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_103; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_104; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_105; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_106; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_107; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_108; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_109; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_110; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_111; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_112; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_113; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_114; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_115; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_116; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_117; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_118; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_119; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_120; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_121; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_122; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_123; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_124; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_125; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_126; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_127; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_128; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_129; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_130; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_131; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_132; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_133; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_134; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_135; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_136; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_137; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_138; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_139; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_140; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_141; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_142; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_143; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_144; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_145; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_146; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_147; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_148; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_149; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_150; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_151; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_152; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_153; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_154; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_155; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_156; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_157; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_158; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_159; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_160; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_161; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_162; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_163; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_164; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_165; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_166; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_167; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_168; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_169; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_170; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_171; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_172; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_173; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_174; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_175; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_176; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_177; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_178; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_179; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_180; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_181; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_182; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_183; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_184; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_185; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_186; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_187; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_188; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_189; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_190; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_191; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_192; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_193; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_194; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_195; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_196; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_197; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_198; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_199; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_200; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_201; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_202; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_203; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_204; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_205; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_206; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_207; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_208; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_209; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_210; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_211; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_212; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_213; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_214; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_215; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_216; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_217; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_218; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_219; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_220; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_221; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_222; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_223; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_224; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_225; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_226; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_227; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_228; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_229; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_230; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_231; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_232; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_233; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_234; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_235; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_236; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_237; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_238; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_239; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_240; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_241; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_242; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_243; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_244; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_245; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_246; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_247; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_248; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_249; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_250; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_251; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_252; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_253; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_254; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_255; // @[pisa.scala 23:21]
  wire [3:0] PAR_io_pipe_phv_out_next_processor_id; // @[pisa.scala 23:21]
  wire  PAR_io_pipe_phv_out_next_config_id; // @[pisa.scala 23:21]
  wire  PAR_io_mod_en; // @[pisa.scala 23:21]
  wire  PAR_io_mod_last_mau_id_mod; // @[pisa.scala 23:21]
  wire [3:0] PAR_io_mod_last_mau_id; // @[pisa.scala 23:21]
  wire [2:0] PAR_io_mod_cs; // @[pisa.scala 23:21]
  wire  PAR_io_mod_module_mod_state_id_mod; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_mod_module_mod_state_id; // @[pisa.scala 23:21]
  wire  PAR_io_mod_module_mod_sram_w_cs; // @[pisa.scala 23:21]
  wire  PAR_io_mod_module_mod_sram_w_en; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_mod_module_mod_sram_w_addr; // @[pisa.scala 23:21]
  wire [63:0] PAR_io_mod_module_mod_sram_w_data; // @[pisa.scala 23:21]
  wire  proc_0_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_160; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_161; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_162; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_163; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_164; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_165; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_166; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_167; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_168; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_169; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_170; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_171; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_172; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_173; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_174; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_175; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_176; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_177; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_178; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_179; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_180; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_181; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_182; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_183; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_184; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_185; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_186; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_187; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_188; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_189; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_190; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_191; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_192; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_193; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_194; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_195; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_196; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_197; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_198; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_199; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_200; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_201; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_202; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_203; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_204; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_205; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_206; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_207; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_208; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_209; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_210; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_211; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_212; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_213; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_214; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_215; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_216; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_217; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_218; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_219; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_220; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_221; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_222; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_223; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_224; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_225; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_226; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_227; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_228; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_229; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_230; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_231; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_232; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_233; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_234; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_235; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_236; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_237; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_238; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_239; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_240; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_241; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_242; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_243; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_244; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_245; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_246; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_247; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_248; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_249; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_250; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_251; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_252; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_253; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_254; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_255; // @[pisa.scala 28:25]
  wire [3:0] proc_0_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_0_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_0_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_160; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_161; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_162; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_163; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_164; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_165; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_166; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_167; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_168; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_169; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_170; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_171; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_172; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_173; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_174; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_175; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_176; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_177; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_178; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_179; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_180; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_181; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_182; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_183; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_184; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_185; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_186; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_187; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_188; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_189; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_190; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_191; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_192; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_193; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_194; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_195; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_196; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_197; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_198; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_199; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_200; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_201; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_202; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_203; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_204; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_205; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_206; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_207; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_208; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_209; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_210; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_211; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_212; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_213; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_214; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_215; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_216; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_217; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_218; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_219; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_220; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_221; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_222; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_223; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_224; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_225; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_226; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_227; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_228; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_229; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_230; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_231; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_232; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_233; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_234; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_235; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_236; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_237; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_238; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_239; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_240; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_241; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_242; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_243; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_244; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_245; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_246; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_247; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_248; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_249; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_250; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_251; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_252; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_253; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_254; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_255; // @[pisa.scala 28:25]
  wire [3:0] proc_0_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_0_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_0_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_0_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_0_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_0_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_0_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_0_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_0_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_0_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_0_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_0_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_0_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_0_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_0_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_0_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_0_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_0_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_0_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_0_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_0_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_0_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_0_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_0_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  wire  proc_1_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_160; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_161; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_162; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_163; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_164; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_165; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_166; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_167; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_168; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_169; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_170; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_171; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_172; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_173; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_174; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_175; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_176; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_177; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_178; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_179; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_180; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_181; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_182; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_183; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_184; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_185; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_186; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_187; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_188; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_189; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_190; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_191; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_192; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_193; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_194; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_195; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_196; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_197; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_198; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_199; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_200; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_201; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_202; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_203; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_204; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_205; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_206; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_207; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_208; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_209; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_210; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_211; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_212; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_213; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_214; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_215; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_216; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_217; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_218; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_219; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_220; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_221; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_222; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_223; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_224; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_225; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_226; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_227; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_228; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_229; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_230; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_231; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_232; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_233; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_234; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_235; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_236; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_237; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_238; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_239; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_240; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_241; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_242; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_243; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_244; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_245; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_246; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_247; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_248; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_249; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_250; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_251; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_252; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_253; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_254; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_255; // @[pisa.scala 28:25]
  wire [3:0] proc_1_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_1_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_1_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_160; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_161; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_162; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_163; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_164; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_165; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_166; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_167; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_168; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_169; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_170; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_171; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_172; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_173; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_174; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_175; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_176; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_177; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_178; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_179; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_180; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_181; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_182; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_183; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_184; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_185; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_186; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_187; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_188; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_189; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_190; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_191; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_192; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_193; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_194; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_195; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_196; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_197; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_198; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_199; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_200; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_201; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_202; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_203; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_204; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_205; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_206; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_207; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_208; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_209; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_210; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_211; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_212; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_213; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_214; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_215; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_216; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_217; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_218; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_219; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_220; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_221; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_222; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_223; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_224; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_225; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_226; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_227; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_228; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_229; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_230; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_231; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_232; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_233; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_234; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_235; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_236; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_237; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_238; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_239; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_240; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_241; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_242; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_243; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_244; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_245; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_246; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_247; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_248; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_249; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_250; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_251; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_252; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_253; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_254; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_255; // @[pisa.scala 28:25]
  wire [3:0] proc_1_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_1_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_1_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_1_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_1_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_1_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_1_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_1_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_1_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_1_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_1_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_1_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_1_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_1_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_1_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_1_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_1_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_1_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_1_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_1_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_1_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_1_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_1_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_1_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  wire  proc_2_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_160; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_161; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_162; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_163; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_164; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_165; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_166; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_167; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_168; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_169; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_170; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_171; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_172; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_173; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_174; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_175; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_176; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_177; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_178; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_179; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_180; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_181; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_182; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_183; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_184; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_185; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_186; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_187; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_188; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_189; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_190; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_191; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_192; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_193; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_194; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_195; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_196; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_197; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_198; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_199; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_200; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_201; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_202; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_203; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_204; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_205; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_206; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_207; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_208; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_209; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_210; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_211; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_212; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_213; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_214; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_215; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_216; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_217; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_218; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_219; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_220; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_221; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_222; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_223; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_224; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_225; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_226; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_227; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_228; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_229; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_230; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_231; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_232; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_233; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_234; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_235; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_236; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_237; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_238; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_239; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_240; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_241; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_242; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_243; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_244; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_245; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_246; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_247; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_248; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_249; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_250; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_251; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_252; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_253; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_254; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_255; // @[pisa.scala 28:25]
  wire [3:0] proc_2_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_2_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_2_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_160; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_161; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_162; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_163; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_164; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_165; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_166; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_167; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_168; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_169; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_170; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_171; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_172; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_173; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_174; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_175; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_176; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_177; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_178; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_179; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_180; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_181; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_182; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_183; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_184; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_185; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_186; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_187; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_188; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_189; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_190; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_191; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_192; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_193; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_194; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_195; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_196; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_197; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_198; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_199; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_200; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_201; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_202; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_203; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_204; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_205; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_206; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_207; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_208; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_209; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_210; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_211; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_212; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_213; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_214; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_215; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_216; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_217; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_218; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_219; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_220; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_221; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_222; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_223; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_224; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_225; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_226; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_227; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_228; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_229; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_230; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_231; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_232; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_233; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_234; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_235; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_236; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_237; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_238; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_239; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_240; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_241; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_242; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_243; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_244; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_245; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_246; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_247; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_248; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_249; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_250; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_251; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_252; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_253; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_254; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_255; // @[pisa.scala 28:25]
  wire [3:0] proc_2_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_2_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_2_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_2_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_2_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_2_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_2_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_2_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_2_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_2_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_2_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_2_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_2_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_2_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_2_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_2_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_2_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_2_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_2_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_2_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_2_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_2_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_2_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_2_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  wire  proc_3_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_160; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_161; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_162; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_163; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_164; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_165; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_166; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_167; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_168; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_169; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_170; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_171; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_172; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_173; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_174; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_175; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_176; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_177; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_178; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_179; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_180; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_181; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_182; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_183; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_184; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_185; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_186; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_187; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_188; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_189; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_190; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_191; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_192; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_193; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_194; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_195; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_196; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_197; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_198; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_199; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_200; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_201; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_202; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_203; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_204; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_205; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_206; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_207; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_208; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_209; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_210; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_211; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_212; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_213; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_214; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_215; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_216; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_217; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_218; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_219; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_220; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_221; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_222; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_223; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_224; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_225; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_226; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_227; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_228; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_229; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_230; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_231; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_232; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_233; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_234; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_235; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_236; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_237; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_238; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_239; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_240; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_241; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_242; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_243; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_244; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_245; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_246; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_247; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_248; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_249; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_250; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_251; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_252; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_253; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_254; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_255; // @[pisa.scala 28:25]
  wire [3:0] proc_3_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_3_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_3_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_160; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_161; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_162; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_163; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_164; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_165; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_166; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_167; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_168; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_169; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_170; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_171; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_172; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_173; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_174; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_175; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_176; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_177; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_178; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_179; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_180; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_181; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_182; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_183; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_184; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_185; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_186; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_187; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_188; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_189; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_190; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_191; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_192; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_193; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_194; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_195; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_196; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_197; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_198; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_199; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_200; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_201; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_202; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_203; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_204; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_205; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_206; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_207; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_208; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_209; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_210; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_211; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_212; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_213; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_214; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_215; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_216; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_217; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_218; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_219; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_220; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_221; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_222; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_223; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_224; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_225; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_226; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_227; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_228; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_229; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_230; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_231; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_232; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_233; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_234; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_235; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_236; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_237; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_238; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_239; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_240; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_241; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_242; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_243; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_244; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_245; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_246; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_247; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_248; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_249; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_250; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_251; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_252; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_253; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_254; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_255; // @[pisa.scala 28:25]
  wire [3:0] proc_3_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_3_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_3_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_3_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_3_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_3_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_3_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_3_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_3_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_3_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_3_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_3_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_3_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_3_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_3_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_3_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_3_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_3_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_3_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_3_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_3_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_3_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_3_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_3_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  wire  proc_4_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_160; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_161; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_162; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_163; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_164; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_165; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_166; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_167; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_168; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_169; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_170; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_171; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_172; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_173; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_174; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_175; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_176; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_177; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_178; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_179; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_180; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_181; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_182; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_183; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_184; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_185; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_186; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_187; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_188; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_189; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_190; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_191; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_192; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_193; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_194; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_195; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_196; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_197; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_198; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_199; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_200; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_201; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_202; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_203; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_204; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_205; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_206; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_207; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_208; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_209; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_210; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_211; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_212; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_213; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_214; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_215; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_216; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_217; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_218; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_219; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_220; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_221; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_222; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_223; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_224; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_225; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_226; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_227; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_228; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_229; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_230; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_231; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_232; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_233; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_234; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_235; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_236; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_237; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_238; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_239; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_240; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_241; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_242; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_243; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_244; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_245; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_246; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_247; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_248; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_249; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_250; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_251; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_252; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_253; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_254; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_255; // @[pisa.scala 28:25]
  wire [3:0] proc_4_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_4_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_4_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_160; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_161; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_162; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_163; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_164; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_165; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_166; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_167; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_168; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_169; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_170; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_171; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_172; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_173; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_174; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_175; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_176; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_177; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_178; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_179; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_180; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_181; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_182; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_183; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_184; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_185; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_186; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_187; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_188; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_189; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_190; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_191; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_192; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_193; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_194; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_195; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_196; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_197; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_198; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_199; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_200; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_201; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_202; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_203; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_204; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_205; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_206; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_207; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_208; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_209; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_210; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_211; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_212; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_213; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_214; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_215; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_216; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_217; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_218; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_219; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_220; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_221; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_222; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_223; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_224; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_225; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_226; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_227; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_228; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_229; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_230; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_231; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_232; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_233; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_234; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_235; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_236; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_237; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_238; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_239; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_240; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_241; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_242; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_243; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_244; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_245; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_246; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_247; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_248; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_249; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_250; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_251; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_252; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_253; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_254; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_255; // @[pisa.scala 28:25]
  wire [3:0] proc_4_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_4_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_4_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_4_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_4_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_4_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_4_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_4_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_4_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_4_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_4_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_4_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_4_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_4_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_4_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_4_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_4_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_4_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_4_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_4_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_4_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_4_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_4_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_4_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  wire  proc_5_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_160; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_161; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_162; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_163; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_164; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_165; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_166; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_167; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_168; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_169; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_170; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_171; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_172; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_173; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_174; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_175; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_176; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_177; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_178; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_179; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_180; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_181; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_182; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_183; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_184; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_185; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_186; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_187; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_188; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_189; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_190; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_191; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_192; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_193; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_194; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_195; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_196; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_197; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_198; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_199; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_200; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_201; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_202; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_203; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_204; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_205; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_206; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_207; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_208; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_209; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_210; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_211; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_212; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_213; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_214; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_215; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_216; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_217; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_218; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_219; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_220; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_221; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_222; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_223; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_224; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_225; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_226; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_227; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_228; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_229; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_230; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_231; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_232; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_233; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_234; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_235; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_236; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_237; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_238; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_239; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_240; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_241; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_242; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_243; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_244; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_245; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_246; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_247; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_248; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_249; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_250; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_251; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_252; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_253; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_254; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_255; // @[pisa.scala 28:25]
  wire [3:0] proc_5_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_5_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_5_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_160; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_161; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_162; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_163; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_164; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_165; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_166; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_167; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_168; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_169; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_170; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_171; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_172; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_173; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_174; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_175; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_176; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_177; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_178; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_179; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_180; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_181; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_182; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_183; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_184; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_185; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_186; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_187; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_188; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_189; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_190; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_191; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_192; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_193; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_194; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_195; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_196; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_197; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_198; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_199; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_200; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_201; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_202; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_203; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_204; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_205; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_206; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_207; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_208; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_209; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_210; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_211; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_212; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_213; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_214; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_215; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_216; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_217; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_218; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_219; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_220; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_221; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_222; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_223; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_224; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_225; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_226; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_227; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_228; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_229; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_230; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_231; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_232; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_233; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_234; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_235; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_236; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_237; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_238; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_239; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_240; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_241; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_242; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_243; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_244; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_245; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_246; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_247; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_248; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_249; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_250; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_251; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_252; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_253; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_254; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_255; // @[pisa.scala 28:25]
  wire [3:0] proc_5_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_5_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_5_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_5_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_5_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_5_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_5_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_5_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_5_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_5_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_5_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_5_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_5_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_5_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_5_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_5_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_5_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_5_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_5_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_5_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_5_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_5_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_5_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_5_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  wire  proc_6_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_160; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_161; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_162; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_163; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_164; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_165; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_166; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_167; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_168; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_169; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_170; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_171; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_172; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_173; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_174; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_175; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_176; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_177; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_178; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_179; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_180; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_181; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_182; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_183; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_184; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_185; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_186; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_187; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_188; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_189; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_190; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_191; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_192; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_193; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_194; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_195; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_196; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_197; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_198; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_199; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_200; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_201; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_202; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_203; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_204; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_205; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_206; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_207; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_208; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_209; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_210; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_211; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_212; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_213; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_214; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_215; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_216; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_217; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_218; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_219; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_220; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_221; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_222; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_223; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_224; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_225; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_226; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_227; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_228; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_229; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_230; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_231; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_232; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_233; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_234; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_235; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_236; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_237; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_238; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_239; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_240; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_241; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_242; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_243; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_244; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_245; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_246; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_247; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_248; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_249; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_250; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_251; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_252; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_253; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_254; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_255; // @[pisa.scala 28:25]
  wire [3:0] proc_6_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_6_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_6_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_160; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_161; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_162; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_163; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_164; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_165; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_166; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_167; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_168; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_169; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_170; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_171; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_172; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_173; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_174; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_175; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_176; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_177; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_178; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_179; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_180; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_181; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_182; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_183; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_184; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_185; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_186; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_187; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_188; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_189; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_190; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_191; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_192; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_193; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_194; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_195; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_196; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_197; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_198; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_199; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_200; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_201; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_202; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_203; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_204; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_205; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_206; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_207; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_208; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_209; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_210; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_211; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_212; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_213; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_214; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_215; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_216; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_217; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_218; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_219; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_220; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_221; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_222; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_223; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_224; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_225; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_226; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_227; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_228; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_229; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_230; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_231; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_232; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_233; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_234; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_235; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_236; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_237; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_238; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_239; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_240; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_241; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_242; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_243; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_244; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_245; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_246; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_247; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_248; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_249; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_250; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_251; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_252; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_253; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_254; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_255; // @[pisa.scala 28:25]
  wire [3:0] proc_6_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_6_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_6_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_6_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_6_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_6_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_6_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_6_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_6_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_6_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_6_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_6_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_6_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_6_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_6_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_6_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_6_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_6_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_6_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_6_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_6_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_6_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_6_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_6_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  wire  proc_7_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_160; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_161; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_162; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_163; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_164; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_165; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_166; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_167; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_168; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_169; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_170; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_171; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_172; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_173; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_174; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_175; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_176; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_177; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_178; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_179; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_180; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_181; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_182; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_183; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_184; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_185; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_186; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_187; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_188; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_189; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_190; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_191; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_192; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_193; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_194; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_195; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_196; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_197; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_198; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_199; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_200; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_201; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_202; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_203; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_204; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_205; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_206; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_207; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_208; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_209; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_210; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_211; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_212; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_213; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_214; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_215; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_216; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_217; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_218; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_219; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_220; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_221; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_222; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_223; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_224; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_225; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_226; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_227; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_228; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_229; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_230; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_231; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_232; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_233; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_234; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_235; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_236; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_237; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_238; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_239; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_240; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_241; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_242; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_243; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_244; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_245; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_246; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_247; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_248; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_249; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_250; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_251; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_252; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_253; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_254; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_255; // @[pisa.scala 28:25]
  wire [3:0] proc_7_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_7_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_7_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_160; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_161; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_162; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_163; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_164; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_165; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_166; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_167; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_168; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_169; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_170; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_171; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_172; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_173; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_174; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_175; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_176; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_177; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_178; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_179; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_180; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_181; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_182; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_183; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_184; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_185; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_186; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_187; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_188; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_189; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_190; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_191; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_192; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_193; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_194; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_195; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_196; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_197; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_198; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_199; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_200; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_201; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_202; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_203; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_204; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_205; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_206; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_207; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_208; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_209; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_210; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_211; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_212; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_213; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_214; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_215; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_216; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_217; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_218; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_219; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_220; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_221; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_222; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_223; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_224; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_225; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_226; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_227; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_228; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_229; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_230; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_231; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_232; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_233; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_234; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_235; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_236; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_237; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_238; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_239; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_240; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_241; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_242; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_243; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_244; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_245; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_246; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_247; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_248; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_249; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_250; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_251; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_252; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_253; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_254; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_255; // @[pisa.scala 28:25]
  wire [3:0] proc_7_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_7_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_7_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_7_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_7_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_7_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_7_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_7_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_7_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_7_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_7_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_7_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_7_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_7_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_7_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_7_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_7_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_7_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_7_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_7_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_7_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_7_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_7_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_7_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  wire  proc_8_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_160; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_161; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_162; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_163; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_164; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_165; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_166; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_167; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_168; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_169; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_170; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_171; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_172; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_173; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_174; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_175; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_176; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_177; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_178; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_179; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_180; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_181; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_182; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_183; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_184; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_185; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_186; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_187; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_188; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_189; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_190; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_191; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_192; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_193; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_194; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_195; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_196; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_197; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_198; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_199; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_200; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_201; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_202; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_203; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_204; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_205; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_206; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_207; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_208; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_209; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_210; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_211; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_212; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_213; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_214; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_215; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_216; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_217; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_218; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_219; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_220; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_221; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_222; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_223; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_224; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_225; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_226; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_227; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_228; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_229; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_230; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_231; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_232; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_233; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_234; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_235; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_236; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_237; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_238; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_239; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_240; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_241; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_242; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_243; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_244; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_245; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_246; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_247; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_248; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_249; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_250; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_251; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_252; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_253; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_254; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_255; // @[pisa.scala 28:25]
  wire [3:0] proc_8_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_8_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_8_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_160; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_161; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_162; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_163; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_164; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_165; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_166; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_167; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_168; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_169; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_170; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_171; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_172; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_173; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_174; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_175; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_176; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_177; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_178; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_179; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_180; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_181; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_182; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_183; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_184; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_185; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_186; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_187; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_188; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_189; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_190; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_191; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_192; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_193; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_194; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_195; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_196; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_197; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_198; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_199; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_200; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_201; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_202; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_203; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_204; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_205; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_206; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_207; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_208; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_209; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_210; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_211; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_212; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_213; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_214; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_215; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_216; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_217; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_218; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_219; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_220; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_221; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_222; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_223; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_224; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_225; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_226; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_227; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_228; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_229; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_230; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_231; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_232; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_233; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_234; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_235; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_236; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_237; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_238; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_239; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_240; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_241; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_242; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_243; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_244; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_245; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_246; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_247; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_248; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_249; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_250; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_251; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_252; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_253; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_254; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_255; // @[pisa.scala 28:25]
  wire [3:0] proc_8_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_8_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_8_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_8_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_8_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_8_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_8_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_8_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_8_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_8_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_8_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_8_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_8_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_8_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_8_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_8_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_8_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_8_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_8_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_8_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_8_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_8_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_8_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_8_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  wire  proc_9_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_160; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_161; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_162; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_163; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_164; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_165; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_166; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_167; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_168; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_169; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_170; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_171; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_172; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_173; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_174; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_175; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_176; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_177; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_178; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_179; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_180; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_181; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_182; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_183; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_184; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_185; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_186; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_187; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_188; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_189; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_190; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_191; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_192; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_193; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_194; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_195; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_196; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_197; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_198; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_199; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_200; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_201; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_202; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_203; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_204; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_205; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_206; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_207; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_208; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_209; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_210; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_211; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_212; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_213; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_214; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_215; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_216; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_217; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_218; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_219; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_220; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_221; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_222; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_223; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_224; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_225; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_226; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_227; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_228; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_229; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_230; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_231; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_232; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_233; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_234; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_235; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_236; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_237; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_238; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_239; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_240; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_241; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_242; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_243; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_244; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_245; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_246; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_247; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_248; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_249; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_250; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_251; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_252; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_253; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_254; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_255; // @[pisa.scala 28:25]
  wire [3:0] proc_9_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_9_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_9_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_160; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_161; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_162; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_163; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_164; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_165; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_166; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_167; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_168; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_169; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_170; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_171; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_172; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_173; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_174; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_175; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_176; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_177; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_178; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_179; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_180; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_181; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_182; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_183; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_184; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_185; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_186; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_187; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_188; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_189; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_190; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_191; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_192; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_193; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_194; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_195; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_196; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_197; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_198; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_199; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_200; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_201; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_202; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_203; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_204; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_205; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_206; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_207; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_208; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_209; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_210; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_211; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_212; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_213; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_214; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_215; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_216; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_217; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_218; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_219; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_220; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_221; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_222; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_223; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_224; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_225; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_226; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_227; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_228; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_229; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_230; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_231; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_232; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_233; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_234; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_235; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_236; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_237; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_238; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_239; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_240; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_241; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_242; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_243; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_244; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_245; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_246; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_247; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_248; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_249; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_250; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_251; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_252; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_253; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_254; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_255; // @[pisa.scala 28:25]
  wire [3:0] proc_9_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_9_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_9_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_9_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_9_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_9_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_9_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_9_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_9_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_9_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_9_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_9_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_9_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_9_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_9_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_9_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_9_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_9_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_9_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_9_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_9_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_9_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_9_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_9_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  wire  proc_10_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_160; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_161; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_162; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_163; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_164; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_165; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_166; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_167; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_168; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_169; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_170; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_171; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_172; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_173; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_174; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_175; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_176; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_177; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_178; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_179; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_180; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_181; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_182; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_183; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_184; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_185; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_186; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_187; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_188; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_189; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_190; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_191; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_192; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_193; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_194; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_195; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_196; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_197; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_198; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_199; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_200; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_201; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_202; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_203; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_204; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_205; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_206; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_207; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_208; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_209; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_210; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_211; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_212; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_213; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_214; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_215; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_216; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_217; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_218; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_219; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_220; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_221; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_222; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_223; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_224; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_225; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_226; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_227; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_228; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_229; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_230; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_231; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_232; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_233; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_234; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_235; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_236; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_237; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_238; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_239; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_240; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_241; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_242; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_243; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_244; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_245; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_246; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_247; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_248; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_249; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_250; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_251; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_252; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_253; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_254; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_255; // @[pisa.scala 28:25]
  wire [3:0] proc_10_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_10_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_10_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_160; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_161; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_162; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_163; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_164; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_165; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_166; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_167; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_168; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_169; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_170; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_171; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_172; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_173; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_174; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_175; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_176; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_177; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_178; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_179; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_180; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_181; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_182; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_183; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_184; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_185; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_186; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_187; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_188; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_189; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_190; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_191; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_192; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_193; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_194; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_195; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_196; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_197; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_198; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_199; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_200; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_201; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_202; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_203; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_204; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_205; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_206; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_207; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_208; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_209; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_210; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_211; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_212; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_213; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_214; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_215; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_216; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_217; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_218; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_219; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_220; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_221; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_222; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_223; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_224; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_225; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_226; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_227; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_228; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_229; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_230; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_231; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_232; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_233; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_234; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_235; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_236; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_237; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_238; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_239; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_240; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_241; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_242; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_243; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_244; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_245; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_246; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_247; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_248; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_249; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_250; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_251; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_252; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_253; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_254; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_255; // @[pisa.scala 28:25]
  wire [3:0] proc_10_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_10_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_10_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_10_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_10_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_10_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_10_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_10_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_10_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_10_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_10_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_10_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_10_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_10_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_10_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_10_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_10_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_10_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_10_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_10_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_10_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_10_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_10_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_10_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  wire  proc_11_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_160; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_161; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_162; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_163; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_164; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_165; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_166; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_167; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_168; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_169; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_170; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_171; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_172; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_173; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_174; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_175; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_176; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_177; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_178; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_179; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_180; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_181; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_182; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_183; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_184; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_185; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_186; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_187; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_188; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_189; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_190; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_191; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_192; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_193; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_194; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_195; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_196; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_197; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_198; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_199; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_200; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_201; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_202; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_203; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_204; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_205; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_206; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_207; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_208; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_209; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_210; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_211; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_212; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_213; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_214; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_215; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_216; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_217; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_218; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_219; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_220; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_221; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_222; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_223; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_224; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_225; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_226; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_227; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_228; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_229; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_230; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_231; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_232; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_233; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_234; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_235; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_236; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_237; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_238; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_239; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_240; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_241; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_242; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_243; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_244; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_245; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_246; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_247; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_248; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_249; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_250; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_251; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_252; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_253; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_254; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_255; // @[pisa.scala 28:25]
  wire [3:0] proc_11_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_11_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_11_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_160; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_161; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_162; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_163; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_164; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_165; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_166; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_167; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_168; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_169; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_170; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_171; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_172; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_173; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_174; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_175; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_176; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_177; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_178; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_179; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_180; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_181; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_182; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_183; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_184; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_185; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_186; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_187; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_188; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_189; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_190; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_191; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_192; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_193; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_194; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_195; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_196; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_197; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_198; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_199; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_200; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_201; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_202; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_203; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_204; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_205; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_206; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_207; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_208; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_209; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_210; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_211; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_212; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_213; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_214; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_215; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_216; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_217; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_218; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_219; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_220; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_221; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_222; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_223; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_224; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_225; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_226; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_227; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_228; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_229; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_230; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_231; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_232; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_233; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_234; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_235; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_236; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_237; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_238; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_239; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_240; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_241; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_242; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_243; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_244; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_245; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_246; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_247; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_248; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_249; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_250; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_251; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_252; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_253; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_254; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_255; // @[pisa.scala 28:25]
  wire [3:0] proc_11_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_11_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_11_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_11_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_11_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_11_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_11_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_11_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_11_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_11_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_11_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_11_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_11_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_11_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_11_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_11_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_11_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_11_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_11_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_11_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_11_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_11_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_11_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_11_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  Initializer init ( // @[pisa.scala 19:22]
    .clock(init_clock),
    .io_pipe_phv_in_data_0(init_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(init_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(init_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(init_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(init_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(init_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(init_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(init_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(init_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(init_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(init_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(init_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(init_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(init_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(init_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(init_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(init_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(init_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(init_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(init_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(init_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(init_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(init_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(init_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(init_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(init_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(init_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(init_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(init_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(init_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(init_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(init_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(init_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(init_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(init_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(init_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(init_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(init_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(init_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(init_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(init_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(init_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(init_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(init_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(init_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(init_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(init_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(init_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(init_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(init_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(init_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(init_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(init_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(init_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(init_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(init_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(init_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(init_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(init_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(init_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(init_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(init_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(init_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(init_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(init_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(init_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(init_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(init_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(init_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(init_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(init_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(init_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(init_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(init_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(init_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(init_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(init_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(init_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(init_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(init_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(init_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(init_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(init_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(init_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(init_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(init_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(init_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(init_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(init_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(init_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(init_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(init_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(init_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(init_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(init_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(init_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(init_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(init_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(init_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(init_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(init_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(init_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(init_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(init_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(init_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(init_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(init_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(init_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(init_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(init_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(init_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(init_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(init_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(init_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(init_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(init_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(init_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(init_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(init_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(init_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(init_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(init_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(init_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(init_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(init_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(init_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(init_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(init_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(init_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(init_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(init_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(init_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(init_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(init_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(init_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(init_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(init_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(init_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(init_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(init_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(init_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(init_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(init_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(init_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(init_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(init_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(init_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(init_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(init_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(init_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(init_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(init_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(init_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(init_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(init_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(init_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(init_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(init_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(init_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(init_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(init_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(init_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(init_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(init_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(init_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(init_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(init_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(init_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(init_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(init_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(init_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(init_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(init_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(init_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(init_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(init_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(init_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(init_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(init_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(init_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(init_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(init_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(init_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(init_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(init_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(init_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(init_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(init_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(init_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(init_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(init_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(init_io_pipe_phv_in_data_191),
    .io_pipe_phv_out_data_0(init_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(init_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(init_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(init_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(init_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(init_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(init_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(init_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(init_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(init_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(init_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(init_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(init_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(init_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(init_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(init_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(init_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(init_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(init_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(init_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(init_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(init_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(init_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(init_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(init_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(init_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(init_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(init_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(init_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(init_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(init_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(init_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(init_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(init_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(init_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(init_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(init_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(init_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(init_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(init_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(init_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(init_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(init_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(init_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(init_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(init_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(init_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(init_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(init_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(init_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(init_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(init_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(init_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(init_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(init_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(init_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(init_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(init_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(init_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(init_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(init_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(init_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(init_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(init_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(init_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(init_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(init_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(init_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(init_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(init_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(init_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(init_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(init_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(init_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(init_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(init_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(init_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(init_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(init_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(init_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(init_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(init_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(init_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(init_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(init_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(init_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(init_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(init_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(init_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(init_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(init_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(init_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(init_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(init_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(init_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(init_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(init_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(init_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(init_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(init_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(init_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(init_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(init_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(init_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(init_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(init_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(init_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(init_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(init_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(init_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(init_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(init_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(init_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(init_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(init_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(init_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(init_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(init_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(init_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(init_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(init_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(init_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(init_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(init_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(init_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(init_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(init_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(init_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(init_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(init_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(init_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(init_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(init_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(init_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(init_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(init_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(init_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(init_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(init_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(init_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(init_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(init_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(init_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(init_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(init_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(init_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(init_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(init_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(init_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(init_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(init_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(init_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(init_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(init_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(init_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(init_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(init_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(init_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(init_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(init_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(init_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(init_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(init_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(init_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(init_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(init_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(init_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(init_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(init_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(init_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(init_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(init_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(init_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(init_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(init_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(init_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(init_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(init_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(init_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(init_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(init_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(init_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(init_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(init_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(init_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(init_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(init_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(init_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(init_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(init_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(init_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(init_io_pipe_phv_out_data_191)
  );
  ParserPISA PAR ( // @[pisa.scala 23:21]
    .clock(PAR_clock),
    .io_pipe_phv_in_data_0(PAR_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(PAR_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(PAR_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(PAR_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(PAR_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(PAR_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(PAR_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(PAR_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(PAR_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(PAR_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(PAR_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(PAR_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(PAR_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(PAR_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(PAR_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(PAR_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(PAR_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(PAR_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(PAR_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(PAR_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(PAR_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(PAR_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(PAR_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(PAR_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(PAR_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(PAR_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(PAR_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(PAR_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(PAR_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(PAR_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(PAR_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(PAR_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(PAR_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(PAR_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(PAR_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(PAR_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(PAR_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(PAR_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(PAR_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(PAR_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(PAR_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(PAR_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(PAR_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(PAR_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(PAR_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(PAR_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(PAR_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(PAR_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(PAR_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(PAR_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(PAR_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(PAR_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(PAR_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(PAR_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(PAR_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(PAR_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(PAR_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(PAR_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(PAR_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(PAR_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(PAR_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(PAR_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(PAR_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(PAR_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(PAR_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(PAR_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(PAR_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(PAR_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(PAR_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(PAR_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(PAR_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(PAR_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(PAR_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(PAR_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(PAR_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(PAR_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(PAR_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(PAR_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(PAR_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(PAR_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(PAR_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(PAR_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(PAR_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(PAR_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(PAR_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(PAR_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(PAR_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(PAR_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(PAR_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(PAR_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(PAR_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(PAR_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(PAR_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(PAR_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(PAR_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(PAR_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(PAR_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(PAR_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(PAR_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(PAR_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(PAR_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(PAR_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(PAR_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(PAR_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(PAR_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(PAR_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(PAR_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(PAR_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(PAR_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(PAR_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(PAR_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(PAR_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(PAR_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(PAR_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(PAR_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(PAR_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(PAR_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(PAR_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(PAR_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(PAR_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(PAR_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(PAR_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(PAR_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(PAR_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(PAR_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(PAR_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(PAR_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(PAR_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(PAR_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(PAR_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(PAR_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(PAR_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(PAR_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(PAR_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(PAR_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(PAR_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(PAR_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(PAR_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(PAR_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(PAR_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(PAR_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(PAR_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(PAR_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(PAR_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(PAR_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(PAR_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(PAR_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(PAR_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(PAR_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(PAR_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(PAR_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(PAR_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(PAR_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(PAR_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(PAR_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(PAR_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(PAR_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(PAR_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(PAR_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(PAR_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(PAR_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(PAR_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(PAR_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(PAR_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(PAR_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(PAR_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(PAR_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(PAR_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(PAR_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(PAR_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(PAR_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(PAR_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(PAR_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(PAR_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(PAR_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(PAR_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(PAR_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(PAR_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(PAR_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(PAR_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(PAR_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(PAR_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(PAR_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(PAR_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(PAR_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(PAR_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(PAR_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(PAR_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(PAR_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(PAR_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(PAR_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(PAR_io_pipe_phv_in_data_191),
    .io_pipe_phv_out_data_0(PAR_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(PAR_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(PAR_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(PAR_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(PAR_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(PAR_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(PAR_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(PAR_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(PAR_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(PAR_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(PAR_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(PAR_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(PAR_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(PAR_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(PAR_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(PAR_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(PAR_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(PAR_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(PAR_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(PAR_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(PAR_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(PAR_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(PAR_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(PAR_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(PAR_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(PAR_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(PAR_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(PAR_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(PAR_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(PAR_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(PAR_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(PAR_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(PAR_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(PAR_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(PAR_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(PAR_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(PAR_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(PAR_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(PAR_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(PAR_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(PAR_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(PAR_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(PAR_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(PAR_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(PAR_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(PAR_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(PAR_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(PAR_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(PAR_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(PAR_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(PAR_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(PAR_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(PAR_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(PAR_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(PAR_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(PAR_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(PAR_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(PAR_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(PAR_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(PAR_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(PAR_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(PAR_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(PAR_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(PAR_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(PAR_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(PAR_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(PAR_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(PAR_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(PAR_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(PAR_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(PAR_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(PAR_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(PAR_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(PAR_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(PAR_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(PAR_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(PAR_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(PAR_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(PAR_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(PAR_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(PAR_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(PAR_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(PAR_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(PAR_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(PAR_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(PAR_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(PAR_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(PAR_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(PAR_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(PAR_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(PAR_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(PAR_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(PAR_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(PAR_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(PAR_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(PAR_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(PAR_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(PAR_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(PAR_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(PAR_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(PAR_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(PAR_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(PAR_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(PAR_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(PAR_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(PAR_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(PAR_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(PAR_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(PAR_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(PAR_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(PAR_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(PAR_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(PAR_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(PAR_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(PAR_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(PAR_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(PAR_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(PAR_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(PAR_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(PAR_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(PAR_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(PAR_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(PAR_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(PAR_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(PAR_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(PAR_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(PAR_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(PAR_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(PAR_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(PAR_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(PAR_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(PAR_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(PAR_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(PAR_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(PAR_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(PAR_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(PAR_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(PAR_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(PAR_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(PAR_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(PAR_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(PAR_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(PAR_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(PAR_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(PAR_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(PAR_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(PAR_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(PAR_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(PAR_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(PAR_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(PAR_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(PAR_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(PAR_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(PAR_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(PAR_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(PAR_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(PAR_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(PAR_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(PAR_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(PAR_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(PAR_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(PAR_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(PAR_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(PAR_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(PAR_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(PAR_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(PAR_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(PAR_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(PAR_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(PAR_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(PAR_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(PAR_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(PAR_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(PAR_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(PAR_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(PAR_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(PAR_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(PAR_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(PAR_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(PAR_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(PAR_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(PAR_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(PAR_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(PAR_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(PAR_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(PAR_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(PAR_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(PAR_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(PAR_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(PAR_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(PAR_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(PAR_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(PAR_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(PAR_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(PAR_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(PAR_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(PAR_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(PAR_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(PAR_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(PAR_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(PAR_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(PAR_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(PAR_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(PAR_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(PAR_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(PAR_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(PAR_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(PAR_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(PAR_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(PAR_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(PAR_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(PAR_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(PAR_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(PAR_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(PAR_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(PAR_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(PAR_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(PAR_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(PAR_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(PAR_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(PAR_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(PAR_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(PAR_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(PAR_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(PAR_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(PAR_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(PAR_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(PAR_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(PAR_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(PAR_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(PAR_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(PAR_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(PAR_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(PAR_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(PAR_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(PAR_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(PAR_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(PAR_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(PAR_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(PAR_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(PAR_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(PAR_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(PAR_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(PAR_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(PAR_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(PAR_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(PAR_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(PAR_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(PAR_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(PAR_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(PAR_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(PAR_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(PAR_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(PAR_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(PAR_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(PAR_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_next_processor_id(PAR_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(PAR_io_pipe_phv_out_next_config_id),
    .io_mod_en(PAR_io_mod_en),
    .io_mod_last_mau_id_mod(PAR_io_mod_last_mau_id_mod),
    .io_mod_last_mau_id(PAR_io_mod_last_mau_id),
    .io_mod_cs(PAR_io_mod_cs),
    .io_mod_module_mod_state_id_mod(PAR_io_mod_module_mod_state_id_mod),
    .io_mod_module_mod_state_id(PAR_io_mod_module_mod_state_id),
    .io_mod_module_mod_sram_w_cs(PAR_io_mod_module_mod_sram_w_cs),
    .io_mod_module_mod_sram_w_en(PAR_io_mod_module_mod_sram_w_en),
    .io_mod_module_mod_sram_w_addr(PAR_io_mod_module_mod_sram_w_addr),
    .io_mod_module_mod_sram_w_data(PAR_io_mod_module_mod_sram_w_data)
  );
  ProcessorPISA proc_0 ( // @[pisa.scala 28:25]
    .clock(proc_0_clock),
    .io_pipe_phv_in_data_0(proc_0_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_0_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_0_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_0_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_0_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_0_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_0_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_0_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_0_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_0_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_0_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_0_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_0_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_0_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_0_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_0_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_0_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_0_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_0_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_0_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_0_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_0_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_0_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_0_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_0_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_0_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_0_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_0_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_0_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_0_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_0_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_0_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_0_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_0_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_0_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_0_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_0_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_0_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_0_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_0_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_0_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_0_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_0_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_0_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_0_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_0_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_0_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_0_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_0_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_0_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_0_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_0_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_0_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_0_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_0_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_0_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_0_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_0_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_0_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_0_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_0_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_0_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_0_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_0_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_0_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_0_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_0_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_0_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_0_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_0_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_0_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_0_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_0_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_0_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_0_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_0_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_0_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_0_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_0_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_0_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_0_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_0_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_0_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_0_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_0_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_0_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_0_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_0_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_0_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_0_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_0_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_0_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_0_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_0_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_0_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_0_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_0_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_0_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_0_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_0_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_0_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_0_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_0_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_0_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_0_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_0_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_0_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_0_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_0_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_0_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_0_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_0_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_0_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_0_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_0_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_0_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_0_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_0_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_0_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_0_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_0_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_0_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_0_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_0_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_0_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_0_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_0_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_0_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_0_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_0_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_0_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_0_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_0_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_0_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_0_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_0_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_0_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_0_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_0_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_0_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_0_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_0_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_0_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_0_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_0_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_0_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_0_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_0_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_0_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_0_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_0_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_0_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_0_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_0_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_0_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_0_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_0_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_0_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_0_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_0_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(proc_0_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(proc_0_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(proc_0_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(proc_0_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(proc_0_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(proc_0_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(proc_0_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(proc_0_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(proc_0_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(proc_0_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(proc_0_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(proc_0_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(proc_0_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(proc_0_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(proc_0_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(proc_0_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(proc_0_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(proc_0_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(proc_0_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(proc_0_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(proc_0_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(proc_0_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(proc_0_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(proc_0_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(proc_0_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(proc_0_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(proc_0_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(proc_0_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(proc_0_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(proc_0_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(proc_0_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(proc_0_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(proc_0_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(proc_0_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(proc_0_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(proc_0_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(proc_0_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(proc_0_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(proc_0_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(proc_0_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(proc_0_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(proc_0_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(proc_0_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(proc_0_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(proc_0_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(proc_0_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(proc_0_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(proc_0_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(proc_0_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(proc_0_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(proc_0_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(proc_0_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(proc_0_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(proc_0_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(proc_0_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(proc_0_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(proc_0_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(proc_0_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(proc_0_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(proc_0_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(proc_0_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(proc_0_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(proc_0_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(proc_0_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(proc_0_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(proc_0_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(proc_0_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(proc_0_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(proc_0_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(proc_0_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(proc_0_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(proc_0_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(proc_0_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(proc_0_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(proc_0_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(proc_0_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(proc_0_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(proc_0_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(proc_0_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(proc_0_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(proc_0_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(proc_0_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(proc_0_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(proc_0_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(proc_0_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(proc_0_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(proc_0_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(proc_0_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(proc_0_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(proc_0_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(proc_0_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(proc_0_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(proc_0_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(proc_0_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(proc_0_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(proc_0_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_next_processor_id(proc_0_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_0_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_0_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(proc_0_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_0_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_0_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_0_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_0_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_0_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_0_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_0_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_0_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_0_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_0_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_0_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_0_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_0_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_0_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_0_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_0_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_0_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_0_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_0_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_0_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_0_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_0_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_0_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_0_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_0_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_0_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_0_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_0_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_0_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_0_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_0_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_0_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_0_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_0_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_0_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_0_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_0_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_0_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_0_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_0_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_0_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_0_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_0_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_0_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_0_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_0_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_0_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_0_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_0_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_0_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_0_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_0_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_0_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_0_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_0_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_0_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_0_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_0_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_0_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_0_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_0_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_0_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_0_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_0_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_0_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_0_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_0_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_0_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_0_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_0_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_0_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_0_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_0_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_0_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_0_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_0_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_0_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_0_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_0_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_0_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_0_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_0_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_0_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_0_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_0_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_0_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_0_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_0_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_0_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_0_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_0_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_0_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_0_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_0_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_0_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_0_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_0_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_0_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_0_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_0_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_0_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_0_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_0_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_0_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_0_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_0_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_0_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_0_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_0_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_0_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_0_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_0_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_0_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_0_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_0_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_0_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_0_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_0_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_0_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_0_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_0_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_0_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_0_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_0_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_0_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_0_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_0_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_0_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_0_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_0_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_0_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_0_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_0_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_0_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_0_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_0_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_0_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_0_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_0_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_0_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_0_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_0_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_0_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_0_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_0_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_0_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_0_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_0_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_0_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_0_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_0_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_0_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_0_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_0_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_0_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_0_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_0_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_0_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_0_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(proc_0_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(proc_0_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(proc_0_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(proc_0_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(proc_0_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(proc_0_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(proc_0_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(proc_0_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(proc_0_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(proc_0_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(proc_0_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(proc_0_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(proc_0_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(proc_0_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(proc_0_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(proc_0_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(proc_0_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(proc_0_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(proc_0_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(proc_0_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(proc_0_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(proc_0_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(proc_0_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(proc_0_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(proc_0_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(proc_0_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(proc_0_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(proc_0_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(proc_0_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(proc_0_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(proc_0_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(proc_0_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(proc_0_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(proc_0_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(proc_0_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(proc_0_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(proc_0_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(proc_0_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(proc_0_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(proc_0_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(proc_0_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(proc_0_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(proc_0_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(proc_0_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(proc_0_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(proc_0_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(proc_0_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(proc_0_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(proc_0_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(proc_0_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(proc_0_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(proc_0_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(proc_0_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(proc_0_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(proc_0_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(proc_0_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(proc_0_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(proc_0_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(proc_0_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(proc_0_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(proc_0_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(proc_0_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(proc_0_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(proc_0_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(proc_0_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(proc_0_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(proc_0_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(proc_0_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(proc_0_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(proc_0_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(proc_0_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(proc_0_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(proc_0_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(proc_0_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(proc_0_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(proc_0_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(proc_0_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(proc_0_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(proc_0_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(proc_0_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(proc_0_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(proc_0_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(proc_0_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(proc_0_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(proc_0_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(proc_0_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(proc_0_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(proc_0_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(proc_0_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(proc_0_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(proc_0_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(proc_0_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(proc_0_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(proc_0_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(proc_0_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(proc_0_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_next_processor_id(proc_0_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_0_io_pipe_phv_out_next_config_id),
    .io_mod_mat_mod_en(proc_0_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_0_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_0_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_0_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_0_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_0_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_0_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_0_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_0_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_0_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_0_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_0_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_0_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_0_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_0_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_0_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_0_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_0_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_0_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_0_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_0_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_0_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_0_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_0_io_mod_exe_mod_data_1)
  );
  ProcessorPISA proc_1 ( // @[pisa.scala 28:25]
    .clock(proc_1_clock),
    .io_pipe_phv_in_data_0(proc_1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_1_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_1_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_1_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_1_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_1_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_1_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_1_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_1_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_1_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_1_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_1_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_1_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_1_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_1_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_1_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_1_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_1_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_1_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_1_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_1_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_1_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_1_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_1_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_1_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_1_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_1_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_1_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_1_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_1_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_1_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_1_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_1_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_1_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_1_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_1_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_1_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_1_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_1_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_1_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_1_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_1_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_1_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_1_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_1_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_1_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_1_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_1_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_1_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_1_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_1_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_1_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_1_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_1_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_1_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_1_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_1_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_1_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_1_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_1_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_1_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_1_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_1_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_1_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_1_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(proc_1_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(proc_1_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(proc_1_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(proc_1_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(proc_1_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(proc_1_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(proc_1_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(proc_1_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(proc_1_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(proc_1_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(proc_1_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(proc_1_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(proc_1_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(proc_1_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(proc_1_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(proc_1_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(proc_1_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(proc_1_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(proc_1_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(proc_1_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(proc_1_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(proc_1_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(proc_1_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(proc_1_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(proc_1_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(proc_1_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(proc_1_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(proc_1_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(proc_1_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(proc_1_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(proc_1_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(proc_1_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(proc_1_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(proc_1_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(proc_1_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(proc_1_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(proc_1_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(proc_1_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(proc_1_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(proc_1_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(proc_1_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(proc_1_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(proc_1_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(proc_1_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(proc_1_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(proc_1_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(proc_1_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(proc_1_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(proc_1_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(proc_1_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(proc_1_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(proc_1_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(proc_1_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(proc_1_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(proc_1_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(proc_1_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(proc_1_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(proc_1_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(proc_1_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(proc_1_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(proc_1_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(proc_1_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(proc_1_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(proc_1_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(proc_1_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(proc_1_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(proc_1_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(proc_1_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(proc_1_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(proc_1_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(proc_1_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(proc_1_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(proc_1_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(proc_1_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(proc_1_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(proc_1_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(proc_1_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(proc_1_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(proc_1_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(proc_1_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(proc_1_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(proc_1_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(proc_1_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(proc_1_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(proc_1_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(proc_1_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(proc_1_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(proc_1_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(proc_1_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(proc_1_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(proc_1_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(proc_1_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(proc_1_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(proc_1_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(proc_1_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(proc_1_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_next_processor_id(proc_1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_1_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(proc_1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_1_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_1_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_1_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_1_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_1_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_1_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_1_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_1_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_1_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_1_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_1_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_1_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_1_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_1_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_1_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_1_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_1_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_1_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_1_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_1_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_1_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_1_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_1_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_1_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_1_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_1_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_1_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_1_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_1_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_1_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_1_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_1_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_1_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_1_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_1_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_1_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_1_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_1_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_1_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_1_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_1_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_1_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_1_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_1_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_1_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_1_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_1_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_1_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_1_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_1_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_1_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_1_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_1_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_1_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_1_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_1_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_1_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_1_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_1_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_1_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_1_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_1_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_1_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_1_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(proc_1_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(proc_1_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(proc_1_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(proc_1_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(proc_1_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(proc_1_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(proc_1_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(proc_1_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(proc_1_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(proc_1_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(proc_1_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(proc_1_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(proc_1_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(proc_1_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(proc_1_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(proc_1_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(proc_1_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(proc_1_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(proc_1_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(proc_1_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(proc_1_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(proc_1_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(proc_1_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(proc_1_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(proc_1_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(proc_1_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(proc_1_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(proc_1_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(proc_1_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(proc_1_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(proc_1_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(proc_1_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(proc_1_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(proc_1_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(proc_1_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(proc_1_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(proc_1_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(proc_1_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(proc_1_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(proc_1_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(proc_1_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(proc_1_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(proc_1_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(proc_1_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(proc_1_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(proc_1_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(proc_1_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(proc_1_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(proc_1_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(proc_1_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(proc_1_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(proc_1_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(proc_1_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(proc_1_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(proc_1_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(proc_1_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(proc_1_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(proc_1_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(proc_1_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(proc_1_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(proc_1_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(proc_1_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(proc_1_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(proc_1_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(proc_1_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(proc_1_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(proc_1_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(proc_1_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(proc_1_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(proc_1_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(proc_1_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(proc_1_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(proc_1_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(proc_1_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(proc_1_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(proc_1_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(proc_1_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(proc_1_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(proc_1_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(proc_1_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(proc_1_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(proc_1_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(proc_1_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(proc_1_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(proc_1_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(proc_1_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(proc_1_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(proc_1_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(proc_1_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(proc_1_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(proc_1_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(proc_1_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(proc_1_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(proc_1_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(proc_1_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(proc_1_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_next_processor_id(proc_1_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_1_io_pipe_phv_out_next_config_id),
    .io_mod_mat_mod_en(proc_1_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_1_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_1_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_1_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_1_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_1_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_1_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_1_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_1_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_1_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_1_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_1_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_1_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_1_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_1_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_1_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_1_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_1_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_1_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_1_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_1_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_1_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_1_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_1_io_mod_exe_mod_data_1)
  );
  ProcessorPISA proc_2 ( // @[pisa.scala 28:25]
    .clock(proc_2_clock),
    .io_pipe_phv_in_data_0(proc_2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_2_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_2_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_2_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_2_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_2_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_2_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_2_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_2_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_2_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_2_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_2_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_2_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_2_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_2_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_2_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_2_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_2_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_2_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_2_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_2_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_2_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_2_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_2_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_2_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_2_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_2_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_2_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_2_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_2_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_2_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_2_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_2_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_2_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_2_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_2_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_2_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_2_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_2_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_2_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_2_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_2_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_2_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_2_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_2_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_2_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_2_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_2_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_2_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_2_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_2_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_2_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_2_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_2_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_2_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_2_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_2_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_2_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_2_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_2_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_2_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_2_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_2_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_2_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_2_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(proc_2_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(proc_2_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(proc_2_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(proc_2_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(proc_2_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(proc_2_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(proc_2_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(proc_2_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(proc_2_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(proc_2_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(proc_2_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(proc_2_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(proc_2_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(proc_2_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(proc_2_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(proc_2_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(proc_2_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(proc_2_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(proc_2_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(proc_2_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(proc_2_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(proc_2_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(proc_2_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(proc_2_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(proc_2_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(proc_2_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(proc_2_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(proc_2_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(proc_2_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(proc_2_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(proc_2_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(proc_2_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(proc_2_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(proc_2_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(proc_2_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(proc_2_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(proc_2_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(proc_2_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(proc_2_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(proc_2_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(proc_2_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(proc_2_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(proc_2_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(proc_2_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(proc_2_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(proc_2_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(proc_2_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(proc_2_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(proc_2_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(proc_2_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(proc_2_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(proc_2_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(proc_2_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(proc_2_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(proc_2_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(proc_2_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(proc_2_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(proc_2_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(proc_2_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(proc_2_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(proc_2_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(proc_2_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(proc_2_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(proc_2_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(proc_2_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(proc_2_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(proc_2_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(proc_2_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(proc_2_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(proc_2_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(proc_2_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(proc_2_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(proc_2_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(proc_2_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(proc_2_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(proc_2_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(proc_2_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(proc_2_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(proc_2_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(proc_2_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(proc_2_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(proc_2_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(proc_2_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(proc_2_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(proc_2_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(proc_2_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(proc_2_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(proc_2_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(proc_2_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(proc_2_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(proc_2_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(proc_2_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(proc_2_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(proc_2_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(proc_2_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(proc_2_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_next_processor_id(proc_2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_2_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(proc_2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_2_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_2_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_2_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_2_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_2_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_2_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_2_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_2_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_2_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_2_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_2_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_2_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_2_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_2_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_2_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_2_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_2_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_2_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_2_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_2_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_2_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_2_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_2_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_2_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_2_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_2_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_2_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_2_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_2_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_2_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_2_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_2_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_2_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_2_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_2_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_2_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_2_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_2_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_2_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_2_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_2_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_2_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_2_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_2_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_2_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_2_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_2_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_2_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_2_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_2_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_2_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_2_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_2_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_2_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_2_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_2_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_2_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_2_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_2_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_2_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_2_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_2_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_2_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_2_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(proc_2_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(proc_2_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(proc_2_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(proc_2_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(proc_2_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(proc_2_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(proc_2_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(proc_2_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(proc_2_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(proc_2_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(proc_2_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(proc_2_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(proc_2_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(proc_2_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(proc_2_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(proc_2_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(proc_2_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(proc_2_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(proc_2_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(proc_2_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(proc_2_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(proc_2_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(proc_2_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(proc_2_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(proc_2_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(proc_2_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(proc_2_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(proc_2_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(proc_2_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(proc_2_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(proc_2_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(proc_2_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(proc_2_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(proc_2_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(proc_2_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(proc_2_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(proc_2_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(proc_2_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(proc_2_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(proc_2_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(proc_2_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(proc_2_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(proc_2_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(proc_2_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(proc_2_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(proc_2_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(proc_2_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(proc_2_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(proc_2_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(proc_2_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(proc_2_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(proc_2_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(proc_2_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(proc_2_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(proc_2_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(proc_2_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(proc_2_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(proc_2_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(proc_2_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(proc_2_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(proc_2_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(proc_2_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(proc_2_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(proc_2_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(proc_2_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(proc_2_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(proc_2_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(proc_2_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(proc_2_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(proc_2_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(proc_2_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(proc_2_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(proc_2_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(proc_2_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(proc_2_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(proc_2_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(proc_2_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(proc_2_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(proc_2_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(proc_2_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(proc_2_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(proc_2_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(proc_2_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(proc_2_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(proc_2_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(proc_2_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(proc_2_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(proc_2_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(proc_2_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(proc_2_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(proc_2_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(proc_2_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(proc_2_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(proc_2_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(proc_2_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(proc_2_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_next_processor_id(proc_2_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_2_io_pipe_phv_out_next_config_id),
    .io_mod_mat_mod_en(proc_2_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_2_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_2_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_2_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_2_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_2_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_2_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_2_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_2_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_2_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_2_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_2_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_2_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_2_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_2_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_2_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_2_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_2_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_2_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_2_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_2_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_2_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_2_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_2_io_mod_exe_mod_data_1)
  );
  ProcessorPISA proc_3 ( // @[pisa.scala 28:25]
    .clock(proc_3_clock),
    .io_pipe_phv_in_data_0(proc_3_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_3_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_3_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_3_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_3_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_3_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_3_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_3_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_3_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_3_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_3_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_3_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_3_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_3_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_3_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_3_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_3_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_3_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_3_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_3_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_3_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_3_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_3_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_3_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_3_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_3_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_3_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_3_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_3_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_3_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_3_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_3_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_3_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_3_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_3_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_3_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_3_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_3_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_3_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_3_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_3_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_3_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_3_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_3_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_3_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_3_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_3_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_3_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_3_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_3_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_3_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_3_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_3_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_3_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_3_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_3_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_3_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_3_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_3_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_3_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_3_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_3_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_3_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_3_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_3_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_3_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_3_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_3_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_3_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_3_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_3_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_3_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_3_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_3_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_3_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_3_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_3_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_3_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_3_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_3_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_3_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_3_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_3_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_3_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_3_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_3_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_3_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_3_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_3_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_3_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_3_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_3_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_3_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_3_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_3_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_3_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_3_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_3_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_3_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_3_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_3_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_3_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_3_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_3_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_3_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_3_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_3_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_3_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_3_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_3_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_3_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_3_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_3_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_3_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_3_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_3_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_3_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_3_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_3_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_3_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_3_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_3_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_3_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_3_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_3_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_3_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_3_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_3_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_3_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_3_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_3_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_3_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_3_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_3_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_3_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_3_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_3_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_3_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_3_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_3_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_3_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_3_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_3_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_3_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_3_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_3_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_3_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_3_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_3_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_3_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_3_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_3_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_3_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_3_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_3_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_3_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_3_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_3_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_3_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_3_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(proc_3_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(proc_3_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(proc_3_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(proc_3_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(proc_3_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(proc_3_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(proc_3_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(proc_3_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(proc_3_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(proc_3_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(proc_3_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(proc_3_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(proc_3_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(proc_3_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(proc_3_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(proc_3_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(proc_3_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(proc_3_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(proc_3_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(proc_3_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(proc_3_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(proc_3_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(proc_3_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(proc_3_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(proc_3_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(proc_3_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(proc_3_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(proc_3_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(proc_3_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(proc_3_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(proc_3_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(proc_3_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(proc_3_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(proc_3_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(proc_3_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(proc_3_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(proc_3_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(proc_3_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(proc_3_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(proc_3_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(proc_3_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(proc_3_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(proc_3_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(proc_3_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(proc_3_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(proc_3_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(proc_3_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(proc_3_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(proc_3_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(proc_3_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(proc_3_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(proc_3_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(proc_3_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(proc_3_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(proc_3_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(proc_3_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(proc_3_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(proc_3_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(proc_3_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(proc_3_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(proc_3_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(proc_3_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(proc_3_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(proc_3_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(proc_3_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(proc_3_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(proc_3_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(proc_3_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(proc_3_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(proc_3_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(proc_3_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(proc_3_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(proc_3_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(proc_3_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(proc_3_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(proc_3_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(proc_3_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(proc_3_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(proc_3_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(proc_3_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(proc_3_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(proc_3_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(proc_3_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(proc_3_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(proc_3_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(proc_3_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(proc_3_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(proc_3_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(proc_3_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(proc_3_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(proc_3_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(proc_3_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(proc_3_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(proc_3_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(proc_3_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(proc_3_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_next_processor_id(proc_3_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_3_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_3_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(proc_3_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_3_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_3_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_3_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_3_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_3_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_3_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_3_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_3_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_3_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_3_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_3_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_3_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_3_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_3_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_3_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_3_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_3_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_3_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_3_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_3_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_3_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_3_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_3_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_3_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_3_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_3_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_3_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_3_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_3_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_3_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_3_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_3_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_3_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_3_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_3_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_3_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_3_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_3_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_3_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_3_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_3_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_3_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_3_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_3_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_3_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_3_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_3_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_3_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_3_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_3_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_3_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_3_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_3_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_3_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_3_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_3_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_3_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_3_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_3_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_3_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_3_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_3_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_3_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_3_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_3_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_3_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_3_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_3_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_3_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_3_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_3_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_3_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_3_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_3_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_3_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_3_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_3_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_3_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_3_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_3_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_3_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_3_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_3_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_3_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_3_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_3_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_3_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_3_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_3_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_3_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_3_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_3_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_3_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_3_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_3_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_3_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_3_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_3_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_3_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_3_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_3_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_3_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_3_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_3_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_3_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_3_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_3_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_3_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_3_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_3_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_3_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_3_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_3_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_3_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_3_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_3_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_3_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_3_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_3_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_3_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_3_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_3_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_3_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_3_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_3_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_3_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_3_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_3_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_3_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_3_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_3_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_3_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_3_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_3_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_3_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_3_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_3_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_3_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_3_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_3_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_3_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_3_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_3_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_3_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_3_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_3_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_3_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_3_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_3_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_3_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_3_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_3_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_3_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_3_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_3_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_3_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_3_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_3_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_3_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(proc_3_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(proc_3_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(proc_3_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(proc_3_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(proc_3_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(proc_3_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(proc_3_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(proc_3_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(proc_3_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(proc_3_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(proc_3_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(proc_3_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(proc_3_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(proc_3_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(proc_3_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(proc_3_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(proc_3_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(proc_3_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(proc_3_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(proc_3_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(proc_3_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(proc_3_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(proc_3_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(proc_3_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(proc_3_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(proc_3_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(proc_3_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(proc_3_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(proc_3_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(proc_3_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(proc_3_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(proc_3_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(proc_3_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(proc_3_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(proc_3_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(proc_3_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(proc_3_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(proc_3_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(proc_3_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(proc_3_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(proc_3_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(proc_3_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(proc_3_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(proc_3_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(proc_3_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(proc_3_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(proc_3_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(proc_3_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(proc_3_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(proc_3_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(proc_3_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(proc_3_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(proc_3_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(proc_3_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(proc_3_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(proc_3_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(proc_3_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(proc_3_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(proc_3_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(proc_3_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(proc_3_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(proc_3_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(proc_3_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(proc_3_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(proc_3_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(proc_3_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(proc_3_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(proc_3_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(proc_3_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(proc_3_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(proc_3_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(proc_3_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(proc_3_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(proc_3_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(proc_3_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(proc_3_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(proc_3_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(proc_3_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(proc_3_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(proc_3_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(proc_3_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(proc_3_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(proc_3_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(proc_3_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(proc_3_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(proc_3_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(proc_3_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(proc_3_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(proc_3_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(proc_3_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(proc_3_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(proc_3_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(proc_3_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(proc_3_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(proc_3_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(proc_3_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_next_processor_id(proc_3_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_3_io_pipe_phv_out_next_config_id),
    .io_mod_mat_mod_en(proc_3_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_3_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_3_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_3_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_3_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_3_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_3_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_3_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_3_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_3_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_3_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_3_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_3_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_3_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_3_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_3_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_3_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_3_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_3_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_3_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_3_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_3_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_3_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_3_io_mod_exe_mod_data_1)
  );
  ProcessorPISA proc_4 ( // @[pisa.scala 28:25]
    .clock(proc_4_clock),
    .io_pipe_phv_in_data_0(proc_4_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_4_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_4_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_4_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_4_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_4_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_4_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_4_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_4_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_4_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_4_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_4_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_4_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_4_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_4_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_4_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_4_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_4_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_4_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_4_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_4_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_4_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_4_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_4_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_4_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_4_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_4_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_4_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_4_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_4_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_4_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_4_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_4_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_4_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_4_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_4_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_4_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_4_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_4_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_4_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_4_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_4_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_4_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_4_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_4_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_4_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_4_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_4_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_4_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_4_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_4_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_4_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_4_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_4_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_4_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_4_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_4_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_4_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_4_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_4_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_4_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_4_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_4_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_4_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_4_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_4_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_4_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_4_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_4_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_4_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_4_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_4_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_4_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_4_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_4_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_4_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_4_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_4_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_4_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_4_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_4_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_4_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_4_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_4_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_4_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_4_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_4_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_4_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_4_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_4_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_4_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_4_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_4_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_4_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_4_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_4_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_4_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_4_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_4_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_4_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_4_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_4_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_4_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_4_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_4_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_4_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_4_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_4_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_4_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_4_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_4_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_4_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_4_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_4_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_4_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_4_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_4_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_4_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_4_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_4_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_4_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_4_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_4_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_4_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_4_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_4_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_4_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_4_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_4_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_4_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_4_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_4_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_4_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_4_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_4_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_4_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_4_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_4_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_4_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_4_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_4_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_4_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_4_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_4_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_4_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_4_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_4_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_4_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_4_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_4_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_4_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_4_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_4_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_4_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_4_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_4_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_4_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_4_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_4_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_4_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(proc_4_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(proc_4_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(proc_4_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(proc_4_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(proc_4_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(proc_4_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(proc_4_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(proc_4_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(proc_4_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(proc_4_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(proc_4_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(proc_4_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(proc_4_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(proc_4_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(proc_4_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(proc_4_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(proc_4_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(proc_4_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(proc_4_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(proc_4_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(proc_4_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(proc_4_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(proc_4_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(proc_4_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(proc_4_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(proc_4_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(proc_4_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(proc_4_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(proc_4_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(proc_4_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(proc_4_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(proc_4_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(proc_4_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(proc_4_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(proc_4_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(proc_4_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(proc_4_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(proc_4_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(proc_4_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(proc_4_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(proc_4_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(proc_4_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(proc_4_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(proc_4_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(proc_4_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(proc_4_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(proc_4_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(proc_4_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(proc_4_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(proc_4_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(proc_4_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(proc_4_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(proc_4_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(proc_4_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(proc_4_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(proc_4_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(proc_4_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(proc_4_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(proc_4_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(proc_4_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(proc_4_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(proc_4_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(proc_4_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(proc_4_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(proc_4_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(proc_4_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(proc_4_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(proc_4_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(proc_4_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(proc_4_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(proc_4_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(proc_4_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(proc_4_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(proc_4_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(proc_4_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(proc_4_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(proc_4_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(proc_4_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(proc_4_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(proc_4_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(proc_4_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(proc_4_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(proc_4_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(proc_4_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(proc_4_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(proc_4_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(proc_4_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(proc_4_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(proc_4_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(proc_4_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(proc_4_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(proc_4_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(proc_4_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(proc_4_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(proc_4_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(proc_4_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_next_processor_id(proc_4_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_4_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_4_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(proc_4_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_4_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_4_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_4_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_4_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_4_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_4_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_4_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_4_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_4_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_4_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_4_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_4_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_4_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_4_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_4_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_4_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_4_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_4_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_4_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_4_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_4_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_4_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_4_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_4_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_4_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_4_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_4_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_4_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_4_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_4_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_4_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_4_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_4_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_4_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_4_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_4_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_4_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_4_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_4_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_4_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_4_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_4_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_4_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_4_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_4_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_4_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_4_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_4_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_4_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_4_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_4_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_4_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_4_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_4_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_4_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_4_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_4_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_4_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_4_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_4_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_4_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_4_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_4_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_4_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_4_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_4_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_4_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_4_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_4_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_4_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_4_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_4_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_4_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_4_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_4_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_4_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_4_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_4_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_4_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_4_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_4_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_4_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_4_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_4_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_4_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_4_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_4_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_4_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_4_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_4_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_4_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_4_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_4_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_4_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_4_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_4_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_4_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_4_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_4_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_4_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_4_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_4_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_4_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_4_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_4_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_4_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_4_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_4_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_4_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_4_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_4_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_4_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_4_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_4_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_4_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_4_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_4_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_4_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_4_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_4_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_4_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_4_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_4_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_4_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_4_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_4_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_4_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_4_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_4_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_4_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_4_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_4_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_4_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_4_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_4_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_4_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_4_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_4_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_4_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_4_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_4_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_4_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_4_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_4_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_4_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_4_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_4_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_4_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_4_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_4_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_4_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_4_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_4_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_4_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_4_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_4_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_4_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_4_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_4_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(proc_4_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(proc_4_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(proc_4_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(proc_4_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(proc_4_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(proc_4_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(proc_4_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(proc_4_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(proc_4_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(proc_4_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(proc_4_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(proc_4_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(proc_4_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(proc_4_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(proc_4_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(proc_4_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(proc_4_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(proc_4_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(proc_4_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(proc_4_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(proc_4_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(proc_4_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(proc_4_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(proc_4_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(proc_4_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(proc_4_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(proc_4_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(proc_4_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(proc_4_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(proc_4_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(proc_4_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(proc_4_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(proc_4_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(proc_4_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(proc_4_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(proc_4_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(proc_4_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(proc_4_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(proc_4_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(proc_4_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(proc_4_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(proc_4_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(proc_4_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(proc_4_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(proc_4_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(proc_4_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(proc_4_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(proc_4_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(proc_4_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(proc_4_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(proc_4_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(proc_4_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(proc_4_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(proc_4_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(proc_4_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(proc_4_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(proc_4_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(proc_4_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(proc_4_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(proc_4_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(proc_4_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(proc_4_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(proc_4_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(proc_4_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(proc_4_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(proc_4_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(proc_4_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(proc_4_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(proc_4_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(proc_4_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(proc_4_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(proc_4_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(proc_4_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(proc_4_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(proc_4_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(proc_4_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(proc_4_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(proc_4_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(proc_4_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(proc_4_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(proc_4_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(proc_4_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(proc_4_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(proc_4_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(proc_4_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(proc_4_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(proc_4_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(proc_4_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(proc_4_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(proc_4_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(proc_4_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(proc_4_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(proc_4_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(proc_4_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(proc_4_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(proc_4_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_next_processor_id(proc_4_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_4_io_pipe_phv_out_next_config_id),
    .io_mod_mat_mod_en(proc_4_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_4_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_4_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_4_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_4_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_4_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_4_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_4_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_4_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_4_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_4_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_4_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_4_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_4_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_4_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_4_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_4_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_4_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_4_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_4_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_4_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_4_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_4_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_4_io_mod_exe_mod_data_1)
  );
  ProcessorPISA proc_5 ( // @[pisa.scala 28:25]
    .clock(proc_5_clock),
    .io_pipe_phv_in_data_0(proc_5_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_5_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_5_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_5_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_5_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_5_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_5_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_5_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_5_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_5_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_5_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_5_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_5_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_5_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_5_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_5_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_5_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_5_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_5_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_5_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_5_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_5_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_5_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_5_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_5_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_5_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_5_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_5_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_5_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_5_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_5_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_5_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_5_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_5_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_5_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_5_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_5_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_5_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_5_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_5_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_5_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_5_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_5_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_5_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_5_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_5_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_5_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_5_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_5_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_5_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_5_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_5_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_5_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_5_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_5_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_5_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_5_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_5_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_5_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_5_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_5_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_5_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_5_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_5_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_5_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_5_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_5_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_5_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_5_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_5_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_5_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_5_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_5_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_5_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_5_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_5_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_5_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_5_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_5_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_5_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_5_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_5_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_5_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_5_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_5_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_5_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_5_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_5_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_5_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_5_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_5_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_5_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_5_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_5_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_5_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_5_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_5_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_5_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_5_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_5_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_5_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_5_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_5_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_5_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_5_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_5_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_5_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_5_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_5_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_5_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_5_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_5_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_5_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_5_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_5_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_5_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_5_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_5_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_5_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_5_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_5_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_5_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_5_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_5_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_5_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_5_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_5_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_5_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_5_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_5_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_5_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_5_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_5_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_5_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_5_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_5_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_5_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_5_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_5_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_5_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_5_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_5_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_5_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_5_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_5_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_5_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_5_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_5_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_5_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_5_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_5_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_5_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_5_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_5_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_5_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_5_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_5_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_5_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_5_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_5_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(proc_5_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(proc_5_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(proc_5_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(proc_5_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(proc_5_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(proc_5_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(proc_5_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(proc_5_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(proc_5_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(proc_5_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(proc_5_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(proc_5_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(proc_5_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(proc_5_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(proc_5_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(proc_5_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(proc_5_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(proc_5_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(proc_5_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(proc_5_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(proc_5_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(proc_5_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(proc_5_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(proc_5_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(proc_5_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(proc_5_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(proc_5_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(proc_5_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(proc_5_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(proc_5_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(proc_5_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(proc_5_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(proc_5_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(proc_5_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(proc_5_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(proc_5_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(proc_5_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(proc_5_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(proc_5_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(proc_5_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(proc_5_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(proc_5_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(proc_5_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(proc_5_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(proc_5_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(proc_5_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(proc_5_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(proc_5_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(proc_5_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(proc_5_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(proc_5_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(proc_5_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(proc_5_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(proc_5_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(proc_5_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(proc_5_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(proc_5_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(proc_5_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(proc_5_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(proc_5_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(proc_5_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(proc_5_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(proc_5_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(proc_5_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(proc_5_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(proc_5_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(proc_5_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(proc_5_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(proc_5_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(proc_5_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(proc_5_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(proc_5_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(proc_5_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(proc_5_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(proc_5_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(proc_5_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(proc_5_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(proc_5_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(proc_5_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(proc_5_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(proc_5_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(proc_5_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(proc_5_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(proc_5_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(proc_5_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(proc_5_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(proc_5_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(proc_5_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(proc_5_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(proc_5_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(proc_5_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(proc_5_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(proc_5_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(proc_5_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(proc_5_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(proc_5_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_next_processor_id(proc_5_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_5_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_5_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(proc_5_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_5_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_5_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_5_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_5_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_5_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_5_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_5_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_5_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_5_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_5_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_5_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_5_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_5_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_5_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_5_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_5_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_5_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_5_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_5_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_5_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_5_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_5_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_5_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_5_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_5_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_5_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_5_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_5_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_5_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_5_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_5_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_5_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_5_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_5_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_5_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_5_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_5_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_5_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_5_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_5_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_5_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_5_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_5_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_5_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_5_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_5_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_5_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_5_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_5_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_5_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_5_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_5_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_5_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_5_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_5_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_5_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_5_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_5_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_5_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_5_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_5_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_5_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_5_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_5_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_5_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_5_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_5_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_5_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_5_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_5_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_5_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_5_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_5_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_5_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_5_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_5_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_5_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_5_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_5_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_5_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_5_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_5_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_5_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_5_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_5_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_5_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_5_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_5_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_5_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_5_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_5_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_5_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_5_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_5_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_5_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_5_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_5_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_5_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_5_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_5_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_5_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_5_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_5_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_5_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_5_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_5_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_5_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_5_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_5_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_5_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_5_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_5_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_5_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_5_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_5_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_5_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_5_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_5_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_5_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_5_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_5_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_5_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_5_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_5_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_5_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_5_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_5_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_5_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_5_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_5_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_5_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_5_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_5_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_5_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_5_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_5_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_5_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_5_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_5_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_5_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_5_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_5_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_5_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_5_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_5_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_5_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_5_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_5_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_5_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_5_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_5_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_5_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_5_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_5_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_5_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_5_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_5_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_5_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_5_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(proc_5_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(proc_5_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(proc_5_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(proc_5_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(proc_5_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(proc_5_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(proc_5_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(proc_5_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(proc_5_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(proc_5_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(proc_5_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(proc_5_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(proc_5_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(proc_5_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(proc_5_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(proc_5_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(proc_5_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(proc_5_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(proc_5_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(proc_5_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(proc_5_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(proc_5_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(proc_5_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(proc_5_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(proc_5_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(proc_5_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(proc_5_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(proc_5_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(proc_5_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(proc_5_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(proc_5_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(proc_5_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(proc_5_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(proc_5_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(proc_5_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(proc_5_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(proc_5_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(proc_5_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(proc_5_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(proc_5_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(proc_5_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(proc_5_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(proc_5_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(proc_5_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(proc_5_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(proc_5_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(proc_5_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(proc_5_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(proc_5_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(proc_5_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(proc_5_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(proc_5_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(proc_5_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(proc_5_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(proc_5_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(proc_5_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(proc_5_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(proc_5_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(proc_5_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(proc_5_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(proc_5_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(proc_5_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(proc_5_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(proc_5_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(proc_5_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(proc_5_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(proc_5_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(proc_5_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(proc_5_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(proc_5_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(proc_5_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(proc_5_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(proc_5_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(proc_5_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(proc_5_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(proc_5_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(proc_5_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(proc_5_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(proc_5_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(proc_5_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(proc_5_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(proc_5_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(proc_5_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(proc_5_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(proc_5_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(proc_5_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(proc_5_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(proc_5_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(proc_5_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(proc_5_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(proc_5_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(proc_5_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(proc_5_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(proc_5_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(proc_5_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(proc_5_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_next_processor_id(proc_5_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_5_io_pipe_phv_out_next_config_id),
    .io_mod_mat_mod_en(proc_5_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_5_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_5_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_5_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_5_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_5_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_5_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_5_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_5_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_5_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_5_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_5_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_5_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_5_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_5_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_5_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_5_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_5_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_5_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_5_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_5_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_5_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_5_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_5_io_mod_exe_mod_data_1)
  );
  ProcessorPISA proc_6 ( // @[pisa.scala 28:25]
    .clock(proc_6_clock),
    .io_pipe_phv_in_data_0(proc_6_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_6_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_6_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_6_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_6_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_6_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_6_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_6_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_6_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_6_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_6_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_6_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_6_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_6_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_6_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_6_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_6_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_6_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_6_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_6_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_6_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_6_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_6_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_6_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_6_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_6_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_6_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_6_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_6_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_6_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_6_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_6_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_6_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_6_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_6_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_6_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_6_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_6_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_6_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_6_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_6_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_6_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_6_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_6_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_6_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_6_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_6_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_6_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_6_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_6_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_6_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_6_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_6_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_6_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_6_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_6_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_6_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_6_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_6_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_6_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_6_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_6_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_6_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_6_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_6_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_6_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_6_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_6_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_6_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_6_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_6_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_6_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_6_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_6_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_6_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_6_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_6_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_6_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_6_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_6_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_6_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_6_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_6_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_6_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_6_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_6_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_6_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_6_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_6_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_6_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_6_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_6_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_6_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_6_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_6_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_6_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_6_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_6_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_6_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_6_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_6_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_6_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_6_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_6_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_6_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_6_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_6_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_6_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_6_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_6_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_6_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_6_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_6_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_6_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_6_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_6_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_6_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_6_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_6_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_6_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_6_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_6_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_6_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_6_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_6_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_6_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_6_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_6_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_6_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_6_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_6_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_6_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_6_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_6_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_6_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_6_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_6_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_6_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_6_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_6_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_6_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_6_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_6_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_6_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_6_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_6_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_6_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_6_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_6_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_6_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_6_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_6_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_6_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_6_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_6_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_6_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_6_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_6_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_6_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_6_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(proc_6_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(proc_6_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(proc_6_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(proc_6_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(proc_6_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(proc_6_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(proc_6_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(proc_6_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(proc_6_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(proc_6_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(proc_6_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(proc_6_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(proc_6_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(proc_6_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(proc_6_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(proc_6_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(proc_6_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(proc_6_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(proc_6_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(proc_6_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(proc_6_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(proc_6_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(proc_6_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(proc_6_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(proc_6_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(proc_6_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(proc_6_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(proc_6_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(proc_6_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(proc_6_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(proc_6_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(proc_6_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(proc_6_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(proc_6_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(proc_6_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(proc_6_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(proc_6_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(proc_6_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(proc_6_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(proc_6_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(proc_6_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(proc_6_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(proc_6_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(proc_6_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(proc_6_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(proc_6_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(proc_6_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(proc_6_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(proc_6_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(proc_6_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(proc_6_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(proc_6_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(proc_6_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(proc_6_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(proc_6_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(proc_6_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(proc_6_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(proc_6_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(proc_6_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(proc_6_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(proc_6_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(proc_6_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(proc_6_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(proc_6_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(proc_6_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(proc_6_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(proc_6_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(proc_6_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(proc_6_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(proc_6_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(proc_6_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(proc_6_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(proc_6_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(proc_6_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(proc_6_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(proc_6_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(proc_6_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(proc_6_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(proc_6_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(proc_6_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(proc_6_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(proc_6_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(proc_6_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(proc_6_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(proc_6_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(proc_6_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(proc_6_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(proc_6_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(proc_6_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(proc_6_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(proc_6_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(proc_6_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(proc_6_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(proc_6_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(proc_6_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(proc_6_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_next_processor_id(proc_6_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_6_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_6_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(proc_6_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_6_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_6_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_6_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_6_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_6_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_6_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_6_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_6_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_6_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_6_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_6_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_6_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_6_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_6_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_6_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_6_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_6_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_6_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_6_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_6_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_6_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_6_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_6_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_6_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_6_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_6_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_6_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_6_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_6_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_6_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_6_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_6_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_6_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_6_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_6_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_6_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_6_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_6_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_6_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_6_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_6_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_6_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_6_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_6_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_6_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_6_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_6_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_6_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_6_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_6_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_6_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_6_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_6_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_6_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_6_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_6_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_6_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_6_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_6_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_6_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_6_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_6_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_6_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_6_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_6_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_6_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_6_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_6_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_6_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_6_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_6_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_6_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_6_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_6_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_6_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_6_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_6_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_6_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_6_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_6_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_6_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_6_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_6_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_6_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_6_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_6_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_6_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_6_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_6_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_6_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_6_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_6_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_6_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_6_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_6_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_6_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_6_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_6_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_6_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_6_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_6_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_6_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_6_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_6_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_6_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_6_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_6_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_6_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_6_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_6_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_6_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_6_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_6_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_6_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_6_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_6_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_6_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_6_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_6_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_6_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_6_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_6_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_6_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_6_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_6_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_6_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_6_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_6_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_6_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_6_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_6_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_6_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_6_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_6_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_6_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_6_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_6_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_6_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_6_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_6_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_6_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_6_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_6_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_6_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_6_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_6_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_6_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_6_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_6_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_6_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_6_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_6_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_6_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_6_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_6_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_6_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_6_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_6_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_6_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(proc_6_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(proc_6_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(proc_6_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(proc_6_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(proc_6_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(proc_6_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(proc_6_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(proc_6_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(proc_6_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(proc_6_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(proc_6_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(proc_6_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(proc_6_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(proc_6_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(proc_6_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(proc_6_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(proc_6_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(proc_6_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(proc_6_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(proc_6_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(proc_6_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(proc_6_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(proc_6_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(proc_6_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(proc_6_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(proc_6_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(proc_6_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(proc_6_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(proc_6_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(proc_6_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(proc_6_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(proc_6_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(proc_6_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(proc_6_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(proc_6_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(proc_6_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(proc_6_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(proc_6_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(proc_6_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(proc_6_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(proc_6_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(proc_6_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(proc_6_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(proc_6_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(proc_6_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(proc_6_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(proc_6_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(proc_6_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(proc_6_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(proc_6_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(proc_6_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(proc_6_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(proc_6_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(proc_6_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(proc_6_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(proc_6_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(proc_6_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(proc_6_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(proc_6_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(proc_6_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(proc_6_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(proc_6_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(proc_6_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(proc_6_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(proc_6_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(proc_6_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(proc_6_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(proc_6_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(proc_6_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(proc_6_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(proc_6_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(proc_6_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(proc_6_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(proc_6_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(proc_6_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(proc_6_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(proc_6_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(proc_6_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(proc_6_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(proc_6_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(proc_6_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(proc_6_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(proc_6_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(proc_6_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(proc_6_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(proc_6_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(proc_6_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(proc_6_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(proc_6_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(proc_6_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(proc_6_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(proc_6_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(proc_6_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(proc_6_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(proc_6_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(proc_6_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_next_processor_id(proc_6_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_6_io_pipe_phv_out_next_config_id),
    .io_mod_mat_mod_en(proc_6_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_6_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_6_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_6_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_6_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_6_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_6_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_6_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_6_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_6_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_6_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_6_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_6_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_6_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_6_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_6_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_6_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_6_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_6_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_6_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_6_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_6_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_6_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_6_io_mod_exe_mod_data_1)
  );
  ProcessorPISA proc_7 ( // @[pisa.scala 28:25]
    .clock(proc_7_clock),
    .io_pipe_phv_in_data_0(proc_7_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_7_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_7_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_7_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_7_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_7_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_7_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_7_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_7_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_7_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_7_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_7_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_7_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_7_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_7_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_7_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_7_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_7_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_7_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_7_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_7_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_7_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_7_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_7_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_7_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_7_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_7_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_7_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_7_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_7_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_7_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_7_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_7_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_7_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_7_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_7_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_7_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_7_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_7_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_7_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_7_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_7_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_7_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_7_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_7_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_7_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_7_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_7_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_7_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_7_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_7_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_7_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_7_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_7_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_7_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_7_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_7_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_7_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_7_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_7_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_7_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_7_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_7_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_7_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_7_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_7_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_7_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_7_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_7_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_7_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_7_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_7_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_7_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_7_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_7_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_7_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_7_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_7_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_7_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_7_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_7_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_7_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_7_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_7_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_7_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_7_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_7_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_7_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_7_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_7_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_7_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_7_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_7_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_7_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_7_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_7_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_7_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_7_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_7_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_7_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_7_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_7_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_7_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_7_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_7_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_7_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_7_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_7_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_7_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_7_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_7_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_7_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_7_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_7_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_7_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_7_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_7_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_7_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_7_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_7_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_7_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_7_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_7_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_7_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_7_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_7_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_7_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_7_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_7_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_7_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_7_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_7_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_7_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_7_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_7_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_7_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_7_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_7_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_7_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_7_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_7_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_7_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_7_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_7_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_7_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_7_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_7_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_7_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_7_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_7_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_7_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_7_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_7_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_7_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_7_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_7_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_7_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_7_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_7_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_7_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(proc_7_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(proc_7_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(proc_7_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(proc_7_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(proc_7_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(proc_7_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(proc_7_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(proc_7_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(proc_7_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(proc_7_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(proc_7_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(proc_7_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(proc_7_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(proc_7_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(proc_7_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(proc_7_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(proc_7_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(proc_7_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(proc_7_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(proc_7_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(proc_7_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(proc_7_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(proc_7_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(proc_7_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(proc_7_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(proc_7_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(proc_7_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(proc_7_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(proc_7_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(proc_7_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(proc_7_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(proc_7_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(proc_7_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(proc_7_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(proc_7_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(proc_7_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(proc_7_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(proc_7_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(proc_7_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(proc_7_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(proc_7_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(proc_7_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(proc_7_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(proc_7_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(proc_7_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(proc_7_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(proc_7_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(proc_7_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(proc_7_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(proc_7_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(proc_7_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(proc_7_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(proc_7_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(proc_7_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(proc_7_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(proc_7_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(proc_7_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(proc_7_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(proc_7_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(proc_7_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(proc_7_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(proc_7_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(proc_7_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(proc_7_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(proc_7_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(proc_7_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(proc_7_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(proc_7_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(proc_7_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(proc_7_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(proc_7_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(proc_7_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(proc_7_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(proc_7_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(proc_7_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(proc_7_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(proc_7_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(proc_7_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(proc_7_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(proc_7_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(proc_7_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(proc_7_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(proc_7_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(proc_7_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(proc_7_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(proc_7_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(proc_7_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(proc_7_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(proc_7_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(proc_7_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(proc_7_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(proc_7_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(proc_7_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(proc_7_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(proc_7_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(proc_7_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_next_processor_id(proc_7_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_7_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_7_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(proc_7_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_7_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_7_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_7_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_7_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_7_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_7_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_7_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_7_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_7_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_7_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_7_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_7_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_7_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_7_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_7_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_7_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_7_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_7_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_7_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_7_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_7_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_7_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_7_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_7_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_7_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_7_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_7_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_7_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_7_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_7_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_7_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_7_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_7_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_7_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_7_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_7_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_7_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_7_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_7_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_7_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_7_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_7_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_7_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_7_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_7_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_7_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_7_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_7_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_7_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_7_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_7_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_7_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_7_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_7_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_7_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_7_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_7_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_7_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_7_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_7_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_7_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_7_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_7_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_7_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_7_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_7_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_7_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_7_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_7_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_7_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_7_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_7_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_7_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_7_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_7_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_7_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_7_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_7_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_7_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_7_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_7_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_7_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_7_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_7_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_7_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_7_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_7_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_7_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_7_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_7_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_7_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_7_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_7_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_7_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_7_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_7_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_7_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_7_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_7_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_7_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_7_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_7_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_7_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_7_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_7_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_7_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_7_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_7_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_7_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_7_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_7_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_7_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_7_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_7_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_7_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_7_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_7_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_7_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_7_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_7_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_7_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_7_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_7_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_7_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_7_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_7_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_7_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_7_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_7_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_7_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_7_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_7_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_7_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_7_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_7_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_7_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_7_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_7_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_7_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_7_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_7_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_7_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_7_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_7_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_7_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_7_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_7_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_7_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_7_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_7_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_7_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_7_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_7_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_7_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_7_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_7_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_7_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_7_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_7_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(proc_7_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(proc_7_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(proc_7_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(proc_7_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(proc_7_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(proc_7_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(proc_7_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(proc_7_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(proc_7_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(proc_7_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(proc_7_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(proc_7_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(proc_7_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(proc_7_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(proc_7_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(proc_7_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(proc_7_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(proc_7_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(proc_7_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(proc_7_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(proc_7_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(proc_7_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(proc_7_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(proc_7_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(proc_7_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(proc_7_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(proc_7_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(proc_7_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(proc_7_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(proc_7_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(proc_7_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(proc_7_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(proc_7_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(proc_7_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(proc_7_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(proc_7_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(proc_7_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(proc_7_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(proc_7_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(proc_7_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(proc_7_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(proc_7_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(proc_7_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(proc_7_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(proc_7_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(proc_7_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(proc_7_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(proc_7_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(proc_7_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(proc_7_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(proc_7_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(proc_7_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(proc_7_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(proc_7_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(proc_7_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(proc_7_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(proc_7_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(proc_7_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(proc_7_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(proc_7_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(proc_7_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(proc_7_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(proc_7_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(proc_7_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(proc_7_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(proc_7_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(proc_7_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(proc_7_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(proc_7_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(proc_7_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(proc_7_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(proc_7_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(proc_7_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(proc_7_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(proc_7_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(proc_7_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(proc_7_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(proc_7_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(proc_7_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(proc_7_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(proc_7_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(proc_7_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(proc_7_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(proc_7_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(proc_7_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(proc_7_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(proc_7_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(proc_7_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(proc_7_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(proc_7_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(proc_7_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(proc_7_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(proc_7_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(proc_7_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(proc_7_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(proc_7_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_next_processor_id(proc_7_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_7_io_pipe_phv_out_next_config_id),
    .io_mod_mat_mod_en(proc_7_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_7_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_7_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_7_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_7_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_7_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_7_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_7_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_7_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_7_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_7_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_7_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_7_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_7_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_7_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_7_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_7_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_7_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_7_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_7_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_7_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_7_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_7_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_7_io_mod_exe_mod_data_1)
  );
  ProcessorPISA proc_8 ( // @[pisa.scala 28:25]
    .clock(proc_8_clock),
    .io_pipe_phv_in_data_0(proc_8_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_8_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_8_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_8_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_8_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_8_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_8_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_8_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_8_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_8_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_8_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_8_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_8_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_8_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_8_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_8_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_8_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_8_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_8_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_8_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_8_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_8_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_8_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_8_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_8_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_8_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_8_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_8_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_8_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_8_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_8_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_8_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_8_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_8_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_8_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_8_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_8_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_8_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_8_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_8_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_8_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_8_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_8_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_8_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_8_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_8_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_8_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_8_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_8_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_8_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_8_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_8_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_8_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_8_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_8_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_8_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_8_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_8_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_8_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_8_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_8_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_8_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_8_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_8_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_8_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_8_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_8_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_8_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_8_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_8_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_8_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_8_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_8_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_8_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_8_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_8_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_8_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_8_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_8_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_8_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_8_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_8_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_8_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_8_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_8_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_8_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_8_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_8_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_8_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_8_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_8_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_8_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_8_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_8_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_8_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_8_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_8_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_8_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_8_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_8_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_8_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_8_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_8_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_8_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_8_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_8_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_8_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_8_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_8_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_8_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_8_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_8_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_8_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_8_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_8_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_8_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_8_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_8_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_8_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_8_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_8_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_8_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_8_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_8_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_8_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_8_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_8_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_8_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_8_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_8_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_8_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_8_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_8_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_8_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_8_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_8_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_8_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_8_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_8_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_8_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_8_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_8_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_8_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_8_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_8_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_8_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_8_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_8_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_8_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_8_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_8_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_8_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_8_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_8_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_8_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_8_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_8_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_8_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_8_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_8_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(proc_8_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(proc_8_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(proc_8_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(proc_8_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(proc_8_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(proc_8_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(proc_8_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(proc_8_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(proc_8_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(proc_8_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(proc_8_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(proc_8_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(proc_8_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(proc_8_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(proc_8_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(proc_8_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(proc_8_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(proc_8_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(proc_8_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(proc_8_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(proc_8_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(proc_8_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(proc_8_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(proc_8_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(proc_8_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(proc_8_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(proc_8_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(proc_8_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(proc_8_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(proc_8_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(proc_8_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(proc_8_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(proc_8_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(proc_8_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(proc_8_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(proc_8_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(proc_8_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(proc_8_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(proc_8_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(proc_8_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(proc_8_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(proc_8_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(proc_8_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(proc_8_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(proc_8_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(proc_8_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(proc_8_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(proc_8_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(proc_8_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(proc_8_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(proc_8_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(proc_8_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(proc_8_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(proc_8_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(proc_8_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(proc_8_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(proc_8_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(proc_8_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(proc_8_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(proc_8_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(proc_8_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(proc_8_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(proc_8_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(proc_8_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(proc_8_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(proc_8_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(proc_8_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(proc_8_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(proc_8_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(proc_8_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(proc_8_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(proc_8_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(proc_8_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(proc_8_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(proc_8_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(proc_8_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(proc_8_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(proc_8_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(proc_8_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(proc_8_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(proc_8_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(proc_8_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(proc_8_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(proc_8_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(proc_8_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(proc_8_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(proc_8_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(proc_8_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(proc_8_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(proc_8_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(proc_8_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(proc_8_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(proc_8_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(proc_8_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(proc_8_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(proc_8_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_next_processor_id(proc_8_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_8_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_8_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(proc_8_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_8_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_8_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_8_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_8_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_8_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_8_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_8_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_8_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_8_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_8_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_8_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_8_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_8_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_8_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_8_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_8_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_8_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_8_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_8_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_8_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_8_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_8_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_8_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_8_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_8_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_8_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_8_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_8_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_8_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_8_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_8_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_8_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_8_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_8_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_8_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_8_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_8_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_8_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_8_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_8_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_8_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_8_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_8_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_8_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_8_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_8_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_8_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_8_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_8_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_8_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_8_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_8_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_8_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_8_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_8_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_8_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_8_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_8_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_8_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_8_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_8_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_8_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_8_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_8_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_8_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_8_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_8_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_8_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_8_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_8_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_8_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_8_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_8_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_8_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_8_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_8_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_8_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_8_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_8_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_8_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_8_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_8_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_8_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_8_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_8_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_8_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_8_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_8_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_8_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_8_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_8_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_8_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_8_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_8_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_8_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_8_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_8_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_8_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_8_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_8_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_8_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_8_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_8_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_8_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_8_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_8_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_8_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_8_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_8_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_8_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_8_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_8_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_8_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_8_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_8_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_8_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_8_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_8_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_8_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_8_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_8_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_8_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_8_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_8_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_8_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_8_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_8_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_8_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_8_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_8_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_8_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_8_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_8_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_8_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_8_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_8_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_8_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_8_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_8_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_8_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_8_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_8_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_8_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_8_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_8_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_8_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_8_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_8_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_8_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_8_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_8_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_8_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_8_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_8_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_8_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_8_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_8_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_8_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_8_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(proc_8_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(proc_8_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(proc_8_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(proc_8_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(proc_8_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(proc_8_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(proc_8_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(proc_8_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(proc_8_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(proc_8_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(proc_8_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(proc_8_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(proc_8_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(proc_8_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(proc_8_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(proc_8_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(proc_8_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(proc_8_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(proc_8_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(proc_8_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(proc_8_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(proc_8_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(proc_8_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(proc_8_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(proc_8_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(proc_8_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(proc_8_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(proc_8_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(proc_8_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(proc_8_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(proc_8_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(proc_8_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(proc_8_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(proc_8_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(proc_8_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(proc_8_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(proc_8_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(proc_8_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(proc_8_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(proc_8_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(proc_8_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(proc_8_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(proc_8_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(proc_8_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(proc_8_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(proc_8_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(proc_8_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(proc_8_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(proc_8_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(proc_8_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(proc_8_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(proc_8_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(proc_8_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(proc_8_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(proc_8_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(proc_8_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(proc_8_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(proc_8_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(proc_8_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(proc_8_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(proc_8_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(proc_8_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(proc_8_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(proc_8_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(proc_8_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(proc_8_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(proc_8_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(proc_8_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(proc_8_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(proc_8_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(proc_8_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(proc_8_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(proc_8_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(proc_8_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(proc_8_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(proc_8_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(proc_8_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(proc_8_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(proc_8_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(proc_8_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(proc_8_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(proc_8_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(proc_8_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(proc_8_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(proc_8_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(proc_8_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(proc_8_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(proc_8_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(proc_8_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(proc_8_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(proc_8_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(proc_8_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(proc_8_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(proc_8_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(proc_8_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(proc_8_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_next_processor_id(proc_8_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_8_io_pipe_phv_out_next_config_id),
    .io_mod_mat_mod_en(proc_8_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_8_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_8_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_8_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_8_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_8_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_8_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_8_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_8_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_8_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_8_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_8_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_8_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_8_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_8_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_8_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_8_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_8_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_8_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_8_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_8_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_8_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_8_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_8_io_mod_exe_mod_data_1)
  );
  ProcessorPISA proc_9 ( // @[pisa.scala 28:25]
    .clock(proc_9_clock),
    .io_pipe_phv_in_data_0(proc_9_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_9_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_9_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_9_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_9_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_9_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_9_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_9_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_9_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_9_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_9_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_9_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_9_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_9_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_9_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_9_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_9_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_9_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_9_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_9_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_9_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_9_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_9_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_9_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_9_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_9_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_9_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_9_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_9_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_9_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_9_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_9_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_9_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_9_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_9_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_9_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_9_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_9_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_9_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_9_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_9_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_9_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_9_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_9_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_9_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_9_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_9_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_9_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_9_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_9_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_9_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_9_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_9_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_9_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_9_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_9_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_9_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_9_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_9_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_9_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_9_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_9_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_9_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_9_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_9_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_9_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_9_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_9_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_9_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_9_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_9_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_9_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_9_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_9_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_9_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_9_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_9_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_9_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_9_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_9_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_9_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_9_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_9_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_9_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_9_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_9_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_9_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_9_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_9_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_9_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_9_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_9_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_9_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_9_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_9_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_9_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_9_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_9_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_9_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_9_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_9_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_9_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_9_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_9_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_9_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_9_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_9_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_9_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_9_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_9_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_9_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_9_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_9_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_9_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_9_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_9_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_9_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_9_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_9_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_9_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_9_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_9_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_9_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_9_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_9_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_9_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_9_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_9_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_9_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_9_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_9_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_9_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_9_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_9_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_9_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_9_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_9_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_9_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_9_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_9_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_9_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_9_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_9_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_9_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_9_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_9_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_9_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_9_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_9_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_9_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_9_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_9_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_9_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_9_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_9_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_9_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_9_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_9_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_9_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_9_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(proc_9_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(proc_9_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(proc_9_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(proc_9_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(proc_9_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(proc_9_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(proc_9_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(proc_9_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(proc_9_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(proc_9_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(proc_9_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(proc_9_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(proc_9_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(proc_9_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(proc_9_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(proc_9_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(proc_9_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(proc_9_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(proc_9_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(proc_9_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(proc_9_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(proc_9_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(proc_9_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(proc_9_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(proc_9_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(proc_9_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(proc_9_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(proc_9_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(proc_9_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(proc_9_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(proc_9_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(proc_9_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(proc_9_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(proc_9_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(proc_9_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(proc_9_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(proc_9_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(proc_9_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(proc_9_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(proc_9_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(proc_9_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(proc_9_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(proc_9_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(proc_9_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(proc_9_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(proc_9_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(proc_9_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(proc_9_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(proc_9_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(proc_9_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(proc_9_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(proc_9_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(proc_9_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(proc_9_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(proc_9_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(proc_9_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(proc_9_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(proc_9_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(proc_9_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(proc_9_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(proc_9_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(proc_9_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(proc_9_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(proc_9_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(proc_9_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(proc_9_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(proc_9_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(proc_9_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(proc_9_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(proc_9_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(proc_9_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(proc_9_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(proc_9_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(proc_9_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(proc_9_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(proc_9_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(proc_9_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(proc_9_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(proc_9_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(proc_9_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(proc_9_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(proc_9_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(proc_9_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(proc_9_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(proc_9_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(proc_9_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(proc_9_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(proc_9_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(proc_9_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(proc_9_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(proc_9_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(proc_9_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(proc_9_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(proc_9_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(proc_9_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(proc_9_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_next_processor_id(proc_9_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_9_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_9_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(proc_9_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_9_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_9_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_9_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_9_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_9_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_9_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_9_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_9_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_9_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_9_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_9_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_9_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_9_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_9_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_9_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_9_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_9_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_9_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_9_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_9_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_9_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_9_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_9_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_9_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_9_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_9_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_9_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_9_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_9_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_9_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_9_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_9_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_9_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_9_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_9_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_9_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_9_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_9_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_9_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_9_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_9_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_9_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_9_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_9_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_9_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_9_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_9_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_9_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_9_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_9_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_9_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_9_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_9_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_9_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_9_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_9_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_9_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_9_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_9_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_9_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_9_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_9_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_9_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_9_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_9_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_9_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_9_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_9_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_9_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_9_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_9_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_9_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_9_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_9_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_9_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_9_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_9_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_9_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_9_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_9_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_9_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_9_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_9_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_9_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_9_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_9_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_9_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_9_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_9_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_9_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_9_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_9_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_9_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_9_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_9_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_9_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_9_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_9_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_9_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_9_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_9_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_9_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_9_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_9_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_9_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_9_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_9_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_9_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_9_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_9_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_9_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_9_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_9_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_9_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_9_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_9_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_9_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_9_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_9_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_9_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_9_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_9_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_9_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_9_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_9_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_9_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_9_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_9_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_9_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_9_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_9_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_9_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_9_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_9_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_9_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_9_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_9_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_9_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_9_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_9_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_9_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_9_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_9_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_9_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_9_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_9_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_9_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_9_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_9_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_9_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_9_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_9_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_9_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_9_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_9_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_9_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_9_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_9_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_9_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(proc_9_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(proc_9_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(proc_9_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(proc_9_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(proc_9_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(proc_9_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(proc_9_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(proc_9_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(proc_9_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(proc_9_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(proc_9_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(proc_9_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(proc_9_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(proc_9_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(proc_9_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(proc_9_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(proc_9_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(proc_9_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(proc_9_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(proc_9_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(proc_9_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(proc_9_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(proc_9_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(proc_9_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(proc_9_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(proc_9_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(proc_9_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(proc_9_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(proc_9_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(proc_9_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(proc_9_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(proc_9_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(proc_9_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(proc_9_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(proc_9_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(proc_9_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(proc_9_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(proc_9_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(proc_9_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(proc_9_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(proc_9_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(proc_9_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(proc_9_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(proc_9_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(proc_9_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(proc_9_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(proc_9_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(proc_9_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(proc_9_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(proc_9_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(proc_9_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(proc_9_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(proc_9_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(proc_9_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(proc_9_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(proc_9_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(proc_9_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(proc_9_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(proc_9_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(proc_9_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(proc_9_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(proc_9_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(proc_9_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(proc_9_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(proc_9_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(proc_9_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(proc_9_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(proc_9_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(proc_9_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(proc_9_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(proc_9_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(proc_9_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(proc_9_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(proc_9_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(proc_9_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(proc_9_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(proc_9_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(proc_9_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(proc_9_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(proc_9_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(proc_9_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(proc_9_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(proc_9_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(proc_9_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(proc_9_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(proc_9_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(proc_9_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(proc_9_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(proc_9_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(proc_9_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(proc_9_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(proc_9_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(proc_9_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(proc_9_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(proc_9_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(proc_9_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_next_processor_id(proc_9_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_9_io_pipe_phv_out_next_config_id),
    .io_mod_mat_mod_en(proc_9_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_9_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_9_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_9_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_9_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_9_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_9_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_9_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_9_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_9_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_9_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_9_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_9_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_9_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_9_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_9_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_9_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_9_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_9_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_9_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_9_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_9_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_9_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_9_io_mod_exe_mod_data_1)
  );
  ProcessorPISA proc_10 ( // @[pisa.scala 28:25]
    .clock(proc_10_clock),
    .io_pipe_phv_in_data_0(proc_10_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_10_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_10_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_10_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_10_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_10_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_10_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_10_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_10_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_10_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_10_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_10_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_10_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_10_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_10_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_10_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_10_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_10_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_10_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_10_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_10_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_10_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_10_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_10_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_10_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_10_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_10_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_10_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_10_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_10_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_10_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_10_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_10_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_10_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_10_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_10_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_10_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_10_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_10_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_10_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_10_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_10_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_10_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_10_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_10_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_10_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_10_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_10_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_10_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_10_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_10_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_10_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_10_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_10_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_10_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_10_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_10_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_10_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_10_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_10_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_10_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_10_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_10_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_10_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_10_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_10_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_10_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_10_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_10_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_10_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_10_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_10_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_10_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_10_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_10_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_10_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_10_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_10_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_10_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_10_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_10_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_10_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_10_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_10_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_10_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_10_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_10_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_10_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_10_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_10_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_10_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_10_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_10_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_10_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_10_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_10_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_10_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_10_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_10_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_10_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_10_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_10_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_10_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_10_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_10_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_10_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_10_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_10_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_10_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_10_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_10_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_10_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_10_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_10_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_10_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_10_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_10_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_10_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_10_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_10_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_10_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_10_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_10_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_10_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_10_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_10_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_10_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_10_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_10_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_10_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_10_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_10_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_10_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_10_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_10_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_10_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_10_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_10_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_10_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_10_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_10_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_10_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_10_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_10_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_10_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_10_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_10_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_10_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_10_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_10_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_10_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_10_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_10_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_10_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_10_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_10_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_10_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_10_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_10_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_10_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(proc_10_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(proc_10_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(proc_10_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(proc_10_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(proc_10_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(proc_10_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(proc_10_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(proc_10_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(proc_10_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(proc_10_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(proc_10_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(proc_10_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(proc_10_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(proc_10_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(proc_10_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(proc_10_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(proc_10_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(proc_10_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(proc_10_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(proc_10_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(proc_10_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(proc_10_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(proc_10_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(proc_10_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(proc_10_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(proc_10_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(proc_10_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(proc_10_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(proc_10_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(proc_10_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(proc_10_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(proc_10_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(proc_10_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(proc_10_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(proc_10_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(proc_10_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(proc_10_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(proc_10_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(proc_10_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(proc_10_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(proc_10_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(proc_10_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(proc_10_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(proc_10_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(proc_10_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(proc_10_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(proc_10_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(proc_10_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(proc_10_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(proc_10_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(proc_10_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(proc_10_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(proc_10_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(proc_10_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(proc_10_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(proc_10_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(proc_10_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(proc_10_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(proc_10_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(proc_10_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(proc_10_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(proc_10_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(proc_10_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(proc_10_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(proc_10_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(proc_10_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(proc_10_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(proc_10_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(proc_10_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(proc_10_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(proc_10_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(proc_10_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(proc_10_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(proc_10_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(proc_10_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(proc_10_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(proc_10_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(proc_10_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(proc_10_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(proc_10_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(proc_10_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(proc_10_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(proc_10_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(proc_10_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(proc_10_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(proc_10_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(proc_10_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(proc_10_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(proc_10_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(proc_10_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(proc_10_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(proc_10_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(proc_10_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(proc_10_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(proc_10_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(proc_10_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_next_processor_id(proc_10_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_10_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_10_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(proc_10_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_10_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_10_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_10_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_10_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_10_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_10_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_10_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_10_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_10_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_10_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_10_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_10_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_10_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_10_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_10_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_10_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_10_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_10_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_10_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_10_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_10_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_10_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_10_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_10_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_10_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_10_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_10_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_10_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_10_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_10_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_10_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_10_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_10_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_10_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_10_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_10_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_10_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_10_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_10_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_10_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_10_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_10_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_10_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_10_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_10_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_10_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_10_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_10_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_10_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_10_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_10_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_10_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_10_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_10_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_10_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_10_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_10_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_10_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_10_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_10_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_10_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_10_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_10_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_10_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_10_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_10_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_10_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_10_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_10_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_10_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_10_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_10_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_10_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_10_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_10_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_10_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_10_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_10_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_10_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_10_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_10_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_10_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_10_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_10_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_10_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_10_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_10_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_10_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_10_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_10_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_10_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_10_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_10_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_10_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_10_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_10_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_10_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_10_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_10_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_10_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_10_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_10_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_10_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_10_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_10_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_10_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_10_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_10_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_10_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_10_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_10_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_10_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_10_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_10_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_10_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_10_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_10_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_10_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_10_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_10_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_10_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_10_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_10_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_10_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_10_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_10_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_10_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_10_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_10_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_10_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_10_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_10_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_10_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_10_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_10_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_10_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_10_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_10_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_10_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_10_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_10_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_10_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_10_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_10_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_10_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_10_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_10_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_10_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_10_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_10_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_10_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_10_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_10_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_10_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_10_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_10_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_10_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_10_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_10_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(proc_10_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(proc_10_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(proc_10_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(proc_10_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(proc_10_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(proc_10_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(proc_10_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(proc_10_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(proc_10_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(proc_10_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(proc_10_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(proc_10_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(proc_10_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(proc_10_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(proc_10_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(proc_10_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(proc_10_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(proc_10_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(proc_10_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(proc_10_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(proc_10_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(proc_10_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(proc_10_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(proc_10_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(proc_10_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(proc_10_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(proc_10_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(proc_10_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(proc_10_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(proc_10_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(proc_10_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(proc_10_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(proc_10_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(proc_10_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(proc_10_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(proc_10_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(proc_10_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(proc_10_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(proc_10_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(proc_10_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(proc_10_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(proc_10_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(proc_10_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(proc_10_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(proc_10_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(proc_10_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(proc_10_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(proc_10_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(proc_10_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(proc_10_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(proc_10_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(proc_10_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(proc_10_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(proc_10_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(proc_10_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(proc_10_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(proc_10_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(proc_10_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(proc_10_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(proc_10_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(proc_10_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(proc_10_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(proc_10_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(proc_10_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(proc_10_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(proc_10_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(proc_10_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(proc_10_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(proc_10_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(proc_10_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(proc_10_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(proc_10_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(proc_10_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(proc_10_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(proc_10_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(proc_10_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(proc_10_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(proc_10_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(proc_10_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(proc_10_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(proc_10_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(proc_10_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(proc_10_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(proc_10_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(proc_10_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(proc_10_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(proc_10_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(proc_10_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(proc_10_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(proc_10_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(proc_10_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(proc_10_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(proc_10_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(proc_10_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(proc_10_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(proc_10_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_next_processor_id(proc_10_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_10_io_pipe_phv_out_next_config_id),
    .io_mod_mat_mod_en(proc_10_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_10_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_10_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_10_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_10_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_10_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_10_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_10_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_10_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_10_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_10_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_10_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_10_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_10_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_10_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_10_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_10_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_10_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_10_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_10_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_10_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_10_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_10_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_10_io_mod_exe_mod_data_1)
  );
  ProcessorPISA proc_11 ( // @[pisa.scala 28:25]
    .clock(proc_11_clock),
    .io_pipe_phv_in_data_0(proc_11_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_11_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_11_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_11_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_11_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_11_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_11_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_11_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_11_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_11_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_11_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_11_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_11_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_11_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_11_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_11_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_11_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_11_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_11_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_11_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_11_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_11_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_11_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_11_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_11_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_11_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_11_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_11_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_11_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_11_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_11_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_11_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_11_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_11_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_11_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_11_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_11_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_11_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_11_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_11_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_11_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_11_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_11_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_11_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_11_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_11_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_11_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_11_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_11_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_11_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_11_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_11_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_11_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_11_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_11_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_11_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_11_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_11_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_11_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_11_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_11_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_11_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_11_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_11_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_11_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_11_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_11_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_11_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_11_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_11_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_11_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_11_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_11_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_11_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_11_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_11_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_11_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_11_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_11_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_11_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_11_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_11_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_11_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_11_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_11_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_11_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_11_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_11_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_11_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_11_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_11_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_11_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_11_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_11_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_11_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_11_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_11_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_11_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_11_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_11_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_11_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_11_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_11_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_11_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_11_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_11_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_11_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_11_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_11_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_11_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_11_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_11_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_11_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_11_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_11_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_11_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_11_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_11_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_11_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_11_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_11_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_11_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_11_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_11_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_11_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_11_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_11_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_11_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_11_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_11_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_11_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_11_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_11_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_11_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_11_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_11_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_11_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_11_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_11_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_11_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_11_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_11_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_11_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_11_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_11_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_11_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_11_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_11_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_11_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_11_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_11_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_11_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_11_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_11_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_11_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_11_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_11_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_11_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_11_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_11_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(proc_11_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(proc_11_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(proc_11_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(proc_11_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(proc_11_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(proc_11_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(proc_11_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(proc_11_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(proc_11_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(proc_11_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(proc_11_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(proc_11_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(proc_11_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(proc_11_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(proc_11_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(proc_11_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(proc_11_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(proc_11_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(proc_11_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(proc_11_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(proc_11_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(proc_11_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(proc_11_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(proc_11_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(proc_11_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(proc_11_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(proc_11_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(proc_11_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(proc_11_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(proc_11_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(proc_11_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(proc_11_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(proc_11_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(proc_11_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(proc_11_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(proc_11_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(proc_11_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(proc_11_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(proc_11_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(proc_11_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(proc_11_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(proc_11_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(proc_11_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(proc_11_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(proc_11_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(proc_11_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(proc_11_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(proc_11_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(proc_11_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(proc_11_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(proc_11_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(proc_11_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(proc_11_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(proc_11_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(proc_11_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(proc_11_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(proc_11_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(proc_11_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(proc_11_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(proc_11_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(proc_11_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(proc_11_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(proc_11_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(proc_11_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(proc_11_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(proc_11_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(proc_11_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(proc_11_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(proc_11_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(proc_11_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(proc_11_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(proc_11_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(proc_11_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(proc_11_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(proc_11_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(proc_11_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(proc_11_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(proc_11_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(proc_11_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(proc_11_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(proc_11_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(proc_11_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(proc_11_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(proc_11_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(proc_11_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(proc_11_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(proc_11_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(proc_11_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(proc_11_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(proc_11_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(proc_11_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(proc_11_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(proc_11_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(proc_11_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(proc_11_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(proc_11_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_next_processor_id(proc_11_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_11_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_11_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(proc_11_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_11_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_11_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_11_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_11_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_11_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_11_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_11_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_11_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_11_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_11_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_11_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_11_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_11_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_11_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_11_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_11_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_11_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_11_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_11_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_11_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_11_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_11_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_11_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_11_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_11_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_11_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_11_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_11_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_11_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_11_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_11_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_11_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_11_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_11_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_11_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_11_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_11_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_11_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_11_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_11_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_11_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_11_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_11_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_11_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_11_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_11_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_11_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_11_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_11_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_11_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_11_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_11_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_11_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_11_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_11_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_11_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_11_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_11_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_11_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_11_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_11_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_11_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_11_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_11_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_11_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_11_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_11_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_11_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_11_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_11_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_11_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_11_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_11_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_11_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_11_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_11_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_11_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_11_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_11_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_11_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_11_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_11_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_11_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_11_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_11_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_11_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_11_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_11_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_11_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_11_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_11_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_11_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_11_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_11_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_11_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_11_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_11_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_11_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_11_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_11_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_11_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_11_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_11_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_11_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_11_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_11_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_11_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_11_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_11_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_11_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_11_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_11_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_11_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_11_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_11_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_11_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_11_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_11_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_11_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_11_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_11_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_11_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_11_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_11_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_11_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_11_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_11_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_11_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_11_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_11_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_11_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_11_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_11_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_11_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_11_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_11_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_11_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_11_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_11_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_11_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_11_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_11_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_11_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_11_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_11_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_11_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_11_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_11_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_11_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_11_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_11_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_11_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_11_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_11_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_11_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_11_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_11_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_11_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_11_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(proc_11_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(proc_11_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(proc_11_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(proc_11_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(proc_11_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(proc_11_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(proc_11_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(proc_11_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(proc_11_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(proc_11_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(proc_11_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(proc_11_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(proc_11_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(proc_11_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(proc_11_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(proc_11_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(proc_11_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(proc_11_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(proc_11_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(proc_11_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(proc_11_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(proc_11_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(proc_11_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(proc_11_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(proc_11_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(proc_11_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(proc_11_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(proc_11_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(proc_11_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(proc_11_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(proc_11_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(proc_11_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(proc_11_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(proc_11_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(proc_11_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(proc_11_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(proc_11_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(proc_11_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(proc_11_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(proc_11_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(proc_11_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(proc_11_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(proc_11_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(proc_11_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(proc_11_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(proc_11_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(proc_11_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(proc_11_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(proc_11_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(proc_11_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(proc_11_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(proc_11_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(proc_11_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(proc_11_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(proc_11_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(proc_11_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(proc_11_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(proc_11_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(proc_11_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(proc_11_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(proc_11_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(proc_11_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(proc_11_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(proc_11_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(proc_11_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(proc_11_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(proc_11_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(proc_11_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(proc_11_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(proc_11_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(proc_11_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(proc_11_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(proc_11_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(proc_11_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(proc_11_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(proc_11_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(proc_11_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(proc_11_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(proc_11_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(proc_11_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(proc_11_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(proc_11_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(proc_11_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(proc_11_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(proc_11_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(proc_11_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(proc_11_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(proc_11_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(proc_11_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(proc_11_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(proc_11_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(proc_11_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(proc_11_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(proc_11_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(proc_11_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(proc_11_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_next_processor_id(proc_11_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_11_io_pipe_phv_out_next_config_id),
    .io_mod_mat_mod_en(proc_11_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_11_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_11_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_11_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_11_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_11_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_11_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_11_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_11_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_11_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_11_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_11_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_11_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_11_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_11_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_11_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_11_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_11_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_11_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_11_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_11_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_11_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_11_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_11_io_mod_exe_mod_data_1)
  );
  assign io_pipe_phv_out_data_0 = proc_11_io_pipe_phv_out_data_0; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_1 = proc_11_io_pipe_phv_out_data_1; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_2 = proc_11_io_pipe_phv_out_data_2; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_3 = proc_11_io_pipe_phv_out_data_3; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_4 = proc_11_io_pipe_phv_out_data_4; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_5 = proc_11_io_pipe_phv_out_data_5; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_6 = proc_11_io_pipe_phv_out_data_6; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_7 = proc_11_io_pipe_phv_out_data_7; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_8 = proc_11_io_pipe_phv_out_data_8; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_9 = proc_11_io_pipe_phv_out_data_9; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_10 = proc_11_io_pipe_phv_out_data_10; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_11 = proc_11_io_pipe_phv_out_data_11; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_12 = proc_11_io_pipe_phv_out_data_12; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_13 = proc_11_io_pipe_phv_out_data_13; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_14 = proc_11_io_pipe_phv_out_data_14; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_15 = proc_11_io_pipe_phv_out_data_15; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_16 = proc_11_io_pipe_phv_out_data_16; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_17 = proc_11_io_pipe_phv_out_data_17; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_18 = proc_11_io_pipe_phv_out_data_18; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_19 = proc_11_io_pipe_phv_out_data_19; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_20 = proc_11_io_pipe_phv_out_data_20; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_21 = proc_11_io_pipe_phv_out_data_21; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_22 = proc_11_io_pipe_phv_out_data_22; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_23 = proc_11_io_pipe_phv_out_data_23; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_24 = proc_11_io_pipe_phv_out_data_24; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_25 = proc_11_io_pipe_phv_out_data_25; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_26 = proc_11_io_pipe_phv_out_data_26; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_27 = proc_11_io_pipe_phv_out_data_27; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_28 = proc_11_io_pipe_phv_out_data_28; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_29 = proc_11_io_pipe_phv_out_data_29; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_30 = proc_11_io_pipe_phv_out_data_30; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_31 = proc_11_io_pipe_phv_out_data_31; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_32 = proc_11_io_pipe_phv_out_data_32; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_33 = proc_11_io_pipe_phv_out_data_33; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_34 = proc_11_io_pipe_phv_out_data_34; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_35 = proc_11_io_pipe_phv_out_data_35; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_36 = proc_11_io_pipe_phv_out_data_36; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_37 = proc_11_io_pipe_phv_out_data_37; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_38 = proc_11_io_pipe_phv_out_data_38; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_39 = proc_11_io_pipe_phv_out_data_39; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_40 = proc_11_io_pipe_phv_out_data_40; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_41 = proc_11_io_pipe_phv_out_data_41; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_42 = proc_11_io_pipe_phv_out_data_42; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_43 = proc_11_io_pipe_phv_out_data_43; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_44 = proc_11_io_pipe_phv_out_data_44; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_45 = proc_11_io_pipe_phv_out_data_45; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_46 = proc_11_io_pipe_phv_out_data_46; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_47 = proc_11_io_pipe_phv_out_data_47; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_48 = proc_11_io_pipe_phv_out_data_48; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_49 = proc_11_io_pipe_phv_out_data_49; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_50 = proc_11_io_pipe_phv_out_data_50; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_51 = proc_11_io_pipe_phv_out_data_51; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_52 = proc_11_io_pipe_phv_out_data_52; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_53 = proc_11_io_pipe_phv_out_data_53; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_54 = proc_11_io_pipe_phv_out_data_54; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_55 = proc_11_io_pipe_phv_out_data_55; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_56 = proc_11_io_pipe_phv_out_data_56; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_57 = proc_11_io_pipe_phv_out_data_57; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_58 = proc_11_io_pipe_phv_out_data_58; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_59 = proc_11_io_pipe_phv_out_data_59; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_60 = proc_11_io_pipe_phv_out_data_60; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_61 = proc_11_io_pipe_phv_out_data_61; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_62 = proc_11_io_pipe_phv_out_data_62; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_63 = proc_11_io_pipe_phv_out_data_63; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_64 = proc_11_io_pipe_phv_out_data_64; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_65 = proc_11_io_pipe_phv_out_data_65; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_66 = proc_11_io_pipe_phv_out_data_66; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_67 = proc_11_io_pipe_phv_out_data_67; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_68 = proc_11_io_pipe_phv_out_data_68; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_69 = proc_11_io_pipe_phv_out_data_69; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_70 = proc_11_io_pipe_phv_out_data_70; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_71 = proc_11_io_pipe_phv_out_data_71; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_72 = proc_11_io_pipe_phv_out_data_72; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_73 = proc_11_io_pipe_phv_out_data_73; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_74 = proc_11_io_pipe_phv_out_data_74; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_75 = proc_11_io_pipe_phv_out_data_75; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_76 = proc_11_io_pipe_phv_out_data_76; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_77 = proc_11_io_pipe_phv_out_data_77; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_78 = proc_11_io_pipe_phv_out_data_78; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_79 = proc_11_io_pipe_phv_out_data_79; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_80 = proc_11_io_pipe_phv_out_data_80; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_81 = proc_11_io_pipe_phv_out_data_81; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_82 = proc_11_io_pipe_phv_out_data_82; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_83 = proc_11_io_pipe_phv_out_data_83; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_84 = proc_11_io_pipe_phv_out_data_84; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_85 = proc_11_io_pipe_phv_out_data_85; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_86 = proc_11_io_pipe_phv_out_data_86; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_87 = proc_11_io_pipe_phv_out_data_87; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_88 = proc_11_io_pipe_phv_out_data_88; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_89 = proc_11_io_pipe_phv_out_data_89; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_90 = proc_11_io_pipe_phv_out_data_90; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_91 = proc_11_io_pipe_phv_out_data_91; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_92 = proc_11_io_pipe_phv_out_data_92; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_93 = proc_11_io_pipe_phv_out_data_93; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_94 = proc_11_io_pipe_phv_out_data_94; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_95 = proc_11_io_pipe_phv_out_data_95; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_96 = proc_11_io_pipe_phv_out_data_96; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_97 = proc_11_io_pipe_phv_out_data_97; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_98 = proc_11_io_pipe_phv_out_data_98; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_99 = proc_11_io_pipe_phv_out_data_99; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_100 = proc_11_io_pipe_phv_out_data_100; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_101 = proc_11_io_pipe_phv_out_data_101; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_102 = proc_11_io_pipe_phv_out_data_102; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_103 = proc_11_io_pipe_phv_out_data_103; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_104 = proc_11_io_pipe_phv_out_data_104; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_105 = proc_11_io_pipe_phv_out_data_105; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_106 = proc_11_io_pipe_phv_out_data_106; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_107 = proc_11_io_pipe_phv_out_data_107; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_108 = proc_11_io_pipe_phv_out_data_108; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_109 = proc_11_io_pipe_phv_out_data_109; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_110 = proc_11_io_pipe_phv_out_data_110; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_111 = proc_11_io_pipe_phv_out_data_111; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_112 = proc_11_io_pipe_phv_out_data_112; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_113 = proc_11_io_pipe_phv_out_data_113; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_114 = proc_11_io_pipe_phv_out_data_114; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_115 = proc_11_io_pipe_phv_out_data_115; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_116 = proc_11_io_pipe_phv_out_data_116; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_117 = proc_11_io_pipe_phv_out_data_117; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_118 = proc_11_io_pipe_phv_out_data_118; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_119 = proc_11_io_pipe_phv_out_data_119; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_120 = proc_11_io_pipe_phv_out_data_120; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_121 = proc_11_io_pipe_phv_out_data_121; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_122 = proc_11_io_pipe_phv_out_data_122; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_123 = proc_11_io_pipe_phv_out_data_123; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_124 = proc_11_io_pipe_phv_out_data_124; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_125 = proc_11_io_pipe_phv_out_data_125; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_126 = proc_11_io_pipe_phv_out_data_126; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_127 = proc_11_io_pipe_phv_out_data_127; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_128 = proc_11_io_pipe_phv_out_data_128; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_129 = proc_11_io_pipe_phv_out_data_129; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_130 = proc_11_io_pipe_phv_out_data_130; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_131 = proc_11_io_pipe_phv_out_data_131; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_132 = proc_11_io_pipe_phv_out_data_132; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_133 = proc_11_io_pipe_phv_out_data_133; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_134 = proc_11_io_pipe_phv_out_data_134; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_135 = proc_11_io_pipe_phv_out_data_135; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_136 = proc_11_io_pipe_phv_out_data_136; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_137 = proc_11_io_pipe_phv_out_data_137; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_138 = proc_11_io_pipe_phv_out_data_138; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_139 = proc_11_io_pipe_phv_out_data_139; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_140 = proc_11_io_pipe_phv_out_data_140; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_141 = proc_11_io_pipe_phv_out_data_141; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_142 = proc_11_io_pipe_phv_out_data_142; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_143 = proc_11_io_pipe_phv_out_data_143; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_144 = proc_11_io_pipe_phv_out_data_144; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_145 = proc_11_io_pipe_phv_out_data_145; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_146 = proc_11_io_pipe_phv_out_data_146; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_147 = proc_11_io_pipe_phv_out_data_147; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_148 = proc_11_io_pipe_phv_out_data_148; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_149 = proc_11_io_pipe_phv_out_data_149; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_150 = proc_11_io_pipe_phv_out_data_150; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_151 = proc_11_io_pipe_phv_out_data_151; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_152 = proc_11_io_pipe_phv_out_data_152; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_153 = proc_11_io_pipe_phv_out_data_153; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_154 = proc_11_io_pipe_phv_out_data_154; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_155 = proc_11_io_pipe_phv_out_data_155; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_156 = proc_11_io_pipe_phv_out_data_156; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_157 = proc_11_io_pipe_phv_out_data_157; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_158 = proc_11_io_pipe_phv_out_data_158; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_159 = proc_11_io_pipe_phv_out_data_159; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_160 = proc_11_io_pipe_phv_out_data_160; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_161 = proc_11_io_pipe_phv_out_data_161; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_162 = proc_11_io_pipe_phv_out_data_162; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_163 = proc_11_io_pipe_phv_out_data_163; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_164 = proc_11_io_pipe_phv_out_data_164; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_165 = proc_11_io_pipe_phv_out_data_165; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_166 = proc_11_io_pipe_phv_out_data_166; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_167 = proc_11_io_pipe_phv_out_data_167; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_168 = proc_11_io_pipe_phv_out_data_168; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_169 = proc_11_io_pipe_phv_out_data_169; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_170 = proc_11_io_pipe_phv_out_data_170; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_171 = proc_11_io_pipe_phv_out_data_171; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_172 = proc_11_io_pipe_phv_out_data_172; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_173 = proc_11_io_pipe_phv_out_data_173; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_174 = proc_11_io_pipe_phv_out_data_174; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_175 = proc_11_io_pipe_phv_out_data_175; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_176 = proc_11_io_pipe_phv_out_data_176; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_177 = proc_11_io_pipe_phv_out_data_177; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_178 = proc_11_io_pipe_phv_out_data_178; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_179 = proc_11_io_pipe_phv_out_data_179; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_180 = proc_11_io_pipe_phv_out_data_180; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_181 = proc_11_io_pipe_phv_out_data_181; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_182 = proc_11_io_pipe_phv_out_data_182; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_183 = proc_11_io_pipe_phv_out_data_183; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_184 = proc_11_io_pipe_phv_out_data_184; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_185 = proc_11_io_pipe_phv_out_data_185; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_186 = proc_11_io_pipe_phv_out_data_186; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_187 = proc_11_io_pipe_phv_out_data_187; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_188 = proc_11_io_pipe_phv_out_data_188; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_189 = proc_11_io_pipe_phv_out_data_189; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_190 = proc_11_io_pipe_phv_out_data_190; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_191 = proc_11_io_pipe_phv_out_data_191; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_192 = proc_11_io_pipe_phv_out_data_192; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_193 = proc_11_io_pipe_phv_out_data_193; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_194 = proc_11_io_pipe_phv_out_data_194; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_195 = proc_11_io_pipe_phv_out_data_195; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_196 = proc_11_io_pipe_phv_out_data_196; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_197 = proc_11_io_pipe_phv_out_data_197; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_198 = proc_11_io_pipe_phv_out_data_198; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_199 = proc_11_io_pipe_phv_out_data_199; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_200 = proc_11_io_pipe_phv_out_data_200; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_201 = proc_11_io_pipe_phv_out_data_201; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_202 = proc_11_io_pipe_phv_out_data_202; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_203 = proc_11_io_pipe_phv_out_data_203; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_204 = proc_11_io_pipe_phv_out_data_204; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_205 = proc_11_io_pipe_phv_out_data_205; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_206 = proc_11_io_pipe_phv_out_data_206; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_207 = proc_11_io_pipe_phv_out_data_207; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_208 = proc_11_io_pipe_phv_out_data_208; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_209 = proc_11_io_pipe_phv_out_data_209; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_210 = proc_11_io_pipe_phv_out_data_210; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_211 = proc_11_io_pipe_phv_out_data_211; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_212 = proc_11_io_pipe_phv_out_data_212; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_213 = proc_11_io_pipe_phv_out_data_213; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_214 = proc_11_io_pipe_phv_out_data_214; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_215 = proc_11_io_pipe_phv_out_data_215; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_216 = proc_11_io_pipe_phv_out_data_216; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_217 = proc_11_io_pipe_phv_out_data_217; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_218 = proc_11_io_pipe_phv_out_data_218; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_219 = proc_11_io_pipe_phv_out_data_219; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_220 = proc_11_io_pipe_phv_out_data_220; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_221 = proc_11_io_pipe_phv_out_data_221; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_222 = proc_11_io_pipe_phv_out_data_222; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_223 = proc_11_io_pipe_phv_out_data_223; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_224 = proc_11_io_pipe_phv_out_data_224; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_225 = proc_11_io_pipe_phv_out_data_225; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_226 = proc_11_io_pipe_phv_out_data_226; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_227 = proc_11_io_pipe_phv_out_data_227; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_228 = proc_11_io_pipe_phv_out_data_228; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_229 = proc_11_io_pipe_phv_out_data_229; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_230 = proc_11_io_pipe_phv_out_data_230; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_231 = proc_11_io_pipe_phv_out_data_231; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_232 = proc_11_io_pipe_phv_out_data_232; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_233 = proc_11_io_pipe_phv_out_data_233; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_234 = proc_11_io_pipe_phv_out_data_234; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_235 = proc_11_io_pipe_phv_out_data_235; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_236 = proc_11_io_pipe_phv_out_data_236; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_237 = proc_11_io_pipe_phv_out_data_237; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_238 = proc_11_io_pipe_phv_out_data_238; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_239 = proc_11_io_pipe_phv_out_data_239; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_240 = proc_11_io_pipe_phv_out_data_240; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_241 = proc_11_io_pipe_phv_out_data_241; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_242 = proc_11_io_pipe_phv_out_data_242; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_243 = proc_11_io_pipe_phv_out_data_243; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_244 = proc_11_io_pipe_phv_out_data_244; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_245 = proc_11_io_pipe_phv_out_data_245; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_246 = proc_11_io_pipe_phv_out_data_246; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_247 = proc_11_io_pipe_phv_out_data_247; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_248 = proc_11_io_pipe_phv_out_data_248; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_249 = proc_11_io_pipe_phv_out_data_249; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_250 = proc_11_io_pipe_phv_out_data_250; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_251 = proc_11_io_pipe_phv_out_data_251; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_252 = proc_11_io_pipe_phv_out_data_252; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_253 = proc_11_io_pipe_phv_out_data_253; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_254 = proc_11_io_pipe_phv_out_data_254; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_255 = proc_11_io_pipe_phv_out_data_255; // @[pisa.scala 42:52]
  assign init_clock = clock;
  assign init_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_96 = io_pipe_phv_in_data_96; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_97 = io_pipe_phv_in_data_97; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_98 = io_pipe_phv_in_data_98; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_99 = io_pipe_phv_in_data_99; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_100 = io_pipe_phv_in_data_100; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_101 = io_pipe_phv_in_data_101; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_102 = io_pipe_phv_in_data_102; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_103 = io_pipe_phv_in_data_103; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_104 = io_pipe_phv_in_data_104; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_105 = io_pipe_phv_in_data_105; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_106 = io_pipe_phv_in_data_106; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_107 = io_pipe_phv_in_data_107; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_108 = io_pipe_phv_in_data_108; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_109 = io_pipe_phv_in_data_109; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_110 = io_pipe_phv_in_data_110; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_111 = io_pipe_phv_in_data_111; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_112 = io_pipe_phv_in_data_112; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_113 = io_pipe_phv_in_data_113; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_114 = io_pipe_phv_in_data_114; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_115 = io_pipe_phv_in_data_115; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_116 = io_pipe_phv_in_data_116; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_117 = io_pipe_phv_in_data_117; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_118 = io_pipe_phv_in_data_118; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_119 = io_pipe_phv_in_data_119; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_120 = io_pipe_phv_in_data_120; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_121 = io_pipe_phv_in_data_121; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_122 = io_pipe_phv_in_data_122; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_123 = io_pipe_phv_in_data_123; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_124 = io_pipe_phv_in_data_124; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_125 = io_pipe_phv_in_data_125; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_126 = io_pipe_phv_in_data_126; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_127 = io_pipe_phv_in_data_127; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_128 = io_pipe_phv_in_data_128; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_129 = io_pipe_phv_in_data_129; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_130 = io_pipe_phv_in_data_130; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_131 = io_pipe_phv_in_data_131; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_132 = io_pipe_phv_in_data_132; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_133 = io_pipe_phv_in_data_133; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_134 = io_pipe_phv_in_data_134; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_135 = io_pipe_phv_in_data_135; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_136 = io_pipe_phv_in_data_136; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_137 = io_pipe_phv_in_data_137; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_138 = io_pipe_phv_in_data_138; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_139 = io_pipe_phv_in_data_139; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_140 = io_pipe_phv_in_data_140; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_141 = io_pipe_phv_in_data_141; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_142 = io_pipe_phv_in_data_142; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_143 = io_pipe_phv_in_data_143; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_144 = io_pipe_phv_in_data_144; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_145 = io_pipe_phv_in_data_145; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_146 = io_pipe_phv_in_data_146; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_147 = io_pipe_phv_in_data_147; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_148 = io_pipe_phv_in_data_148; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_149 = io_pipe_phv_in_data_149; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_150 = io_pipe_phv_in_data_150; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_151 = io_pipe_phv_in_data_151; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_152 = io_pipe_phv_in_data_152; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_153 = io_pipe_phv_in_data_153; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_154 = io_pipe_phv_in_data_154; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_155 = io_pipe_phv_in_data_155; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_156 = io_pipe_phv_in_data_156; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_157 = io_pipe_phv_in_data_157; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_158 = io_pipe_phv_in_data_158; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_159 = io_pipe_phv_in_data_159; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_160 = io_pipe_phv_in_data_160; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_161 = io_pipe_phv_in_data_161; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_162 = io_pipe_phv_in_data_162; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_163 = io_pipe_phv_in_data_163; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_164 = io_pipe_phv_in_data_164; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_165 = io_pipe_phv_in_data_165; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_166 = io_pipe_phv_in_data_166; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_167 = io_pipe_phv_in_data_167; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_168 = io_pipe_phv_in_data_168; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_169 = io_pipe_phv_in_data_169; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_170 = io_pipe_phv_in_data_170; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_171 = io_pipe_phv_in_data_171; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_172 = io_pipe_phv_in_data_172; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_173 = io_pipe_phv_in_data_173; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_174 = io_pipe_phv_in_data_174; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_175 = io_pipe_phv_in_data_175; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_176 = io_pipe_phv_in_data_176; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_177 = io_pipe_phv_in_data_177; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_178 = io_pipe_phv_in_data_178; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_179 = io_pipe_phv_in_data_179; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_180 = io_pipe_phv_in_data_180; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_181 = io_pipe_phv_in_data_181; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_182 = io_pipe_phv_in_data_182; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_183 = io_pipe_phv_in_data_183; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_184 = io_pipe_phv_in_data_184; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_185 = io_pipe_phv_in_data_185; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_186 = io_pipe_phv_in_data_186; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_187 = io_pipe_phv_in_data_187; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_188 = io_pipe_phv_in_data_188; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_189 = io_pipe_phv_in_data_189; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_190 = io_pipe_phv_in_data_190; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_191 = io_pipe_phv_in_data_191; // @[pisa.scala 20:25]
  assign PAR_clock = clock;
  assign PAR_io_pipe_phv_in_data_0 = init_io_pipe_phv_out_data_0; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_1 = init_io_pipe_phv_out_data_1; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_2 = init_io_pipe_phv_out_data_2; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_3 = init_io_pipe_phv_out_data_3; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_4 = init_io_pipe_phv_out_data_4; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_5 = init_io_pipe_phv_out_data_5; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_6 = init_io_pipe_phv_out_data_6; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_7 = init_io_pipe_phv_out_data_7; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_8 = init_io_pipe_phv_out_data_8; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_9 = init_io_pipe_phv_out_data_9; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_10 = init_io_pipe_phv_out_data_10; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_11 = init_io_pipe_phv_out_data_11; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_12 = init_io_pipe_phv_out_data_12; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_13 = init_io_pipe_phv_out_data_13; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_14 = init_io_pipe_phv_out_data_14; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_15 = init_io_pipe_phv_out_data_15; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_16 = init_io_pipe_phv_out_data_16; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_17 = init_io_pipe_phv_out_data_17; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_18 = init_io_pipe_phv_out_data_18; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_19 = init_io_pipe_phv_out_data_19; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_20 = init_io_pipe_phv_out_data_20; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_21 = init_io_pipe_phv_out_data_21; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_22 = init_io_pipe_phv_out_data_22; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_23 = init_io_pipe_phv_out_data_23; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_24 = init_io_pipe_phv_out_data_24; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_25 = init_io_pipe_phv_out_data_25; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_26 = init_io_pipe_phv_out_data_26; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_27 = init_io_pipe_phv_out_data_27; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_28 = init_io_pipe_phv_out_data_28; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_29 = init_io_pipe_phv_out_data_29; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_30 = init_io_pipe_phv_out_data_30; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_31 = init_io_pipe_phv_out_data_31; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_32 = init_io_pipe_phv_out_data_32; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_33 = init_io_pipe_phv_out_data_33; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_34 = init_io_pipe_phv_out_data_34; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_35 = init_io_pipe_phv_out_data_35; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_36 = init_io_pipe_phv_out_data_36; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_37 = init_io_pipe_phv_out_data_37; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_38 = init_io_pipe_phv_out_data_38; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_39 = init_io_pipe_phv_out_data_39; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_40 = init_io_pipe_phv_out_data_40; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_41 = init_io_pipe_phv_out_data_41; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_42 = init_io_pipe_phv_out_data_42; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_43 = init_io_pipe_phv_out_data_43; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_44 = init_io_pipe_phv_out_data_44; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_45 = init_io_pipe_phv_out_data_45; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_46 = init_io_pipe_phv_out_data_46; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_47 = init_io_pipe_phv_out_data_47; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_48 = init_io_pipe_phv_out_data_48; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_49 = init_io_pipe_phv_out_data_49; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_50 = init_io_pipe_phv_out_data_50; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_51 = init_io_pipe_phv_out_data_51; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_52 = init_io_pipe_phv_out_data_52; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_53 = init_io_pipe_phv_out_data_53; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_54 = init_io_pipe_phv_out_data_54; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_55 = init_io_pipe_phv_out_data_55; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_56 = init_io_pipe_phv_out_data_56; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_57 = init_io_pipe_phv_out_data_57; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_58 = init_io_pipe_phv_out_data_58; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_59 = init_io_pipe_phv_out_data_59; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_60 = init_io_pipe_phv_out_data_60; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_61 = init_io_pipe_phv_out_data_61; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_62 = init_io_pipe_phv_out_data_62; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_63 = init_io_pipe_phv_out_data_63; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_64 = init_io_pipe_phv_out_data_64; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_65 = init_io_pipe_phv_out_data_65; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_66 = init_io_pipe_phv_out_data_66; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_67 = init_io_pipe_phv_out_data_67; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_68 = init_io_pipe_phv_out_data_68; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_69 = init_io_pipe_phv_out_data_69; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_70 = init_io_pipe_phv_out_data_70; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_71 = init_io_pipe_phv_out_data_71; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_72 = init_io_pipe_phv_out_data_72; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_73 = init_io_pipe_phv_out_data_73; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_74 = init_io_pipe_phv_out_data_74; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_75 = init_io_pipe_phv_out_data_75; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_76 = init_io_pipe_phv_out_data_76; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_77 = init_io_pipe_phv_out_data_77; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_78 = init_io_pipe_phv_out_data_78; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_79 = init_io_pipe_phv_out_data_79; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_80 = init_io_pipe_phv_out_data_80; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_81 = init_io_pipe_phv_out_data_81; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_82 = init_io_pipe_phv_out_data_82; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_83 = init_io_pipe_phv_out_data_83; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_84 = init_io_pipe_phv_out_data_84; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_85 = init_io_pipe_phv_out_data_85; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_86 = init_io_pipe_phv_out_data_86; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_87 = init_io_pipe_phv_out_data_87; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_88 = init_io_pipe_phv_out_data_88; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_89 = init_io_pipe_phv_out_data_89; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_90 = init_io_pipe_phv_out_data_90; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_91 = init_io_pipe_phv_out_data_91; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_92 = init_io_pipe_phv_out_data_92; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_93 = init_io_pipe_phv_out_data_93; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_94 = init_io_pipe_phv_out_data_94; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_95 = init_io_pipe_phv_out_data_95; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_96 = init_io_pipe_phv_out_data_96; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_97 = init_io_pipe_phv_out_data_97; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_98 = init_io_pipe_phv_out_data_98; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_99 = init_io_pipe_phv_out_data_99; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_100 = init_io_pipe_phv_out_data_100; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_101 = init_io_pipe_phv_out_data_101; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_102 = init_io_pipe_phv_out_data_102; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_103 = init_io_pipe_phv_out_data_103; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_104 = init_io_pipe_phv_out_data_104; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_105 = init_io_pipe_phv_out_data_105; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_106 = init_io_pipe_phv_out_data_106; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_107 = init_io_pipe_phv_out_data_107; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_108 = init_io_pipe_phv_out_data_108; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_109 = init_io_pipe_phv_out_data_109; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_110 = init_io_pipe_phv_out_data_110; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_111 = init_io_pipe_phv_out_data_111; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_112 = init_io_pipe_phv_out_data_112; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_113 = init_io_pipe_phv_out_data_113; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_114 = init_io_pipe_phv_out_data_114; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_115 = init_io_pipe_phv_out_data_115; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_116 = init_io_pipe_phv_out_data_116; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_117 = init_io_pipe_phv_out_data_117; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_118 = init_io_pipe_phv_out_data_118; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_119 = init_io_pipe_phv_out_data_119; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_120 = init_io_pipe_phv_out_data_120; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_121 = init_io_pipe_phv_out_data_121; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_122 = init_io_pipe_phv_out_data_122; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_123 = init_io_pipe_phv_out_data_123; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_124 = init_io_pipe_phv_out_data_124; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_125 = init_io_pipe_phv_out_data_125; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_126 = init_io_pipe_phv_out_data_126; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_127 = init_io_pipe_phv_out_data_127; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_128 = init_io_pipe_phv_out_data_128; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_129 = init_io_pipe_phv_out_data_129; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_130 = init_io_pipe_phv_out_data_130; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_131 = init_io_pipe_phv_out_data_131; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_132 = init_io_pipe_phv_out_data_132; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_133 = init_io_pipe_phv_out_data_133; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_134 = init_io_pipe_phv_out_data_134; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_135 = init_io_pipe_phv_out_data_135; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_136 = init_io_pipe_phv_out_data_136; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_137 = init_io_pipe_phv_out_data_137; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_138 = init_io_pipe_phv_out_data_138; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_139 = init_io_pipe_phv_out_data_139; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_140 = init_io_pipe_phv_out_data_140; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_141 = init_io_pipe_phv_out_data_141; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_142 = init_io_pipe_phv_out_data_142; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_143 = init_io_pipe_phv_out_data_143; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_144 = init_io_pipe_phv_out_data_144; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_145 = init_io_pipe_phv_out_data_145; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_146 = init_io_pipe_phv_out_data_146; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_147 = init_io_pipe_phv_out_data_147; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_148 = init_io_pipe_phv_out_data_148; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_149 = init_io_pipe_phv_out_data_149; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_150 = init_io_pipe_phv_out_data_150; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_151 = init_io_pipe_phv_out_data_151; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_152 = init_io_pipe_phv_out_data_152; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_153 = init_io_pipe_phv_out_data_153; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_154 = init_io_pipe_phv_out_data_154; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_155 = init_io_pipe_phv_out_data_155; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_156 = init_io_pipe_phv_out_data_156; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_157 = init_io_pipe_phv_out_data_157; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_158 = init_io_pipe_phv_out_data_158; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_159 = init_io_pipe_phv_out_data_159; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_160 = init_io_pipe_phv_out_data_160; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_161 = init_io_pipe_phv_out_data_161; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_162 = init_io_pipe_phv_out_data_162; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_163 = init_io_pipe_phv_out_data_163; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_164 = init_io_pipe_phv_out_data_164; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_165 = init_io_pipe_phv_out_data_165; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_166 = init_io_pipe_phv_out_data_166; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_167 = init_io_pipe_phv_out_data_167; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_168 = init_io_pipe_phv_out_data_168; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_169 = init_io_pipe_phv_out_data_169; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_170 = init_io_pipe_phv_out_data_170; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_171 = init_io_pipe_phv_out_data_171; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_172 = init_io_pipe_phv_out_data_172; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_173 = init_io_pipe_phv_out_data_173; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_174 = init_io_pipe_phv_out_data_174; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_175 = init_io_pipe_phv_out_data_175; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_176 = init_io_pipe_phv_out_data_176; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_177 = init_io_pipe_phv_out_data_177; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_178 = init_io_pipe_phv_out_data_178; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_179 = init_io_pipe_phv_out_data_179; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_180 = init_io_pipe_phv_out_data_180; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_181 = init_io_pipe_phv_out_data_181; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_182 = init_io_pipe_phv_out_data_182; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_183 = init_io_pipe_phv_out_data_183; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_184 = init_io_pipe_phv_out_data_184; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_185 = init_io_pipe_phv_out_data_185; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_186 = init_io_pipe_phv_out_data_186; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_187 = init_io_pipe_phv_out_data_187; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_188 = init_io_pipe_phv_out_data_188; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_189 = init_io_pipe_phv_out_data_189; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_190 = init_io_pipe_phv_out_data_190; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_191 = init_io_pipe_phv_out_data_191; // @[pisa.scala 24:24]
  assign PAR_io_mod_en = io_mod_par_mod_en; // @[pisa.scala 25:16]
  assign PAR_io_mod_last_mau_id_mod = io_mod_par_mod_last_mau_id_mod; // @[pisa.scala 25:16]
  assign PAR_io_mod_last_mau_id = io_mod_par_mod_last_mau_id; // @[pisa.scala 25:16]
  assign PAR_io_mod_cs = io_mod_par_mod_cs; // @[pisa.scala 25:16]
  assign PAR_io_mod_module_mod_state_id_mod = io_mod_par_mod_module_mod_state_id_mod; // @[pisa.scala 25:16]
  assign PAR_io_mod_module_mod_state_id = io_mod_par_mod_module_mod_state_id; // @[pisa.scala 25:16]
  assign PAR_io_mod_module_mod_sram_w_cs = io_mod_par_mod_module_mod_sram_w_cs; // @[pisa.scala 25:16]
  assign PAR_io_mod_module_mod_sram_w_en = io_mod_par_mod_module_mod_sram_w_en; // @[pisa.scala 25:16]
  assign PAR_io_mod_module_mod_sram_w_addr = io_mod_par_mod_module_mod_sram_w_addr; // @[pisa.scala 25:16]
  assign PAR_io_mod_module_mod_sram_w_data = io_mod_par_mod_module_mod_sram_w_data; // @[pisa.scala 25:16]
  assign proc_0_clock = clock;
  assign proc_0_io_pipe_phv_in_data_0 = PAR_io_pipe_phv_out_data_0; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_1 = PAR_io_pipe_phv_out_data_1; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_2 = PAR_io_pipe_phv_out_data_2; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_3 = PAR_io_pipe_phv_out_data_3; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_4 = PAR_io_pipe_phv_out_data_4; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_5 = PAR_io_pipe_phv_out_data_5; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_6 = PAR_io_pipe_phv_out_data_6; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_7 = PAR_io_pipe_phv_out_data_7; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_8 = PAR_io_pipe_phv_out_data_8; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_9 = PAR_io_pipe_phv_out_data_9; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_10 = PAR_io_pipe_phv_out_data_10; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_11 = PAR_io_pipe_phv_out_data_11; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_12 = PAR_io_pipe_phv_out_data_12; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_13 = PAR_io_pipe_phv_out_data_13; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_14 = PAR_io_pipe_phv_out_data_14; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_15 = PAR_io_pipe_phv_out_data_15; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_16 = PAR_io_pipe_phv_out_data_16; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_17 = PAR_io_pipe_phv_out_data_17; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_18 = PAR_io_pipe_phv_out_data_18; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_19 = PAR_io_pipe_phv_out_data_19; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_20 = PAR_io_pipe_phv_out_data_20; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_21 = PAR_io_pipe_phv_out_data_21; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_22 = PAR_io_pipe_phv_out_data_22; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_23 = PAR_io_pipe_phv_out_data_23; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_24 = PAR_io_pipe_phv_out_data_24; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_25 = PAR_io_pipe_phv_out_data_25; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_26 = PAR_io_pipe_phv_out_data_26; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_27 = PAR_io_pipe_phv_out_data_27; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_28 = PAR_io_pipe_phv_out_data_28; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_29 = PAR_io_pipe_phv_out_data_29; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_30 = PAR_io_pipe_phv_out_data_30; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_31 = PAR_io_pipe_phv_out_data_31; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_32 = PAR_io_pipe_phv_out_data_32; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_33 = PAR_io_pipe_phv_out_data_33; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_34 = PAR_io_pipe_phv_out_data_34; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_35 = PAR_io_pipe_phv_out_data_35; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_36 = PAR_io_pipe_phv_out_data_36; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_37 = PAR_io_pipe_phv_out_data_37; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_38 = PAR_io_pipe_phv_out_data_38; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_39 = PAR_io_pipe_phv_out_data_39; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_40 = PAR_io_pipe_phv_out_data_40; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_41 = PAR_io_pipe_phv_out_data_41; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_42 = PAR_io_pipe_phv_out_data_42; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_43 = PAR_io_pipe_phv_out_data_43; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_44 = PAR_io_pipe_phv_out_data_44; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_45 = PAR_io_pipe_phv_out_data_45; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_46 = PAR_io_pipe_phv_out_data_46; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_47 = PAR_io_pipe_phv_out_data_47; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_48 = PAR_io_pipe_phv_out_data_48; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_49 = PAR_io_pipe_phv_out_data_49; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_50 = PAR_io_pipe_phv_out_data_50; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_51 = PAR_io_pipe_phv_out_data_51; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_52 = PAR_io_pipe_phv_out_data_52; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_53 = PAR_io_pipe_phv_out_data_53; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_54 = PAR_io_pipe_phv_out_data_54; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_55 = PAR_io_pipe_phv_out_data_55; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_56 = PAR_io_pipe_phv_out_data_56; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_57 = PAR_io_pipe_phv_out_data_57; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_58 = PAR_io_pipe_phv_out_data_58; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_59 = PAR_io_pipe_phv_out_data_59; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_60 = PAR_io_pipe_phv_out_data_60; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_61 = PAR_io_pipe_phv_out_data_61; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_62 = PAR_io_pipe_phv_out_data_62; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_63 = PAR_io_pipe_phv_out_data_63; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_64 = PAR_io_pipe_phv_out_data_64; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_65 = PAR_io_pipe_phv_out_data_65; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_66 = PAR_io_pipe_phv_out_data_66; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_67 = PAR_io_pipe_phv_out_data_67; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_68 = PAR_io_pipe_phv_out_data_68; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_69 = PAR_io_pipe_phv_out_data_69; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_70 = PAR_io_pipe_phv_out_data_70; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_71 = PAR_io_pipe_phv_out_data_71; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_72 = PAR_io_pipe_phv_out_data_72; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_73 = PAR_io_pipe_phv_out_data_73; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_74 = PAR_io_pipe_phv_out_data_74; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_75 = PAR_io_pipe_phv_out_data_75; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_76 = PAR_io_pipe_phv_out_data_76; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_77 = PAR_io_pipe_phv_out_data_77; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_78 = PAR_io_pipe_phv_out_data_78; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_79 = PAR_io_pipe_phv_out_data_79; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_80 = PAR_io_pipe_phv_out_data_80; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_81 = PAR_io_pipe_phv_out_data_81; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_82 = PAR_io_pipe_phv_out_data_82; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_83 = PAR_io_pipe_phv_out_data_83; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_84 = PAR_io_pipe_phv_out_data_84; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_85 = PAR_io_pipe_phv_out_data_85; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_86 = PAR_io_pipe_phv_out_data_86; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_87 = PAR_io_pipe_phv_out_data_87; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_88 = PAR_io_pipe_phv_out_data_88; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_89 = PAR_io_pipe_phv_out_data_89; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_90 = PAR_io_pipe_phv_out_data_90; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_91 = PAR_io_pipe_phv_out_data_91; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_92 = PAR_io_pipe_phv_out_data_92; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_93 = PAR_io_pipe_phv_out_data_93; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_94 = PAR_io_pipe_phv_out_data_94; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_95 = PAR_io_pipe_phv_out_data_95; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_96 = PAR_io_pipe_phv_out_data_96; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_97 = PAR_io_pipe_phv_out_data_97; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_98 = PAR_io_pipe_phv_out_data_98; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_99 = PAR_io_pipe_phv_out_data_99; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_100 = PAR_io_pipe_phv_out_data_100; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_101 = PAR_io_pipe_phv_out_data_101; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_102 = PAR_io_pipe_phv_out_data_102; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_103 = PAR_io_pipe_phv_out_data_103; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_104 = PAR_io_pipe_phv_out_data_104; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_105 = PAR_io_pipe_phv_out_data_105; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_106 = PAR_io_pipe_phv_out_data_106; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_107 = PAR_io_pipe_phv_out_data_107; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_108 = PAR_io_pipe_phv_out_data_108; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_109 = PAR_io_pipe_phv_out_data_109; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_110 = PAR_io_pipe_phv_out_data_110; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_111 = PAR_io_pipe_phv_out_data_111; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_112 = PAR_io_pipe_phv_out_data_112; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_113 = PAR_io_pipe_phv_out_data_113; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_114 = PAR_io_pipe_phv_out_data_114; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_115 = PAR_io_pipe_phv_out_data_115; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_116 = PAR_io_pipe_phv_out_data_116; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_117 = PAR_io_pipe_phv_out_data_117; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_118 = PAR_io_pipe_phv_out_data_118; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_119 = PAR_io_pipe_phv_out_data_119; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_120 = PAR_io_pipe_phv_out_data_120; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_121 = PAR_io_pipe_phv_out_data_121; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_122 = PAR_io_pipe_phv_out_data_122; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_123 = PAR_io_pipe_phv_out_data_123; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_124 = PAR_io_pipe_phv_out_data_124; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_125 = PAR_io_pipe_phv_out_data_125; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_126 = PAR_io_pipe_phv_out_data_126; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_127 = PAR_io_pipe_phv_out_data_127; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_128 = PAR_io_pipe_phv_out_data_128; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_129 = PAR_io_pipe_phv_out_data_129; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_130 = PAR_io_pipe_phv_out_data_130; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_131 = PAR_io_pipe_phv_out_data_131; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_132 = PAR_io_pipe_phv_out_data_132; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_133 = PAR_io_pipe_phv_out_data_133; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_134 = PAR_io_pipe_phv_out_data_134; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_135 = PAR_io_pipe_phv_out_data_135; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_136 = PAR_io_pipe_phv_out_data_136; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_137 = PAR_io_pipe_phv_out_data_137; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_138 = PAR_io_pipe_phv_out_data_138; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_139 = PAR_io_pipe_phv_out_data_139; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_140 = PAR_io_pipe_phv_out_data_140; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_141 = PAR_io_pipe_phv_out_data_141; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_142 = PAR_io_pipe_phv_out_data_142; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_143 = PAR_io_pipe_phv_out_data_143; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_144 = PAR_io_pipe_phv_out_data_144; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_145 = PAR_io_pipe_phv_out_data_145; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_146 = PAR_io_pipe_phv_out_data_146; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_147 = PAR_io_pipe_phv_out_data_147; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_148 = PAR_io_pipe_phv_out_data_148; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_149 = PAR_io_pipe_phv_out_data_149; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_150 = PAR_io_pipe_phv_out_data_150; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_151 = PAR_io_pipe_phv_out_data_151; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_152 = PAR_io_pipe_phv_out_data_152; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_153 = PAR_io_pipe_phv_out_data_153; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_154 = PAR_io_pipe_phv_out_data_154; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_155 = PAR_io_pipe_phv_out_data_155; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_156 = PAR_io_pipe_phv_out_data_156; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_157 = PAR_io_pipe_phv_out_data_157; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_158 = PAR_io_pipe_phv_out_data_158; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_159 = PAR_io_pipe_phv_out_data_159; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_160 = PAR_io_pipe_phv_out_data_160; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_161 = PAR_io_pipe_phv_out_data_161; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_162 = PAR_io_pipe_phv_out_data_162; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_163 = PAR_io_pipe_phv_out_data_163; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_164 = PAR_io_pipe_phv_out_data_164; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_165 = PAR_io_pipe_phv_out_data_165; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_166 = PAR_io_pipe_phv_out_data_166; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_167 = PAR_io_pipe_phv_out_data_167; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_168 = PAR_io_pipe_phv_out_data_168; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_169 = PAR_io_pipe_phv_out_data_169; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_170 = PAR_io_pipe_phv_out_data_170; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_171 = PAR_io_pipe_phv_out_data_171; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_172 = PAR_io_pipe_phv_out_data_172; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_173 = PAR_io_pipe_phv_out_data_173; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_174 = PAR_io_pipe_phv_out_data_174; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_175 = PAR_io_pipe_phv_out_data_175; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_176 = PAR_io_pipe_phv_out_data_176; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_177 = PAR_io_pipe_phv_out_data_177; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_178 = PAR_io_pipe_phv_out_data_178; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_179 = PAR_io_pipe_phv_out_data_179; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_180 = PAR_io_pipe_phv_out_data_180; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_181 = PAR_io_pipe_phv_out_data_181; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_182 = PAR_io_pipe_phv_out_data_182; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_183 = PAR_io_pipe_phv_out_data_183; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_184 = PAR_io_pipe_phv_out_data_184; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_185 = PAR_io_pipe_phv_out_data_185; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_186 = PAR_io_pipe_phv_out_data_186; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_187 = PAR_io_pipe_phv_out_data_187; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_188 = PAR_io_pipe_phv_out_data_188; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_189 = PAR_io_pipe_phv_out_data_189; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_190 = PAR_io_pipe_phv_out_data_190; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_191 = PAR_io_pipe_phv_out_data_191; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_192 = PAR_io_pipe_phv_out_data_192; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_193 = PAR_io_pipe_phv_out_data_193; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_194 = PAR_io_pipe_phv_out_data_194; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_195 = PAR_io_pipe_phv_out_data_195; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_196 = PAR_io_pipe_phv_out_data_196; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_197 = PAR_io_pipe_phv_out_data_197; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_198 = PAR_io_pipe_phv_out_data_198; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_199 = PAR_io_pipe_phv_out_data_199; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_200 = PAR_io_pipe_phv_out_data_200; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_201 = PAR_io_pipe_phv_out_data_201; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_202 = PAR_io_pipe_phv_out_data_202; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_203 = PAR_io_pipe_phv_out_data_203; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_204 = PAR_io_pipe_phv_out_data_204; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_205 = PAR_io_pipe_phv_out_data_205; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_206 = PAR_io_pipe_phv_out_data_206; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_207 = PAR_io_pipe_phv_out_data_207; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_208 = PAR_io_pipe_phv_out_data_208; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_209 = PAR_io_pipe_phv_out_data_209; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_210 = PAR_io_pipe_phv_out_data_210; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_211 = PAR_io_pipe_phv_out_data_211; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_212 = PAR_io_pipe_phv_out_data_212; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_213 = PAR_io_pipe_phv_out_data_213; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_214 = PAR_io_pipe_phv_out_data_214; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_215 = PAR_io_pipe_phv_out_data_215; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_216 = PAR_io_pipe_phv_out_data_216; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_217 = PAR_io_pipe_phv_out_data_217; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_218 = PAR_io_pipe_phv_out_data_218; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_219 = PAR_io_pipe_phv_out_data_219; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_220 = PAR_io_pipe_phv_out_data_220; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_221 = PAR_io_pipe_phv_out_data_221; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_222 = PAR_io_pipe_phv_out_data_222; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_223 = PAR_io_pipe_phv_out_data_223; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_224 = PAR_io_pipe_phv_out_data_224; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_225 = PAR_io_pipe_phv_out_data_225; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_226 = PAR_io_pipe_phv_out_data_226; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_227 = PAR_io_pipe_phv_out_data_227; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_228 = PAR_io_pipe_phv_out_data_228; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_229 = PAR_io_pipe_phv_out_data_229; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_230 = PAR_io_pipe_phv_out_data_230; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_231 = PAR_io_pipe_phv_out_data_231; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_232 = PAR_io_pipe_phv_out_data_232; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_233 = PAR_io_pipe_phv_out_data_233; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_234 = PAR_io_pipe_phv_out_data_234; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_235 = PAR_io_pipe_phv_out_data_235; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_236 = PAR_io_pipe_phv_out_data_236; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_237 = PAR_io_pipe_phv_out_data_237; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_238 = PAR_io_pipe_phv_out_data_238; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_239 = PAR_io_pipe_phv_out_data_239; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_240 = PAR_io_pipe_phv_out_data_240; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_241 = PAR_io_pipe_phv_out_data_241; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_242 = PAR_io_pipe_phv_out_data_242; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_243 = PAR_io_pipe_phv_out_data_243; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_244 = PAR_io_pipe_phv_out_data_244; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_245 = PAR_io_pipe_phv_out_data_245; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_246 = PAR_io_pipe_phv_out_data_246; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_247 = PAR_io_pipe_phv_out_data_247; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_248 = PAR_io_pipe_phv_out_data_248; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_249 = PAR_io_pipe_phv_out_data_249; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_250 = PAR_io_pipe_phv_out_data_250; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_251 = PAR_io_pipe_phv_out_data_251; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_252 = PAR_io_pipe_phv_out_data_252; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_253 = PAR_io_pipe_phv_out_data_253; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_254 = PAR_io_pipe_phv_out_data_254; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_255 = PAR_io_pipe_phv_out_data_255; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_next_processor_id = PAR_io_pipe_phv_out_next_processor_id; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_next_config_id = PAR_io_pipe_phv_out_next_config_id; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_is_valid_processor = 1'h1; // @[pisa.scala 39:55]
  assign proc_0_io_mod_mat_mod_en = io_mod_proc_mod_0_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_config_id = io_mod_proc_mod_0_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_0_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_0_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_0_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_0_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_0_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_0_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_0_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_0_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_0_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_0_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_0_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_0_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_0_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_w_en = io_mod_proc_mod_0_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_0_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_w_addr = io_mod_proc_mod_0_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_w_data = io_mod_proc_mod_0_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_0_io_mod_exe_mod_en_0 = io_mod_proc_mod_0_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_0_io_mod_exe_mod_en_1 = io_mod_proc_mod_0_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_0_io_mod_exe_mod_addr = io_mod_proc_mod_0_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_0_io_mod_exe_mod_data_0 = io_mod_proc_mod_0_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_0_io_mod_exe_mod_data_1 = io_mod_proc_mod_0_exe_mod_data_1; // @[pisa.scala 29:20]
  assign proc_1_clock = clock;
  assign proc_1_io_pipe_phv_in_data_0 = proc_0_io_pipe_phv_out_data_0; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_1 = proc_0_io_pipe_phv_out_data_1; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_2 = proc_0_io_pipe_phv_out_data_2; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_3 = proc_0_io_pipe_phv_out_data_3; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_4 = proc_0_io_pipe_phv_out_data_4; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_5 = proc_0_io_pipe_phv_out_data_5; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_6 = proc_0_io_pipe_phv_out_data_6; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_7 = proc_0_io_pipe_phv_out_data_7; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_8 = proc_0_io_pipe_phv_out_data_8; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_9 = proc_0_io_pipe_phv_out_data_9; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_10 = proc_0_io_pipe_phv_out_data_10; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_11 = proc_0_io_pipe_phv_out_data_11; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_12 = proc_0_io_pipe_phv_out_data_12; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_13 = proc_0_io_pipe_phv_out_data_13; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_14 = proc_0_io_pipe_phv_out_data_14; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_15 = proc_0_io_pipe_phv_out_data_15; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_16 = proc_0_io_pipe_phv_out_data_16; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_17 = proc_0_io_pipe_phv_out_data_17; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_18 = proc_0_io_pipe_phv_out_data_18; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_19 = proc_0_io_pipe_phv_out_data_19; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_20 = proc_0_io_pipe_phv_out_data_20; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_21 = proc_0_io_pipe_phv_out_data_21; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_22 = proc_0_io_pipe_phv_out_data_22; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_23 = proc_0_io_pipe_phv_out_data_23; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_24 = proc_0_io_pipe_phv_out_data_24; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_25 = proc_0_io_pipe_phv_out_data_25; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_26 = proc_0_io_pipe_phv_out_data_26; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_27 = proc_0_io_pipe_phv_out_data_27; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_28 = proc_0_io_pipe_phv_out_data_28; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_29 = proc_0_io_pipe_phv_out_data_29; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_30 = proc_0_io_pipe_phv_out_data_30; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_31 = proc_0_io_pipe_phv_out_data_31; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_32 = proc_0_io_pipe_phv_out_data_32; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_33 = proc_0_io_pipe_phv_out_data_33; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_34 = proc_0_io_pipe_phv_out_data_34; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_35 = proc_0_io_pipe_phv_out_data_35; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_36 = proc_0_io_pipe_phv_out_data_36; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_37 = proc_0_io_pipe_phv_out_data_37; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_38 = proc_0_io_pipe_phv_out_data_38; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_39 = proc_0_io_pipe_phv_out_data_39; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_40 = proc_0_io_pipe_phv_out_data_40; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_41 = proc_0_io_pipe_phv_out_data_41; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_42 = proc_0_io_pipe_phv_out_data_42; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_43 = proc_0_io_pipe_phv_out_data_43; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_44 = proc_0_io_pipe_phv_out_data_44; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_45 = proc_0_io_pipe_phv_out_data_45; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_46 = proc_0_io_pipe_phv_out_data_46; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_47 = proc_0_io_pipe_phv_out_data_47; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_48 = proc_0_io_pipe_phv_out_data_48; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_49 = proc_0_io_pipe_phv_out_data_49; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_50 = proc_0_io_pipe_phv_out_data_50; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_51 = proc_0_io_pipe_phv_out_data_51; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_52 = proc_0_io_pipe_phv_out_data_52; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_53 = proc_0_io_pipe_phv_out_data_53; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_54 = proc_0_io_pipe_phv_out_data_54; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_55 = proc_0_io_pipe_phv_out_data_55; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_56 = proc_0_io_pipe_phv_out_data_56; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_57 = proc_0_io_pipe_phv_out_data_57; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_58 = proc_0_io_pipe_phv_out_data_58; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_59 = proc_0_io_pipe_phv_out_data_59; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_60 = proc_0_io_pipe_phv_out_data_60; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_61 = proc_0_io_pipe_phv_out_data_61; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_62 = proc_0_io_pipe_phv_out_data_62; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_63 = proc_0_io_pipe_phv_out_data_63; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_64 = proc_0_io_pipe_phv_out_data_64; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_65 = proc_0_io_pipe_phv_out_data_65; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_66 = proc_0_io_pipe_phv_out_data_66; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_67 = proc_0_io_pipe_phv_out_data_67; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_68 = proc_0_io_pipe_phv_out_data_68; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_69 = proc_0_io_pipe_phv_out_data_69; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_70 = proc_0_io_pipe_phv_out_data_70; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_71 = proc_0_io_pipe_phv_out_data_71; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_72 = proc_0_io_pipe_phv_out_data_72; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_73 = proc_0_io_pipe_phv_out_data_73; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_74 = proc_0_io_pipe_phv_out_data_74; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_75 = proc_0_io_pipe_phv_out_data_75; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_76 = proc_0_io_pipe_phv_out_data_76; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_77 = proc_0_io_pipe_phv_out_data_77; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_78 = proc_0_io_pipe_phv_out_data_78; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_79 = proc_0_io_pipe_phv_out_data_79; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_80 = proc_0_io_pipe_phv_out_data_80; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_81 = proc_0_io_pipe_phv_out_data_81; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_82 = proc_0_io_pipe_phv_out_data_82; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_83 = proc_0_io_pipe_phv_out_data_83; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_84 = proc_0_io_pipe_phv_out_data_84; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_85 = proc_0_io_pipe_phv_out_data_85; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_86 = proc_0_io_pipe_phv_out_data_86; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_87 = proc_0_io_pipe_phv_out_data_87; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_88 = proc_0_io_pipe_phv_out_data_88; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_89 = proc_0_io_pipe_phv_out_data_89; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_90 = proc_0_io_pipe_phv_out_data_90; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_91 = proc_0_io_pipe_phv_out_data_91; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_92 = proc_0_io_pipe_phv_out_data_92; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_93 = proc_0_io_pipe_phv_out_data_93; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_94 = proc_0_io_pipe_phv_out_data_94; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_95 = proc_0_io_pipe_phv_out_data_95; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_96 = proc_0_io_pipe_phv_out_data_96; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_97 = proc_0_io_pipe_phv_out_data_97; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_98 = proc_0_io_pipe_phv_out_data_98; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_99 = proc_0_io_pipe_phv_out_data_99; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_100 = proc_0_io_pipe_phv_out_data_100; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_101 = proc_0_io_pipe_phv_out_data_101; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_102 = proc_0_io_pipe_phv_out_data_102; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_103 = proc_0_io_pipe_phv_out_data_103; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_104 = proc_0_io_pipe_phv_out_data_104; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_105 = proc_0_io_pipe_phv_out_data_105; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_106 = proc_0_io_pipe_phv_out_data_106; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_107 = proc_0_io_pipe_phv_out_data_107; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_108 = proc_0_io_pipe_phv_out_data_108; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_109 = proc_0_io_pipe_phv_out_data_109; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_110 = proc_0_io_pipe_phv_out_data_110; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_111 = proc_0_io_pipe_phv_out_data_111; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_112 = proc_0_io_pipe_phv_out_data_112; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_113 = proc_0_io_pipe_phv_out_data_113; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_114 = proc_0_io_pipe_phv_out_data_114; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_115 = proc_0_io_pipe_phv_out_data_115; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_116 = proc_0_io_pipe_phv_out_data_116; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_117 = proc_0_io_pipe_phv_out_data_117; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_118 = proc_0_io_pipe_phv_out_data_118; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_119 = proc_0_io_pipe_phv_out_data_119; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_120 = proc_0_io_pipe_phv_out_data_120; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_121 = proc_0_io_pipe_phv_out_data_121; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_122 = proc_0_io_pipe_phv_out_data_122; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_123 = proc_0_io_pipe_phv_out_data_123; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_124 = proc_0_io_pipe_phv_out_data_124; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_125 = proc_0_io_pipe_phv_out_data_125; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_126 = proc_0_io_pipe_phv_out_data_126; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_127 = proc_0_io_pipe_phv_out_data_127; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_128 = proc_0_io_pipe_phv_out_data_128; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_129 = proc_0_io_pipe_phv_out_data_129; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_130 = proc_0_io_pipe_phv_out_data_130; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_131 = proc_0_io_pipe_phv_out_data_131; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_132 = proc_0_io_pipe_phv_out_data_132; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_133 = proc_0_io_pipe_phv_out_data_133; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_134 = proc_0_io_pipe_phv_out_data_134; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_135 = proc_0_io_pipe_phv_out_data_135; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_136 = proc_0_io_pipe_phv_out_data_136; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_137 = proc_0_io_pipe_phv_out_data_137; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_138 = proc_0_io_pipe_phv_out_data_138; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_139 = proc_0_io_pipe_phv_out_data_139; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_140 = proc_0_io_pipe_phv_out_data_140; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_141 = proc_0_io_pipe_phv_out_data_141; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_142 = proc_0_io_pipe_phv_out_data_142; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_143 = proc_0_io_pipe_phv_out_data_143; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_144 = proc_0_io_pipe_phv_out_data_144; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_145 = proc_0_io_pipe_phv_out_data_145; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_146 = proc_0_io_pipe_phv_out_data_146; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_147 = proc_0_io_pipe_phv_out_data_147; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_148 = proc_0_io_pipe_phv_out_data_148; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_149 = proc_0_io_pipe_phv_out_data_149; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_150 = proc_0_io_pipe_phv_out_data_150; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_151 = proc_0_io_pipe_phv_out_data_151; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_152 = proc_0_io_pipe_phv_out_data_152; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_153 = proc_0_io_pipe_phv_out_data_153; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_154 = proc_0_io_pipe_phv_out_data_154; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_155 = proc_0_io_pipe_phv_out_data_155; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_156 = proc_0_io_pipe_phv_out_data_156; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_157 = proc_0_io_pipe_phv_out_data_157; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_158 = proc_0_io_pipe_phv_out_data_158; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_159 = proc_0_io_pipe_phv_out_data_159; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_160 = proc_0_io_pipe_phv_out_data_160; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_161 = proc_0_io_pipe_phv_out_data_161; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_162 = proc_0_io_pipe_phv_out_data_162; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_163 = proc_0_io_pipe_phv_out_data_163; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_164 = proc_0_io_pipe_phv_out_data_164; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_165 = proc_0_io_pipe_phv_out_data_165; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_166 = proc_0_io_pipe_phv_out_data_166; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_167 = proc_0_io_pipe_phv_out_data_167; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_168 = proc_0_io_pipe_phv_out_data_168; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_169 = proc_0_io_pipe_phv_out_data_169; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_170 = proc_0_io_pipe_phv_out_data_170; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_171 = proc_0_io_pipe_phv_out_data_171; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_172 = proc_0_io_pipe_phv_out_data_172; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_173 = proc_0_io_pipe_phv_out_data_173; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_174 = proc_0_io_pipe_phv_out_data_174; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_175 = proc_0_io_pipe_phv_out_data_175; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_176 = proc_0_io_pipe_phv_out_data_176; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_177 = proc_0_io_pipe_phv_out_data_177; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_178 = proc_0_io_pipe_phv_out_data_178; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_179 = proc_0_io_pipe_phv_out_data_179; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_180 = proc_0_io_pipe_phv_out_data_180; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_181 = proc_0_io_pipe_phv_out_data_181; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_182 = proc_0_io_pipe_phv_out_data_182; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_183 = proc_0_io_pipe_phv_out_data_183; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_184 = proc_0_io_pipe_phv_out_data_184; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_185 = proc_0_io_pipe_phv_out_data_185; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_186 = proc_0_io_pipe_phv_out_data_186; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_187 = proc_0_io_pipe_phv_out_data_187; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_188 = proc_0_io_pipe_phv_out_data_188; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_189 = proc_0_io_pipe_phv_out_data_189; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_190 = proc_0_io_pipe_phv_out_data_190; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_191 = proc_0_io_pipe_phv_out_data_191; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_192 = proc_0_io_pipe_phv_out_data_192; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_193 = proc_0_io_pipe_phv_out_data_193; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_194 = proc_0_io_pipe_phv_out_data_194; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_195 = proc_0_io_pipe_phv_out_data_195; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_196 = proc_0_io_pipe_phv_out_data_196; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_197 = proc_0_io_pipe_phv_out_data_197; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_198 = proc_0_io_pipe_phv_out_data_198; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_199 = proc_0_io_pipe_phv_out_data_199; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_200 = proc_0_io_pipe_phv_out_data_200; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_201 = proc_0_io_pipe_phv_out_data_201; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_202 = proc_0_io_pipe_phv_out_data_202; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_203 = proc_0_io_pipe_phv_out_data_203; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_204 = proc_0_io_pipe_phv_out_data_204; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_205 = proc_0_io_pipe_phv_out_data_205; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_206 = proc_0_io_pipe_phv_out_data_206; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_207 = proc_0_io_pipe_phv_out_data_207; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_208 = proc_0_io_pipe_phv_out_data_208; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_209 = proc_0_io_pipe_phv_out_data_209; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_210 = proc_0_io_pipe_phv_out_data_210; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_211 = proc_0_io_pipe_phv_out_data_211; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_212 = proc_0_io_pipe_phv_out_data_212; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_213 = proc_0_io_pipe_phv_out_data_213; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_214 = proc_0_io_pipe_phv_out_data_214; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_215 = proc_0_io_pipe_phv_out_data_215; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_216 = proc_0_io_pipe_phv_out_data_216; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_217 = proc_0_io_pipe_phv_out_data_217; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_218 = proc_0_io_pipe_phv_out_data_218; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_219 = proc_0_io_pipe_phv_out_data_219; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_220 = proc_0_io_pipe_phv_out_data_220; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_221 = proc_0_io_pipe_phv_out_data_221; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_222 = proc_0_io_pipe_phv_out_data_222; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_223 = proc_0_io_pipe_phv_out_data_223; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_224 = proc_0_io_pipe_phv_out_data_224; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_225 = proc_0_io_pipe_phv_out_data_225; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_226 = proc_0_io_pipe_phv_out_data_226; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_227 = proc_0_io_pipe_phv_out_data_227; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_228 = proc_0_io_pipe_phv_out_data_228; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_229 = proc_0_io_pipe_phv_out_data_229; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_230 = proc_0_io_pipe_phv_out_data_230; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_231 = proc_0_io_pipe_phv_out_data_231; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_232 = proc_0_io_pipe_phv_out_data_232; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_233 = proc_0_io_pipe_phv_out_data_233; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_234 = proc_0_io_pipe_phv_out_data_234; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_235 = proc_0_io_pipe_phv_out_data_235; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_236 = proc_0_io_pipe_phv_out_data_236; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_237 = proc_0_io_pipe_phv_out_data_237; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_238 = proc_0_io_pipe_phv_out_data_238; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_239 = proc_0_io_pipe_phv_out_data_239; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_240 = proc_0_io_pipe_phv_out_data_240; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_241 = proc_0_io_pipe_phv_out_data_241; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_242 = proc_0_io_pipe_phv_out_data_242; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_243 = proc_0_io_pipe_phv_out_data_243; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_244 = proc_0_io_pipe_phv_out_data_244; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_245 = proc_0_io_pipe_phv_out_data_245; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_246 = proc_0_io_pipe_phv_out_data_246; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_247 = proc_0_io_pipe_phv_out_data_247; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_248 = proc_0_io_pipe_phv_out_data_248; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_249 = proc_0_io_pipe_phv_out_data_249; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_250 = proc_0_io_pipe_phv_out_data_250; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_251 = proc_0_io_pipe_phv_out_data_251; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_252 = proc_0_io_pipe_phv_out_data_252; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_253 = proc_0_io_pipe_phv_out_data_253; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_254 = proc_0_io_pipe_phv_out_data_254; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_255 = proc_0_io_pipe_phv_out_data_255; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_next_processor_id = proc_0_io_pipe_phv_out_next_processor_id; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_next_config_id = proc_0_io_pipe_phv_out_next_config_id; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_is_valid_processor = 4'h1 == proc_0_io_pipe_phv_out_next_processor_id; // @[pisa.scala 36:62]
  assign proc_1_io_mod_mat_mod_en = io_mod_proc_mod_1_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_config_id = io_mod_proc_mod_1_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_1_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_1_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_1_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_1_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_1_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_1_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_1_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_1_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_1_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_1_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_1_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_1_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_1_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_w_en = io_mod_proc_mod_1_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_1_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_w_addr = io_mod_proc_mod_1_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_w_data = io_mod_proc_mod_1_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_1_io_mod_exe_mod_en_0 = io_mod_proc_mod_1_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_1_io_mod_exe_mod_en_1 = io_mod_proc_mod_1_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_1_io_mod_exe_mod_addr = io_mod_proc_mod_1_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_1_io_mod_exe_mod_data_0 = io_mod_proc_mod_1_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_1_io_mod_exe_mod_data_1 = io_mod_proc_mod_1_exe_mod_data_1; // @[pisa.scala 29:20]
  assign proc_2_clock = clock;
  assign proc_2_io_pipe_phv_in_data_0 = proc_1_io_pipe_phv_out_data_0; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_1 = proc_1_io_pipe_phv_out_data_1; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_2 = proc_1_io_pipe_phv_out_data_2; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_3 = proc_1_io_pipe_phv_out_data_3; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_4 = proc_1_io_pipe_phv_out_data_4; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_5 = proc_1_io_pipe_phv_out_data_5; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_6 = proc_1_io_pipe_phv_out_data_6; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_7 = proc_1_io_pipe_phv_out_data_7; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_8 = proc_1_io_pipe_phv_out_data_8; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_9 = proc_1_io_pipe_phv_out_data_9; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_10 = proc_1_io_pipe_phv_out_data_10; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_11 = proc_1_io_pipe_phv_out_data_11; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_12 = proc_1_io_pipe_phv_out_data_12; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_13 = proc_1_io_pipe_phv_out_data_13; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_14 = proc_1_io_pipe_phv_out_data_14; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_15 = proc_1_io_pipe_phv_out_data_15; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_16 = proc_1_io_pipe_phv_out_data_16; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_17 = proc_1_io_pipe_phv_out_data_17; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_18 = proc_1_io_pipe_phv_out_data_18; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_19 = proc_1_io_pipe_phv_out_data_19; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_20 = proc_1_io_pipe_phv_out_data_20; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_21 = proc_1_io_pipe_phv_out_data_21; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_22 = proc_1_io_pipe_phv_out_data_22; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_23 = proc_1_io_pipe_phv_out_data_23; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_24 = proc_1_io_pipe_phv_out_data_24; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_25 = proc_1_io_pipe_phv_out_data_25; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_26 = proc_1_io_pipe_phv_out_data_26; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_27 = proc_1_io_pipe_phv_out_data_27; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_28 = proc_1_io_pipe_phv_out_data_28; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_29 = proc_1_io_pipe_phv_out_data_29; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_30 = proc_1_io_pipe_phv_out_data_30; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_31 = proc_1_io_pipe_phv_out_data_31; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_32 = proc_1_io_pipe_phv_out_data_32; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_33 = proc_1_io_pipe_phv_out_data_33; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_34 = proc_1_io_pipe_phv_out_data_34; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_35 = proc_1_io_pipe_phv_out_data_35; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_36 = proc_1_io_pipe_phv_out_data_36; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_37 = proc_1_io_pipe_phv_out_data_37; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_38 = proc_1_io_pipe_phv_out_data_38; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_39 = proc_1_io_pipe_phv_out_data_39; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_40 = proc_1_io_pipe_phv_out_data_40; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_41 = proc_1_io_pipe_phv_out_data_41; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_42 = proc_1_io_pipe_phv_out_data_42; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_43 = proc_1_io_pipe_phv_out_data_43; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_44 = proc_1_io_pipe_phv_out_data_44; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_45 = proc_1_io_pipe_phv_out_data_45; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_46 = proc_1_io_pipe_phv_out_data_46; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_47 = proc_1_io_pipe_phv_out_data_47; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_48 = proc_1_io_pipe_phv_out_data_48; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_49 = proc_1_io_pipe_phv_out_data_49; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_50 = proc_1_io_pipe_phv_out_data_50; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_51 = proc_1_io_pipe_phv_out_data_51; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_52 = proc_1_io_pipe_phv_out_data_52; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_53 = proc_1_io_pipe_phv_out_data_53; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_54 = proc_1_io_pipe_phv_out_data_54; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_55 = proc_1_io_pipe_phv_out_data_55; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_56 = proc_1_io_pipe_phv_out_data_56; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_57 = proc_1_io_pipe_phv_out_data_57; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_58 = proc_1_io_pipe_phv_out_data_58; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_59 = proc_1_io_pipe_phv_out_data_59; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_60 = proc_1_io_pipe_phv_out_data_60; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_61 = proc_1_io_pipe_phv_out_data_61; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_62 = proc_1_io_pipe_phv_out_data_62; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_63 = proc_1_io_pipe_phv_out_data_63; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_64 = proc_1_io_pipe_phv_out_data_64; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_65 = proc_1_io_pipe_phv_out_data_65; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_66 = proc_1_io_pipe_phv_out_data_66; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_67 = proc_1_io_pipe_phv_out_data_67; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_68 = proc_1_io_pipe_phv_out_data_68; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_69 = proc_1_io_pipe_phv_out_data_69; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_70 = proc_1_io_pipe_phv_out_data_70; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_71 = proc_1_io_pipe_phv_out_data_71; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_72 = proc_1_io_pipe_phv_out_data_72; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_73 = proc_1_io_pipe_phv_out_data_73; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_74 = proc_1_io_pipe_phv_out_data_74; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_75 = proc_1_io_pipe_phv_out_data_75; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_76 = proc_1_io_pipe_phv_out_data_76; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_77 = proc_1_io_pipe_phv_out_data_77; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_78 = proc_1_io_pipe_phv_out_data_78; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_79 = proc_1_io_pipe_phv_out_data_79; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_80 = proc_1_io_pipe_phv_out_data_80; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_81 = proc_1_io_pipe_phv_out_data_81; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_82 = proc_1_io_pipe_phv_out_data_82; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_83 = proc_1_io_pipe_phv_out_data_83; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_84 = proc_1_io_pipe_phv_out_data_84; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_85 = proc_1_io_pipe_phv_out_data_85; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_86 = proc_1_io_pipe_phv_out_data_86; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_87 = proc_1_io_pipe_phv_out_data_87; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_88 = proc_1_io_pipe_phv_out_data_88; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_89 = proc_1_io_pipe_phv_out_data_89; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_90 = proc_1_io_pipe_phv_out_data_90; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_91 = proc_1_io_pipe_phv_out_data_91; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_92 = proc_1_io_pipe_phv_out_data_92; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_93 = proc_1_io_pipe_phv_out_data_93; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_94 = proc_1_io_pipe_phv_out_data_94; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_95 = proc_1_io_pipe_phv_out_data_95; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_96 = proc_1_io_pipe_phv_out_data_96; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_97 = proc_1_io_pipe_phv_out_data_97; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_98 = proc_1_io_pipe_phv_out_data_98; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_99 = proc_1_io_pipe_phv_out_data_99; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_100 = proc_1_io_pipe_phv_out_data_100; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_101 = proc_1_io_pipe_phv_out_data_101; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_102 = proc_1_io_pipe_phv_out_data_102; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_103 = proc_1_io_pipe_phv_out_data_103; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_104 = proc_1_io_pipe_phv_out_data_104; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_105 = proc_1_io_pipe_phv_out_data_105; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_106 = proc_1_io_pipe_phv_out_data_106; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_107 = proc_1_io_pipe_phv_out_data_107; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_108 = proc_1_io_pipe_phv_out_data_108; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_109 = proc_1_io_pipe_phv_out_data_109; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_110 = proc_1_io_pipe_phv_out_data_110; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_111 = proc_1_io_pipe_phv_out_data_111; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_112 = proc_1_io_pipe_phv_out_data_112; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_113 = proc_1_io_pipe_phv_out_data_113; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_114 = proc_1_io_pipe_phv_out_data_114; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_115 = proc_1_io_pipe_phv_out_data_115; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_116 = proc_1_io_pipe_phv_out_data_116; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_117 = proc_1_io_pipe_phv_out_data_117; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_118 = proc_1_io_pipe_phv_out_data_118; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_119 = proc_1_io_pipe_phv_out_data_119; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_120 = proc_1_io_pipe_phv_out_data_120; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_121 = proc_1_io_pipe_phv_out_data_121; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_122 = proc_1_io_pipe_phv_out_data_122; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_123 = proc_1_io_pipe_phv_out_data_123; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_124 = proc_1_io_pipe_phv_out_data_124; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_125 = proc_1_io_pipe_phv_out_data_125; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_126 = proc_1_io_pipe_phv_out_data_126; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_127 = proc_1_io_pipe_phv_out_data_127; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_128 = proc_1_io_pipe_phv_out_data_128; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_129 = proc_1_io_pipe_phv_out_data_129; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_130 = proc_1_io_pipe_phv_out_data_130; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_131 = proc_1_io_pipe_phv_out_data_131; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_132 = proc_1_io_pipe_phv_out_data_132; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_133 = proc_1_io_pipe_phv_out_data_133; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_134 = proc_1_io_pipe_phv_out_data_134; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_135 = proc_1_io_pipe_phv_out_data_135; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_136 = proc_1_io_pipe_phv_out_data_136; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_137 = proc_1_io_pipe_phv_out_data_137; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_138 = proc_1_io_pipe_phv_out_data_138; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_139 = proc_1_io_pipe_phv_out_data_139; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_140 = proc_1_io_pipe_phv_out_data_140; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_141 = proc_1_io_pipe_phv_out_data_141; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_142 = proc_1_io_pipe_phv_out_data_142; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_143 = proc_1_io_pipe_phv_out_data_143; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_144 = proc_1_io_pipe_phv_out_data_144; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_145 = proc_1_io_pipe_phv_out_data_145; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_146 = proc_1_io_pipe_phv_out_data_146; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_147 = proc_1_io_pipe_phv_out_data_147; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_148 = proc_1_io_pipe_phv_out_data_148; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_149 = proc_1_io_pipe_phv_out_data_149; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_150 = proc_1_io_pipe_phv_out_data_150; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_151 = proc_1_io_pipe_phv_out_data_151; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_152 = proc_1_io_pipe_phv_out_data_152; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_153 = proc_1_io_pipe_phv_out_data_153; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_154 = proc_1_io_pipe_phv_out_data_154; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_155 = proc_1_io_pipe_phv_out_data_155; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_156 = proc_1_io_pipe_phv_out_data_156; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_157 = proc_1_io_pipe_phv_out_data_157; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_158 = proc_1_io_pipe_phv_out_data_158; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_159 = proc_1_io_pipe_phv_out_data_159; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_160 = proc_1_io_pipe_phv_out_data_160; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_161 = proc_1_io_pipe_phv_out_data_161; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_162 = proc_1_io_pipe_phv_out_data_162; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_163 = proc_1_io_pipe_phv_out_data_163; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_164 = proc_1_io_pipe_phv_out_data_164; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_165 = proc_1_io_pipe_phv_out_data_165; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_166 = proc_1_io_pipe_phv_out_data_166; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_167 = proc_1_io_pipe_phv_out_data_167; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_168 = proc_1_io_pipe_phv_out_data_168; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_169 = proc_1_io_pipe_phv_out_data_169; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_170 = proc_1_io_pipe_phv_out_data_170; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_171 = proc_1_io_pipe_phv_out_data_171; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_172 = proc_1_io_pipe_phv_out_data_172; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_173 = proc_1_io_pipe_phv_out_data_173; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_174 = proc_1_io_pipe_phv_out_data_174; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_175 = proc_1_io_pipe_phv_out_data_175; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_176 = proc_1_io_pipe_phv_out_data_176; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_177 = proc_1_io_pipe_phv_out_data_177; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_178 = proc_1_io_pipe_phv_out_data_178; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_179 = proc_1_io_pipe_phv_out_data_179; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_180 = proc_1_io_pipe_phv_out_data_180; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_181 = proc_1_io_pipe_phv_out_data_181; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_182 = proc_1_io_pipe_phv_out_data_182; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_183 = proc_1_io_pipe_phv_out_data_183; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_184 = proc_1_io_pipe_phv_out_data_184; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_185 = proc_1_io_pipe_phv_out_data_185; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_186 = proc_1_io_pipe_phv_out_data_186; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_187 = proc_1_io_pipe_phv_out_data_187; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_188 = proc_1_io_pipe_phv_out_data_188; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_189 = proc_1_io_pipe_phv_out_data_189; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_190 = proc_1_io_pipe_phv_out_data_190; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_191 = proc_1_io_pipe_phv_out_data_191; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_192 = proc_1_io_pipe_phv_out_data_192; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_193 = proc_1_io_pipe_phv_out_data_193; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_194 = proc_1_io_pipe_phv_out_data_194; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_195 = proc_1_io_pipe_phv_out_data_195; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_196 = proc_1_io_pipe_phv_out_data_196; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_197 = proc_1_io_pipe_phv_out_data_197; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_198 = proc_1_io_pipe_phv_out_data_198; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_199 = proc_1_io_pipe_phv_out_data_199; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_200 = proc_1_io_pipe_phv_out_data_200; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_201 = proc_1_io_pipe_phv_out_data_201; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_202 = proc_1_io_pipe_phv_out_data_202; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_203 = proc_1_io_pipe_phv_out_data_203; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_204 = proc_1_io_pipe_phv_out_data_204; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_205 = proc_1_io_pipe_phv_out_data_205; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_206 = proc_1_io_pipe_phv_out_data_206; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_207 = proc_1_io_pipe_phv_out_data_207; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_208 = proc_1_io_pipe_phv_out_data_208; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_209 = proc_1_io_pipe_phv_out_data_209; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_210 = proc_1_io_pipe_phv_out_data_210; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_211 = proc_1_io_pipe_phv_out_data_211; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_212 = proc_1_io_pipe_phv_out_data_212; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_213 = proc_1_io_pipe_phv_out_data_213; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_214 = proc_1_io_pipe_phv_out_data_214; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_215 = proc_1_io_pipe_phv_out_data_215; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_216 = proc_1_io_pipe_phv_out_data_216; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_217 = proc_1_io_pipe_phv_out_data_217; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_218 = proc_1_io_pipe_phv_out_data_218; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_219 = proc_1_io_pipe_phv_out_data_219; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_220 = proc_1_io_pipe_phv_out_data_220; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_221 = proc_1_io_pipe_phv_out_data_221; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_222 = proc_1_io_pipe_phv_out_data_222; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_223 = proc_1_io_pipe_phv_out_data_223; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_224 = proc_1_io_pipe_phv_out_data_224; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_225 = proc_1_io_pipe_phv_out_data_225; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_226 = proc_1_io_pipe_phv_out_data_226; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_227 = proc_1_io_pipe_phv_out_data_227; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_228 = proc_1_io_pipe_phv_out_data_228; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_229 = proc_1_io_pipe_phv_out_data_229; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_230 = proc_1_io_pipe_phv_out_data_230; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_231 = proc_1_io_pipe_phv_out_data_231; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_232 = proc_1_io_pipe_phv_out_data_232; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_233 = proc_1_io_pipe_phv_out_data_233; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_234 = proc_1_io_pipe_phv_out_data_234; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_235 = proc_1_io_pipe_phv_out_data_235; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_236 = proc_1_io_pipe_phv_out_data_236; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_237 = proc_1_io_pipe_phv_out_data_237; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_238 = proc_1_io_pipe_phv_out_data_238; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_239 = proc_1_io_pipe_phv_out_data_239; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_240 = proc_1_io_pipe_phv_out_data_240; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_241 = proc_1_io_pipe_phv_out_data_241; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_242 = proc_1_io_pipe_phv_out_data_242; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_243 = proc_1_io_pipe_phv_out_data_243; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_244 = proc_1_io_pipe_phv_out_data_244; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_245 = proc_1_io_pipe_phv_out_data_245; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_246 = proc_1_io_pipe_phv_out_data_246; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_247 = proc_1_io_pipe_phv_out_data_247; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_248 = proc_1_io_pipe_phv_out_data_248; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_249 = proc_1_io_pipe_phv_out_data_249; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_250 = proc_1_io_pipe_phv_out_data_250; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_251 = proc_1_io_pipe_phv_out_data_251; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_252 = proc_1_io_pipe_phv_out_data_252; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_253 = proc_1_io_pipe_phv_out_data_253; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_254 = proc_1_io_pipe_phv_out_data_254; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_255 = proc_1_io_pipe_phv_out_data_255; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_next_processor_id = proc_1_io_pipe_phv_out_next_processor_id; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_next_config_id = proc_1_io_pipe_phv_out_next_config_id; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_is_valid_processor = 4'h2 == proc_1_io_pipe_phv_out_next_processor_id; // @[pisa.scala 36:62]
  assign proc_2_io_mod_mat_mod_en = io_mod_proc_mod_2_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_config_id = io_mod_proc_mod_2_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_2_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_2_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_2_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_2_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_2_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_2_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_2_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_2_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_2_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_2_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_2_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_2_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_2_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_w_en = io_mod_proc_mod_2_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_2_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_w_addr = io_mod_proc_mod_2_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_w_data = io_mod_proc_mod_2_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_2_io_mod_exe_mod_en_0 = io_mod_proc_mod_2_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_2_io_mod_exe_mod_en_1 = io_mod_proc_mod_2_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_2_io_mod_exe_mod_addr = io_mod_proc_mod_2_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_2_io_mod_exe_mod_data_0 = io_mod_proc_mod_2_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_2_io_mod_exe_mod_data_1 = io_mod_proc_mod_2_exe_mod_data_1; // @[pisa.scala 29:20]
  assign proc_3_clock = clock;
  assign proc_3_io_pipe_phv_in_data_0 = proc_2_io_pipe_phv_out_data_0; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_1 = proc_2_io_pipe_phv_out_data_1; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_2 = proc_2_io_pipe_phv_out_data_2; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_3 = proc_2_io_pipe_phv_out_data_3; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_4 = proc_2_io_pipe_phv_out_data_4; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_5 = proc_2_io_pipe_phv_out_data_5; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_6 = proc_2_io_pipe_phv_out_data_6; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_7 = proc_2_io_pipe_phv_out_data_7; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_8 = proc_2_io_pipe_phv_out_data_8; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_9 = proc_2_io_pipe_phv_out_data_9; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_10 = proc_2_io_pipe_phv_out_data_10; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_11 = proc_2_io_pipe_phv_out_data_11; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_12 = proc_2_io_pipe_phv_out_data_12; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_13 = proc_2_io_pipe_phv_out_data_13; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_14 = proc_2_io_pipe_phv_out_data_14; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_15 = proc_2_io_pipe_phv_out_data_15; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_16 = proc_2_io_pipe_phv_out_data_16; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_17 = proc_2_io_pipe_phv_out_data_17; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_18 = proc_2_io_pipe_phv_out_data_18; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_19 = proc_2_io_pipe_phv_out_data_19; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_20 = proc_2_io_pipe_phv_out_data_20; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_21 = proc_2_io_pipe_phv_out_data_21; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_22 = proc_2_io_pipe_phv_out_data_22; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_23 = proc_2_io_pipe_phv_out_data_23; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_24 = proc_2_io_pipe_phv_out_data_24; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_25 = proc_2_io_pipe_phv_out_data_25; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_26 = proc_2_io_pipe_phv_out_data_26; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_27 = proc_2_io_pipe_phv_out_data_27; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_28 = proc_2_io_pipe_phv_out_data_28; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_29 = proc_2_io_pipe_phv_out_data_29; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_30 = proc_2_io_pipe_phv_out_data_30; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_31 = proc_2_io_pipe_phv_out_data_31; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_32 = proc_2_io_pipe_phv_out_data_32; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_33 = proc_2_io_pipe_phv_out_data_33; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_34 = proc_2_io_pipe_phv_out_data_34; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_35 = proc_2_io_pipe_phv_out_data_35; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_36 = proc_2_io_pipe_phv_out_data_36; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_37 = proc_2_io_pipe_phv_out_data_37; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_38 = proc_2_io_pipe_phv_out_data_38; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_39 = proc_2_io_pipe_phv_out_data_39; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_40 = proc_2_io_pipe_phv_out_data_40; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_41 = proc_2_io_pipe_phv_out_data_41; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_42 = proc_2_io_pipe_phv_out_data_42; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_43 = proc_2_io_pipe_phv_out_data_43; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_44 = proc_2_io_pipe_phv_out_data_44; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_45 = proc_2_io_pipe_phv_out_data_45; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_46 = proc_2_io_pipe_phv_out_data_46; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_47 = proc_2_io_pipe_phv_out_data_47; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_48 = proc_2_io_pipe_phv_out_data_48; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_49 = proc_2_io_pipe_phv_out_data_49; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_50 = proc_2_io_pipe_phv_out_data_50; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_51 = proc_2_io_pipe_phv_out_data_51; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_52 = proc_2_io_pipe_phv_out_data_52; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_53 = proc_2_io_pipe_phv_out_data_53; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_54 = proc_2_io_pipe_phv_out_data_54; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_55 = proc_2_io_pipe_phv_out_data_55; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_56 = proc_2_io_pipe_phv_out_data_56; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_57 = proc_2_io_pipe_phv_out_data_57; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_58 = proc_2_io_pipe_phv_out_data_58; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_59 = proc_2_io_pipe_phv_out_data_59; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_60 = proc_2_io_pipe_phv_out_data_60; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_61 = proc_2_io_pipe_phv_out_data_61; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_62 = proc_2_io_pipe_phv_out_data_62; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_63 = proc_2_io_pipe_phv_out_data_63; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_64 = proc_2_io_pipe_phv_out_data_64; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_65 = proc_2_io_pipe_phv_out_data_65; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_66 = proc_2_io_pipe_phv_out_data_66; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_67 = proc_2_io_pipe_phv_out_data_67; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_68 = proc_2_io_pipe_phv_out_data_68; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_69 = proc_2_io_pipe_phv_out_data_69; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_70 = proc_2_io_pipe_phv_out_data_70; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_71 = proc_2_io_pipe_phv_out_data_71; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_72 = proc_2_io_pipe_phv_out_data_72; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_73 = proc_2_io_pipe_phv_out_data_73; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_74 = proc_2_io_pipe_phv_out_data_74; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_75 = proc_2_io_pipe_phv_out_data_75; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_76 = proc_2_io_pipe_phv_out_data_76; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_77 = proc_2_io_pipe_phv_out_data_77; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_78 = proc_2_io_pipe_phv_out_data_78; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_79 = proc_2_io_pipe_phv_out_data_79; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_80 = proc_2_io_pipe_phv_out_data_80; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_81 = proc_2_io_pipe_phv_out_data_81; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_82 = proc_2_io_pipe_phv_out_data_82; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_83 = proc_2_io_pipe_phv_out_data_83; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_84 = proc_2_io_pipe_phv_out_data_84; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_85 = proc_2_io_pipe_phv_out_data_85; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_86 = proc_2_io_pipe_phv_out_data_86; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_87 = proc_2_io_pipe_phv_out_data_87; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_88 = proc_2_io_pipe_phv_out_data_88; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_89 = proc_2_io_pipe_phv_out_data_89; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_90 = proc_2_io_pipe_phv_out_data_90; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_91 = proc_2_io_pipe_phv_out_data_91; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_92 = proc_2_io_pipe_phv_out_data_92; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_93 = proc_2_io_pipe_phv_out_data_93; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_94 = proc_2_io_pipe_phv_out_data_94; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_95 = proc_2_io_pipe_phv_out_data_95; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_96 = proc_2_io_pipe_phv_out_data_96; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_97 = proc_2_io_pipe_phv_out_data_97; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_98 = proc_2_io_pipe_phv_out_data_98; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_99 = proc_2_io_pipe_phv_out_data_99; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_100 = proc_2_io_pipe_phv_out_data_100; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_101 = proc_2_io_pipe_phv_out_data_101; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_102 = proc_2_io_pipe_phv_out_data_102; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_103 = proc_2_io_pipe_phv_out_data_103; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_104 = proc_2_io_pipe_phv_out_data_104; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_105 = proc_2_io_pipe_phv_out_data_105; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_106 = proc_2_io_pipe_phv_out_data_106; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_107 = proc_2_io_pipe_phv_out_data_107; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_108 = proc_2_io_pipe_phv_out_data_108; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_109 = proc_2_io_pipe_phv_out_data_109; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_110 = proc_2_io_pipe_phv_out_data_110; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_111 = proc_2_io_pipe_phv_out_data_111; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_112 = proc_2_io_pipe_phv_out_data_112; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_113 = proc_2_io_pipe_phv_out_data_113; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_114 = proc_2_io_pipe_phv_out_data_114; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_115 = proc_2_io_pipe_phv_out_data_115; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_116 = proc_2_io_pipe_phv_out_data_116; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_117 = proc_2_io_pipe_phv_out_data_117; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_118 = proc_2_io_pipe_phv_out_data_118; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_119 = proc_2_io_pipe_phv_out_data_119; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_120 = proc_2_io_pipe_phv_out_data_120; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_121 = proc_2_io_pipe_phv_out_data_121; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_122 = proc_2_io_pipe_phv_out_data_122; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_123 = proc_2_io_pipe_phv_out_data_123; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_124 = proc_2_io_pipe_phv_out_data_124; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_125 = proc_2_io_pipe_phv_out_data_125; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_126 = proc_2_io_pipe_phv_out_data_126; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_127 = proc_2_io_pipe_phv_out_data_127; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_128 = proc_2_io_pipe_phv_out_data_128; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_129 = proc_2_io_pipe_phv_out_data_129; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_130 = proc_2_io_pipe_phv_out_data_130; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_131 = proc_2_io_pipe_phv_out_data_131; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_132 = proc_2_io_pipe_phv_out_data_132; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_133 = proc_2_io_pipe_phv_out_data_133; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_134 = proc_2_io_pipe_phv_out_data_134; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_135 = proc_2_io_pipe_phv_out_data_135; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_136 = proc_2_io_pipe_phv_out_data_136; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_137 = proc_2_io_pipe_phv_out_data_137; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_138 = proc_2_io_pipe_phv_out_data_138; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_139 = proc_2_io_pipe_phv_out_data_139; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_140 = proc_2_io_pipe_phv_out_data_140; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_141 = proc_2_io_pipe_phv_out_data_141; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_142 = proc_2_io_pipe_phv_out_data_142; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_143 = proc_2_io_pipe_phv_out_data_143; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_144 = proc_2_io_pipe_phv_out_data_144; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_145 = proc_2_io_pipe_phv_out_data_145; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_146 = proc_2_io_pipe_phv_out_data_146; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_147 = proc_2_io_pipe_phv_out_data_147; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_148 = proc_2_io_pipe_phv_out_data_148; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_149 = proc_2_io_pipe_phv_out_data_149; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_150 = proc_2_io_pipe_phv_out_data_150; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_151 = proc_2_io_pipe_phv_out_data_151; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_152 = proc_2_io_pipe_phv_out_data_152; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_153 = proc_2_io_pipe_phv_out_data_153; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_154 = proc_2_io_pipe_phv_out_data_154; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_155 = proc_2_io_pipe_phv_out_data_155; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_156 = proc_2_io_pipe_phv_out_data_156; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_157 = proc_2_io_pipe_phv_out_data_157; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_158 = proc_2_io_pipe_phv_out_data_158; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_159 = proc_2_io_pipe_phv_out_data_159; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_160 = proc_2_io_pipe_phv_out_data_160; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_161 = proc_2_io_pipe_phv_out_data_161; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_162 = proc_2_io_pipe_phv_out_data_162; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_163 = proc_2_io_pipe_phv_out_data_163; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_164 = proc_2_io_pipe_phv_out_data_164; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_165 = proc_2_io_pipe_phv_out_data_165; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_166 = proc_2_io_pipe_phv_out_data_166; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_167 = proc_2_io_pipe_phv_out_data_167; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_168 = proc_2_io_pipe_phv_out_data_168; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_169 = proc_2_io_pipe_phv_out_data_169; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_170 = proc_2_io_pipe_phv_out_data_170; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_171 = proc_2_io_pipe_phv_out_data_171; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_172 = proc_2_io_pipe_phv_out_data_172; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_173 = proc_2_io_pipe_phv_out_data_173; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_174 = proc_2_io_pipe_phv_out_data_174; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_175 = proc_2_io_pipe_phv_out_data_175; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_176 = proc_2_io_pipe_phv_out_data_176; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_177 = proc_2_io_pipe_phv_out_data_177; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_178 = proc_2_io_pipe_phv_out_data_178; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_179 = proc_2_io_pipe_phv_out_data_179; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_180 = proc_2_io_pipe_phv_out_data_180; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_181 = proc_2_io_pipe_phv_out_data_181; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_182 = proc_2_io_pipe_phv_out_data_182; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_183 = proc_2_io_pipe_phv_out_data_183; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_184 = proc_2_io_pipe_phv_out_data_184; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_185 = proc_2_io_pipe_phv_out_data_185; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_186 = proc_2_io_pipe_phv_out_data_186; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_187 = proc_2_io_pipe_phv_out_data_187; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_188 = proc_2_io_pipe_phv_out_data_188; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_189 = proc_2_io_pipe_phv_out_data_189; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_190 = proc_2_io_pipe_phv_out_data_190; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_191 = proc_2_io_pipe_phv_out_data_191; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_192 = proc_2_io_pipe_phv_out_data_192; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_193 = proc_2_io_pipe_phv_out_data_193; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_194 = proc_2_io_pipe_phv_out_data_194; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_195 = proc_2_io_pipe_phv_out_data_195; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_196 = proc_2_io_pipe_phv_out_data_196; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_197 = proc_2_io_pipe_phv_out_data_197; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_198 = proc_2_io_pipe_phv_out_data_198; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_199 = proc_2_io_pipe_phv_out_data_199; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_200 = proc_2_io_pipe_phv_out_data_200; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_201 = proc_2_io_pipe_phv_out_data_201; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_202 = proc_2_io_pipe_phv_out_data_202; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_203 = proc_2_io_pipe_phv_out_data_203; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_204 = proc_2_io_pipe_phv_out_data_204; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_205 = proc_2_io_pipe_phv_out_data_205; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_206 = proc_2_io_pipe_phv_out_data_206; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_207 = proc_2_io_pipe_phv_out_data_207; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_208 = proc_2_io_pipe_phv_out_data_208; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_209 = proc_2_io_pipe_phv_out_data_209; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_210 = proc_2_io_pipe_phv_out_data_210; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_211 = proc_2_io_pipe_phv_out_data_211; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_212 = proc_2_io_pipe_phv_out_data_212; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_213 = proc_2_io_pipe_phv_out_data_213; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_214 = proc_2_io_pipe_phv_out_data_214; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_215 = proc_2_io_pipe_phv_out_data_215; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_216 = proc_2_io_pipe_phv_out_data_216; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_217 = proc_2_io_pipe_phv_out_data_217; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_218 = proc_2_io_pipe_phv_out_data_218; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_219 = proc_2_io_pipe_phv_out_data_219; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_220 = proc_2_io_pipe_phv_out_data_220; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_221 = proc_2_io_pipe_phv_out_data_221; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_222 = proc_2_io_pipe_phv_out_data_222; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_223 = proc_2_io_pipe_phv_out_data_223; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_224 = proc_2_io_pipe_phv_out_data_224; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_225 = proc_2_io_pipe_phv_out_data_225; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_226 = proc_2_io_pipe_phv_out_data_226; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_227 = proc_2_io_pipe_phv_out_data_227; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_228 = proc_2_io_pipe_phv_out_data_228; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_229 = proc_2_io_pipe_phv_out_data_229; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_230 = proc_2_io_pipe_phv_out_data_230; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_231 = proc_2_io_pipe_phv_out_data_231; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_232 = proc_2_io_pipe_phv_out_data_232; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_233 = proc_2_io_pipe_phv_out_data_233; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_234 = proc_2_io_pipe_phv_out_data_234; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_235 = proc_2_io_pipe_phv_out_data_235; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_236 = proc_2_io_pipe_phv_out_data_236; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_237 = proc_2_io_pipe_phv_out_data_237; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_238 = proc_2_io_pipe_phv_out_data_238; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_239 = proc_2_io_pipe_phv_out_data_239; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_240 = proc_2_io_pipe_phv_out_data_240; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_241 = proc_2_io_pipe_phv_out_data_241; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_242 = proc_2_io_pipe_phv_out_data_242; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_243 = proc_2_io_pipe_phv_out_data_243; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_244 = proc_2_io_pipe_phv_out_data_244; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_245 = proc_2_io_pipe_phv_out_data_245; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_246 = proc_2_io_pipe_phv_out_data_246; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_247 = proc_2_io_pipe_phv_out_data_247; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_248 = proc_2_io_pipe_phv_out_data_248; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_249 = proc_2_io_pipe_phv_out_data_249; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_250 = proc_2_io_pipe_phv_out_data_250; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_251 = proc_2_io_pipe_phv_out_data_251; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_252 = proc_2_io_pipe_phv_out_data_252; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_253 = proc_2_io_pipe_phv_out_data_253; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_254 = proc_2_io_pipe_phv_out_data_254; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_255 = proc_2_io_pipe_phv_out_data_255; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_next_processor_id = proc_2_io_pipe_phv_out_next_processor_id; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_next_config_id = proc_2_io_pipe_phv_out_next_config_id; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_is_valid_processor = 4'h3 == proc_2_io_pipe_phv_out_next_processor_id; // @[pisa.scala 36:62]
  assign proc_3_io_mod_mat_mod_en = io_mod_proc_mod_3_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_config_id = io_mod_proc_mod_3_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_3_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_3_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_3_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_3_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_3_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_3_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_3_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_3_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_3_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_3_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_3_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_3_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_3_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_w_en = io_mod_proc_mod_3_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_3_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_w_addr = io_mod_proc_mod_3_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_w_data = io_mod_proc_mod_3_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_3_io_mod_exe_mod_en_0 = io_mod_proc_mod_3_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_3_io_mod_exe_mod_en_1 = io_mod_proc_mod_3_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_3_io_mod_exe_mod_addr = io_mod_proc_mod_3_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_3_io_mod_exe_mod_data_0 = io_mod_proc_mod_3_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_3_io_mod_exe_mod_data_1 = io_mod_proc_mod_3_exe_mod_data_1; // @[pisa.scala 29:20]
  assign proc_4_clock = clock;
  assign proc_4_io_pipe_phv_in_data_0 = proc_3_io_pipe_phv_out_data_0; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_1 = proc_3_io_pipe_phv_out_data_1; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_2 = proc_3_io_pipe_phv_out_data_2; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_3 = proc_3_io_pipe_phv_out_data_3; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_4 = proc_3_io_pipe_phv_out_data_4; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_5 = proc_3_io_pipe_phv_out_data_5; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_6 = proc_3_io_pipe_phv_out_data_6; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_7 = proc_3_io_pipe_phv_out_data_7; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_8 = proc_3_io_pipe_phv_out_data_8; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_9 = proc_3_io_pipe_phv_out_data_9; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_10 = proc_3_io_pipe_phv_out_data_10; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_11 = proc_3_io_pipe_phv_out_data_11; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_12 = proc_3_io_pipe_phv_out_data_12; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_13 = proc_3_io_pipe_phv_out_data_13; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_14 = proc_3_io_pipe_phv_out_data_14; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_15 = proc_3_io_pipe_phv_out_data_15; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_16 = proc_3_io_pipe_phv_out_data_16; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_17 = proc_3_io_pipe_phv_out_data_17; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_18 = proc_3_io_pipe_phv_out_data_18; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_19 = proc_3_io_pipe_phv_out_data_19; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_20 = proc_3_io_pipe_phv_out_data_20; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_21 = proc_3_io_pipe_phv_out_data_21; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_22 = proc_3_io_pipe_phv_out_data_22; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_23 = proc_3_io_pipe_phv_out_data_23; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_24 = proc_3_io_pipe_phv_out_data_24; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_25 = proc_3_io_pipe_phv_out_data_25; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_26 = proc_3_io_pipe_phv_out_data_26; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_27 = proc_3_io_pipe_phv_out_data_27; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_28 = proc_3_io_pipe_phv_out_data_28; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_29 = proc_3_io_pipe_phv_out_data_29; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_30 = proc_3_io_pipe_phv_out_data_30; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_31 = proc_3_io_pipe_phv_out_data_31; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_32 = proc_3_io_pipe_phv_out_data_32; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_33 = proc_3_io_pipe_phv_out_data_33; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_34 = proc_3_io_pipe_phv_out_data_34; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_35 = proc_3_io_pipe_phv_out_data_35; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_36 = proc_3_io_pipe_phv_out_data_36; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_37 = proc_3_io_pipe_phv_out_data_37; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_38 = proc_3_io_pipe_phv_out_data_38; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_39 = proc_3_io_pipe_phv_out_data_39; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_40 = proc_3_io_pipe_phv_out_data_40; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_41 = proc_3_io_pipe_phv_out_data_41; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_42 = proc_3_io_pipe_phv_out_data_42; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_43 = proc_3_io_pipe_phv_out_data_43; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_44 = proc_3_io_pipe_phv_out_data_44; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_45 = proc_3_io_pipe_phv_out_data_45; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_46 = proc_3_io_pipe_phv_out_data_46; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_47 = proc_3_io_pipe_phv_out_data_47; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_48 = proc_3_io_pipe_phv_out_data_48; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_49 = proc_3_io_pipe_phv_out_data_49; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_50 = proc_3_io_pipe_phv_out_data_50; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_51 = proc_3_io_pipe_phv_out_data_51; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_52 = proc_3_io_pipe_phv_out_data_52; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_53 = proc_3_io_pipe_phv_out_data_53; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_54 = proc_3_io_pipe_phv_out_data_54; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_55 = proc_3_io_pipe_phv_out_data_55; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_56 = proc_3_io_pipe_phv_out_data_56; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_57 = proc_3_io_pipe_phv_out_data_57; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_58 = proc_3_io_pipe_phv_out_data_58; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_59 = proc_3_io_pipe_phv_out_data_59; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_60 = proc_3_io_pipe_phv_out_data_60; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_61 = proc_3_io_pipe_phv_out_data_61; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_62 = proc_3_io_pipe_phv_out_data_62; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_63 = proc_3_io_pipe_phv_out_data_63; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_64 = proc_3_io_pipe_phv_out_data_64; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_65 = proc_3_io_pipe_phv_out_data_65; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_66 = proc_3_io_pipe_phv_out_data_66; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_67 = proc_3_io_pipe_phv_out_data_67; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_68 = proc_3_io_pipe_phv_out_data_68; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_69 = proc_3_io_pipe_phv_out_data_69; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_70 = proc_3_io_pipe_phv_out_data_70; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_71 = proc_3_io_pipe_phv_out_data_71; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_72 = proc_3_io_pipe_phv_out_data_72; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_73 = proc_3_io_pipe_phv_out_data_73; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_74 = proc_3_io_pipe_phv_out_data_74; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_75 = proc_3_io_pipe_phv_out_data_75; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_76 = proc_3_io_pipe_phv_out_data_76; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_77 = proc_3_io_pipe_phv_out_data_77; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_78 = proc_3_io_pipe_phv_out_data_78; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_79 = proc_3_io_pipe_phv_out_data_79; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_80 = proc_3_io_pipe_phv_out_data_80; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_81 = proc_3_io_pipe_phv_out_data_81; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_82 = proc_3_io_pipe_phv_out_data_82; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_83 = proc_3_io_pipe_phv_out_data_83; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_84 = proc_3_io_pipe_phv_out_data_84; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_85 = proc_3_io_pipe_phv_out_data_85; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_86 = proc_3_io_pipe_phv_out_data_86; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_87 = proc_3_io_pipe_phv_out_data_87; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_88 = proc_3_io_pipe_phv_out_data_88; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_89 = proc_3_io_pipe_phv_out_data_89; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_90 = proc_3_io_pipe_phv_out_data_90; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_91 = proc_3_io_pipe_phv_out_data_91; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_92 = proc_3_io_pipe_phv_out_data_92; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_93 = proc_3_io_pipe_phv_out_data_93; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_94 = proc_3_io_pipe_phv_out_data_94; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_95 = proc_3_io_pipe_phv_out_data_95; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_96 = proc_3_io_pipe_phv_out_data_96; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_97 = proc_3_io_pipe_phv_out_data_97; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_98 = proc_3_io_pipe_phv_out_data_98; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_99 = proc_3_io_pipe_phv_out_data_99; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_100 = proc_3_io_pipe_phv_out_data_100; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_101 = proc_3_io_pipe_phv_out_data_101; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_102 = proc_3_io_pipe_phv_out_data_102; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_103 = proc_3_io_pipe_phv_out_data_103; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_104 = proc_3_io_pipe_phv_out_data_104; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_105 = proc_3_io_pipe_phv_out_data_105; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_106 = proc_3_io_pipe_phv_out_data_106; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_107 = proc_3_io_pipe_phv_out_data_107; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_108 = proc_3_io_pipe_phv_out_data_108; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_109 = proc_3_io_pipe_phv_out_data_109; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_110 = proc_3_io_pipe_phv_out_data_110; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_111 = proc_3_io_pipe_phv_out_data_111; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_112 = proc_3_io_pipe_phv_out_data_112; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_113 = proc_3_io_pipe_phv_out_data_113; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_114 = proc_3_io_pipe_phv_out_data_114; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_115 = proc_3_io_pipe_phv_out_data_115; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_116 = proc_3_io_pipe_phv_out_data_116; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_117 = proc_3_io_pipe_phv_out_data_117; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_118 = proc_3_io_pipe_phv_out_data_118; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_119 = proc_3_io_pipe_phv_out_data_119; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_120 = proc_3_io_pipe_phv_out_data_120; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_121 = proc_3_io_pipe_phv_out_data_121; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_122 = proc_3_io_pipe_phv_out_data_122; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_123 = proc_3_io_pipe_phv_out_data_123; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_124 = proc_3_io_pipe_phv_out_data_124; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_125 = proc_3_io_pipe_phv_out_data_125; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_126 = proc_3_io_pipe_phv_out_data_126; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_127 = proc_3_io_pipe_phv_out_data_127; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_128 = proc_3_io_pipe_phv_out_data_128; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_129 = proc_3_io_pipe_phv_out_data_129; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_130 = proc_3_io_pipe_phv_out_data_130; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_131 = proc_3_io_pipe_phv_out_data_131; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_132 = proc_3_io_pipe_phv_out_data_132; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_133 = proc_3_io_pipe_phv_out_data_133; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_134 = proc_3_io_pipe_phv_out_data_134; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_135 = proc_3_io_pipe_phv_out_data_135; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_136 = proc_3_io_pipe_phv_out_data_136; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_137 = proc_3_io_pipe_phv_out_data_137; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_138 = proc_3_io_pipe_phv_out_data_138; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_139 = proc_3_io_pipe_phv_out_data_139; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_140 = proc_3_io_pipe_phv_out_data_140; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_141 = proc_3_io_pipe_phv_out_data_141; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_142 = proc_3_io_pipe_phv_out_data_142; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_143 = proc_3_io_pipe_phv_out_data_143; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_144 = proc_3_io_pipe_phv_out_data_144; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_145 = proc_3_io_pipe_phv_out_data_145; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_146 = proc_3_io_pipe_phv_out_data_146; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_147 = proc_3_io_pipe_phv_out_data_147; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_148 = proc_3_io_pipe_phv_out_data_148; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_149 = proc_3_io_pipe_phv_out_data_149; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_150 = proc_3_io_pipe_phv_out_data_150; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_151 = proc_3_io_pipe_phv_out_data_151; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_152 = proc_3_io_pipe_phv_out_data_152; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_153 = proc_3_io_pipe_phv_out_data_153; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_154 = proc_3_io_pipe_phv_out_data_154; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_155 = proc_3_io_pipe_phv_out_data_155; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_156 = proc_3_io_pipe_phv_out_data_156; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_157 = proc_3_io_pipe_phv_out_data_157; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_158 = proc_3_io_pipe_phv_out_data_158; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_159 = proc_3_io_pipe_phv_out_data_159; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_160 = proc_3_io_pipe_phv_out_data_160; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_161 = proc_3_io_pipe_phv_out_data_161; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_162 = proc_3_io_pipe_phv_out_data_162; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_163 = proc_3_io_pipe_phv_out_data_163; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_164 = proc_3_io_pipe_phv_out_data_164; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_165 = proc_3_io_pipe_phv_out_data_165; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_166 = proc_3_io_pipe_phv_out_data_166; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_167 = proc_3_io_pipe_phv_out_data_167; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_168 = proc_3_io_pipe_phv_out_data_168; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_169 = proc_3_io_pipe_phv_out_data_169; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_170 = proc_3_io_pipe_phv_out_data_170; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_171 = proc_3_io_pipe_phv_out_data_171; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_172 = proc_3_io_pipe_phv_out_data_172; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_173 = proc_3_io_pipe_phv_out_data_173; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_174 = proc_3_io_pipe_phv_out_data_174; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_175 = proc_3_io_pipe_phv_out_data_175; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_176 = proc_3_io_pipe_phv_out_data_176; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_177 = proc_3_io_pipe_phv_out_data_177; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_178 = proc_3_io_pipe_phv_out_data_178; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_179 = proc_3_io_pipe_phv_out_data_179; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_180 = proc_3_io_pipe_phv_out_data_180; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_181 = proc_3_io_pipe_phv_out_data_181; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_182 = proc_3_io_pipe_phv_out_data_182; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_183 = proc_3_io_pipe_phv_out_data_183; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_184 = proc_3_io_pipe_phv_out_data_184; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_185 = proc_3_io_pipe_phv_out_data_185; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_186 = proc_3_io_pipe_phv_out_data_186; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_187 = proc_3_io_pipe_phv_out_data_187; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_188 = proc_3_io_pipe_phv_out_data_188; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_189 = proc_3_io_pipe_phv_out_data_189; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_190 = proc_3_io_pipe_phv_out_data_190; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_191 = proc_3_io_pipe_phv_out_data_191; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_192 = proc_3_io_pipe_phv_out_data_192; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_193 = proc_3_io_pipe_phv_out_data_193; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_194 = proc_3_io_pipe_phv_out_data_194; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_195 = proc_3_io_pipe_phv_out_data_195; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_196 = proc_3_io_pipe_phv_out_data_196; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_197 = proc_3_io_pipe_phv_out_data_197; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_198 = proc_3_io_pipe_phv_out_data_198; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_199 = proc_3_io_pipe_phv_out_data_199; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_200 = proc_3_io_pipe_phv_out_data_200; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_201 = proc_3_io_pipe_phv_out_data_201; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_202 = proc_3_io_pipe_phv_out_data_202; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_203 = proc_3_io_pipe_phv_out_data_203; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_204 = proc_3_io_pipe_phv_out_data_204; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_205 = proc_3_io_pipe_phv_out_data_205; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_206 = proc_3_io_pipe_phv_out_data_206; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_207 = proc_3_io_pipe_phv_out_data_207; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_208 = proc_3_io_pipe_phv_out_data_208; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_209 = proc_3_io_pipe_phv_out_data_209; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_210 = proc_3_io_pipe_phv_out_data_210; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_211 = proc_3_io_pipe_phv_out_data_211; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_212 = proc_3_io_pipe_phv_out_data_212; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_213 = proc_3_io_pipe_phv_out_data_213; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_214 = proc_3_io_pipe_phv_out_data_214; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_215 = proc_3_io_pipe_phv_out_data_215; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_216 = proc_3_io_pipe_phv_out_data_216; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_217 = proc_3_io_pipe_phv_out_data_217; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_218 = proc_3_io_pipe_phv_out_data_218; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_219 = proc_3_io_pipe_phv_out_data_219; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_220 = proc_3_io_pipe_phv_out_data_220; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_221 = proc_3_io_pipe_phv_out_data_221; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_222 = proc_3_io_pipe_phv_out_data_222; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_223 = proc_3_io_pipe_phv_out_data_223; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_224 = proc_3_io_pipe_phv_out_data_224; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_225 = proc_3_io_pipe_phv_out_data_225; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_226 = proc_3_io_pipe_phv_out_data_226; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_227 = proc_3_io_pipe_phv_out_data_227; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_228 = proc_3_io_pipe_phv_out_data_228; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_229 = proc_3_io_pipe_phv_out_data_229; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_230 = proc_3_io_pipe_phv_out_data_230; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_231 = proc_3_io_pipe_phv_out_data_231; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_232 = proc_3_io_pipe_phv_out_data_232; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_233 = proc_3_io_pipe_phv_out_data_233; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_234 = proc_3_io_pipe_phv_out_data_234; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_235 = proc_3_io_pipe_phv_out_data_235; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_236 = proc_3_io_pipe_phv_out_data_236; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_237 = proc_3_io_pipe_phv_out_data_237; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_238 = proc_3_io_pipe_phv_out_data_238; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_239 = proc_3_io_pipe_phv_out_data_239; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_240 = proc_3_io_pipe_phv_out_data_240; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_241 = proc_3_io_pipe_phv_out_data_241; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_242 = proc_3_io_pipe_phv_out_data_242; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_243 = proc_3_io_pipe_phv_out_data_243; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_244 = proc_3_io_pipe_phv_out_data_244; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_245 = proc_3_io_pipe_phv_out_data_245; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_246 = proc_3_io_pipe_phv_out_data_246; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_247 = proc_3_io_pipe_phv_out_data_247; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_248 = proc_3_io_pipe_phv_out_data_248; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_249 = proc_3_io_pipe_phv_out_data_249; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_250 = proc_3_io_pipe_phv_out_data_250; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_251 = proc_3_io_pipe_phv_out_data_251; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_252 = proc_3_io_pipe_phv_out_data_252; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_253 = proc_3_io_pipe_phv_out_data_253; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_254 = proc_3_io_pipe_phv_out_data_254; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_255 = proc_3_io_pipe_phv_out_data_255; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_next_processor_id = proc_3_io_pipe_phv_out_next_processor_id; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_next_config_id = proc_3_io_pipe_phv_out_next_config_id; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_is_valid_processor = 4'h4 == proc_3_io_pipe_phv_out_next_processor_id; // @[pisa.scala 36:62]
  assign proc_4_io_mod_mat_mod_en = io_mod_proc_mod_4_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_config_id = io_mod_proc_mod_4_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_4_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_4_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_4_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_4_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_4_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_4_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_4_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_4_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_4_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_4_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_4_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_4_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_4_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_w_en = io_mod_proc_mod_4_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_4_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_w_addr = io_mod_proc_mod_4_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_w_data = io_mod_proc_mod_4_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_4_io_mod_exe_mod_en_0 = io_mod_proc_mod_4_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_4_io_mod_exe_mod_en_1 = io_mod_proc_mod_4_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_4_io_mod_exe_mod_addr = io_mod_proc_mod_4_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_4_io_mod_exe_mod_data_0 = io_mod_proc_mod_4_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_4_io_mod_exe_mod_data_1 = io_mod_proc_mod_4_exe_mod_data_1; // @[pisa.scala 29:20]
  assign proc_5_clock = clock;
  assign proc_5_io_pipe_phv_in_data_0 = proc_4_io_pipe_phv_out_data_0; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_1 = proc_4_io_pipe_phv_out_data_1; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_2 = proc_4_io_pipe_phv_out_data_2; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_3 = proc_4_io_pipe_phv_out_data_3; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_4 = proc_4_io_pipe_phv_out_data_4; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_5 = proc_4_io_pipe_phv_out_data_5; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_6 = proc_4_io_pipe_phv_out_data_6; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_7 = proc_4_io_pipe_phv_out_data_7; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_8 = proc_4_io_pipe_phv_out_data_8; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_9 = proc_4_io_pipe_phv_out_data_9; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_10 = proc_4_io_pipe_phv_out_data_10; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_11 = proc_4_io_pipe_phv_out_data_11; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_12 = proc_4_io_pipe_phv_out_data_12; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_13 = proc_4_io_pipe_phv_out_data_13; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_14 = proc_4_io_pipe_phv_out_data_14; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_15 = proc_4_io_pipe_phv_out_data_15; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_16 = proc_4_io_pipe_phv_out_data_16; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_17 = proc_4_io_pipe_phv_out_data_17; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_18 = proc_4_io_pipe_phv_out_data_18; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_19 = proc_4_io_pipe_phv_out_data_19; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_20 = proc_4_io_pipe_phv_out_data_20; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_21 = proc_4_io_pipe_phv_out_data_21; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_22 = proc_4_io_pipe_phv_out_data_22; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_23 = proc_4_io_pipe_phv_out_data_23; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_24 = proc_4_io_pipe_phv_out_data_24; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_25 = proc_4_io_pipe_phv_out_data_25; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_26 = proc_4_io_pipe_phv_out_data_26; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_27 = proc_4_io_pipe_phv_out_data_27; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_28 = proc_4_io_pipe_phv_out_data_28; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_29 = proc_4_io_pipe_phv_out_data_29; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_30 = proc_4_io_pipe_phv_out_data_30; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_31 = proc_4_io_pipe_phv_out_data_31; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_32 = proc_4_io_pipe_phv_out_data_32; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_33 = proc_4_io_pipe_phv_out_data_33; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_34 = proc_4_io_pipe_phv_out_data_34; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_35 = proc_4_io_pipe_phv_out_data_35; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_36 = proc_4_io_pipe_phv_out_data_36; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_37 = proc_4_io_pipe_phv_out_data_37; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_38 = proc_4_io_pipe_phv_out_data_38; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_39 = proc_4_io_pipe_phv_out_data_39; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_40 = proc_4_io_pipe_phv_out_data_40; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_41 = proc_4_io_pipe_phv_out_data_41; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_42 = proc_4_io_pipe_phv_out_data_42; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_43 = proc_4_io_pipe_phv_out_data_43; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_44 = proc_4_io_pipe_phv_out_data_44; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_45 = proc_4_io_pipe_phv_out_data_45; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_46 = proc_4_io_pipe_phv_out_data_46; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_47 = proc_4_io_pipe_phv_out_data_47; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_48 = proc_4_io_pipe_phv_out_data_48; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_49 = proc_4_io_pipe_phv_out_data_49; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_50 = proc_4_io_pipe_phv_out_data_50; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_51 = proc_4_io_pipe_phv_out_data_51; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_52 = proc_4_io_pipe_phv_out_data_52; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_53 = proc_4_io_pipe_phv_out_data_53; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_54 = proc_4_io_pipe_phv_out_data_54; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_55 = proc_4_io_pipe_phv_out_data_55; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_56 = proc_4_io_pipe_phv_out_data_56; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_57 = proc_4_io_pipe_phv_out_data_57; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_58 = proc_4_io_pipe_phv_out_data_58; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_59 = proc_4_io_pipe_phv_out_data_59; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_60 = proc_4_io_pipe_phv_out_data_60; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_61 = proc_4_io_pipe_phv_out_data_61; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_62 = proc_4_io_pipe_phv_out_data_62; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_63 = proc_4_io_pipe_phv_out_data_63; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_64 = proc_4_io_pipe_phv_out_data_64; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_65 = proc_4_io_pipe_phv_out_data_65; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_66 = proc_4_io_pipe_phv_out_data_66; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_67 = proc_4_io_pipe_phv_out_data_67; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_68 = proc_4_io_pipe_phv_out_data_68; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_69 = proc_4_io_pipe_phv_out_data_69; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_70 = proc_4_io_pipe_phv_out_data_70; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_71 = proc_4_io_pipe_phv_out_data_71; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_72 = proc_4_io_pipe_phv_out_data_72; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_73 = proc_4_io_pipe_phv_out_data_73; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_74 = proc_4_io_pipe_phv_out_data_74; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_75 = proc_4_io_pipe_phv_out_data_75; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_76 = proc_4_io_pipe_phv_out_data_76; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_77 = proc_4_io_pipe_phv_out_data_77; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_78 = proc_4_io_pipe_phv_out_data_78; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_79 = proc_4_io_pipe_phv_out_data_79; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_80 = proc_4_io_pipe_phv_out_data_80; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_81 = proc_4_io_pipe_phv_out_data_81; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_82 = proc_4_io_pipe_phv_out_data_82; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_83 = proc_4_io_pipe_phv_out_data_83; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_84 = proc_4_io_pipe_phv_out_data_84; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_85 = proc_4_io_pipe_phv_out_data_85; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_86 = proc_4_io_pipe_phv_out_data_86; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_87 = proc_4_io_pipe_phv_out_data_87; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_88 = proc_4_io_pipe_phv_out_data_88; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_89 = proc_4_io_pipe_phv_out_data_89; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_90 = proc_4_io_pipe_phv_out_data_90; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_91 = proc_4_io_pipe_phv_out_data_91; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_92 = proc_4_io_pipe_phv_out_data_92; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_93 = proc_4_io_pipe_phv_out_data_93; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_94 = proc_4_io_pipe_phv_out_data_94; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_95 = proc_4_io_pipe_phv_out_data_95; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_96 = proc_4_io_pipe_phv_out_data_96; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_97 = proc_4_io_pipe_phv_out_data_97; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_98 = proc_4_io_pipe_phv_out_data_98; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_99 = proc_4_io_pipe_phv_out_data_99; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_100 = proc_4_io_pipe_phv_out_data_100; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_101 = proc_4_io_pipe_phv_out_data_101; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_102 = proc_4_io_pipe_phv_out_data_102; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_103 = proc_4_io_pipe_phv_out_data_103; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_104 = proc_4_io_pipe_phv_out_data_104; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_105 = proc_4_io_pipe_phv_out_data_105; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_106 = proc_4_io_pipe_phv_out_data_106; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_107 = proc_4_io_pipe_phv_out_data_107; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_108 = proc_4_io_pipe_phv_out_data_108; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_109 = proc_4_io_pipe_phv_out_data_109; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_110 = proc_4_io_pipe_phv_out_data_110; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_111 = proc_4_io_pipe_phv_out_data_111; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_112 = proc_4_io_pipe_phv_out_data_112; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_113 = proc_4_io_pipe_phv_out_data_113; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_114 = proc_4_io_pipe_phv_out_data_114; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_115 = proc_4_io_pipe_phv_out_data_115; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_116 = proc_4_io_pipe_phv_out_data_116; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_117 = proc_4_io_pipe_phv_out_data_117; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_118 = proc_4_io_pipe_phv_out_data_118; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_119 = proc_4_io_pipe_phv_out_data_119; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_120 = proc_4_io_pipe_phv_out_data_120; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_121 = proc_4_io_pipe_phv_out_data_121; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_122 = proc_4_io_pipe_phv_out_data_122; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_123 = proc_4_io_pipe_phv_out_data_123; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_124 = proc_4_io_pipe_phv_out_data_124; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_125 = proc_4_io_pipe_phv_out_data_125; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_126 = proc_4_io_pipe_phv_out_data_126; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_127 = proc_4_io_pipe_phv_out_data_127; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_128 = proc_4_io_pipe_phv_out_data_128; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_129 = proc_4_io_pipe_phv_out_data_129; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_130 = proc_4_io_pipe_phv_out_data_130; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_131 = proc_4_io_pipe_phv_out_data_131; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_132 = proc_4_io_pipe_phv_out_data_132; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_133 = proc_4_io_pipe_phv_out_data_133; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_134 = proc_4_io_pipe_phv_out_data_134; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_135 = proc_4_io_pipe_phv_out_data_135; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_136 = proc_4_io_pipe_phv_out_data_136; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_137 = proc_4_io_pipe_phv_out_data_137; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_138 = proc_4_io_pipe_phv_out_data_138; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_139 = proc_4_io_pipe_phv_out_data_139; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_140 = proc_4_io_pipe_phv_out_data_140; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_141 = proc_4_io_pipe_phv_out_data_141; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_142 = proc_4_io_pipe_phv_out_data_142; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_143 = proc_4_io_pipe_phv_out_data_143; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_144 = proc_4_io_pipe_phv_out_data_144; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_145 = proc_4_io_pipe_phv_out_data_145; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_146 = proc_4_io_pipe_phv_out_data_146; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_147 = proc_4_io_pipe_phv_out_data_147; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_148 = proc_4_io_pipe_phv_out_data_148; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_149 = proc_4_io_pipe_phv_out_data_149; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_150 = proc_4_io_pipe_phv_out_data_150; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_151 = proc_4_io_pipe_phv_out_data_151; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_152 = proc_4_io_pipe_phv_out_data_152; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_153 = proc_4_io_pipe_phv_out_data_153; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_154 = proc_4_io_pipe_phv_out_data_154; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_155 = proc_4_io_pipe_phv_out_data_155; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_156 = proc_4_io_pipe_phv_out_data_156; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_157 = proc_4_io_pipe_phv_out_data_157; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_158 = proc_4_io_pipe_phv_out_data_158; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_159 = proc_4_io_pipe_phv_out_data_159; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_160 = proc_4_io_pipe_phv_out_data_160; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_161 = proc_4_io_pipe_phv_out_data_161; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_162 = proc_4_io_pipe_phv_out_data_162; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_163 = proc_4_io_pipe_phv_out_data_163; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_164 = proc_4_io_pipe_phv_out_data_164; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_165 = proc_4_io_pipe_phv_out_data_165; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_166 = proc_4_io_pipe_phv_out_data_166; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_167 = proc_4_io_pipe_phv_out_data_167; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_168 = proc_4_io_pipe_phv_out_data_168; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_169 = proc_4_io_pipe_phv_out_data_169; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_170 = proc_4_io_pipe_phv_out_data_170; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_171 = proc_4_io_pipe_phv_out_data_171; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_172 = proc_4_io_pipe_phv_out_data_172; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_173 = proc_4_io_pipe_phv_out_data_173; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_174 = proc_4_io_pipe_phv_out_data_174; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_175 = proc_4_io_pipe_phv_out_data_175; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_176 = proc_4_io_pipe_phv_out_data_176; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_177 = proc_4_io_pipe_phv_out_data_177; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_178 = proc_4_io_pipe_phv_out_data_178; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_179 = proc_4_io_pipe_phv_out_data_179; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_180 = proc_4_io_pipe_phv_out_data_180; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_181 = proc_4_io_pipe_phv_out_data_181; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_182 = proc_4_io_pipe_phv_out_data_182; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_183 = proc_4_io_pipe_phv_out_data_183; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_184 = proc_4_io_pipe_phv_out_data_184; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_185 = proc_4_io_pipe_phv_out_data_185; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_186 = proc_4_io_pipe_phv_out_data_186; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_187 = proc_4_io_pipe_phv_out_data_187; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_188 = proc_4_io_pipe_phv_out_data_188; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_189 = proc_4_io_pipe_phv_out_data_189; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_190 = proc_4_io_pipe_phv_out_data_190; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_191 = proc_4_io_pipe_phv_out_data_191; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_192 = proc_4_io_pipe_phv_out_data_192; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_193 = proc_4_io_pipe_phv_out_data_193; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_194 = proc_4_io_pipe_phv_out_data_194; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_195 = proc_4_io_pipe_phv_out_data_195; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_196 = proc_4_io_pipe_phv_out_data_196; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_197 = proc_4_io_pipe_phv_out_data_197; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_198 = proc_4_io_pipe_phv_out_data_198; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_199 = proc_4_io_pipe_phv_out_data_199; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_200 = proc_4_io_pipe_phv_out_data_200; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_201 = proc_4_io_pipe_phv_out_data_201; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_202 = proc_4_io_pipe_phv_out_data_202; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_203 = proc_4_io_pipe_phv_out_data_203; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_204 = proc_4_io_pipe_phv_out_data_204; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_205 = proc_4_io_pipe_phv_out_data_205; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_206 = proc_4_io_pipe_phv_out_data_206; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_207 = proc_4_io_pipe_phv_out_data_207; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_208 = proc_4_io_pipe_phv_out_data_208; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_209 = proc_4_io_pipe_phv_out_data_209; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_210 = proc_4_io_pipe_phv_out_data_210; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_211 = proc_4_io_pipe_phv_out_data_211; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_212 = proc_4_io_pipe_phv_out_data_212; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_213 = proc_4_io_pipe_phv_out_data_213; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_214 = proc_4_io_pipe_phv_out_data_214; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_215 = proc_4_io_pipe_phv_out_data_215; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_216 = proc_4_io_pipe_phv_out_data_216; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_217 = proc_4_io_pipe_phv_out_data_217; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_218 = proc_4_io_pipe_phv_out_data_218; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_219 = proc_4_io_pipe_phv_out_data_219; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_220 = proc_4_io_pipe_phv_out_data_220; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_221 = proc_4_io_pipe_phv_out_data_221; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_222 = proc_4_io_pipe_phv_out_data_222; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_223 = proc_4_io_pipe_phv_out_data_223; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_224 = proc_4_io_pipe_phv_out_data_224; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_225 = proc_4_io_pipe_phv_out_data_225; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_226 = proc_4_io_pipe_phv_out_data_226; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_227 = proc_4_io_pipe_phv_out_data_227; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_228 = proc_4_io_pipe_phv_out_data_228; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_229 = proc_4_io_pipe_phv_out_data_229; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_230 = proc_4_io_pipe_phv_out_data_230; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_231 = proc_4_io_pipe_phv_out_data_231; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_232 = proc_4_io_pipe_phv_out_data_232; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_233 = proc_4_io_pipe_phv_out_data_233; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_234 = proc_4_io_pipe_phv_out_data_234; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_235 = proc_4_io_pipe_phv_out_data_235; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_236 = proc_4_io_pipe_phv_out_data_236; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_237 = proc_4_io_pipe_phv_out_data_237; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_238 = proc_4_io_pipe_phv_out_data_238; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_239 = proc_4_io_pipe_phv_out_data_239; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_240 = proc_4_io_pipe_phv_out_data_240; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_241 = proc_4_io_pipe_phv_out_data_241; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_242 = proc_4_io_pipe_phv_out_data_242; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_243 = proc_4_io_pipe_phv_out_data_243; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_244 = proc_4_io_pipe_phv_out_data_244; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_245 = proc_4_io_pipe_phv_out_data_245; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_246 = proc_4_io_pipe_phv_out_data_246; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_247 = proc_4_io_pipe_phv_out_data_247; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_248 = proc_4_io_pipe_phv_out_data_248; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_249 = proc_4_io_pipe_phv_out_data_249; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_250 = proc_4_io_pipe_phv_out_data_250; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_251 = proc_4_io_pipe_phv_out_data_251; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_252 = proc_4_io_pipe_phv_out_data_252; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_253 = proc_4_io_pipe_phv_out_data_253; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_254 = proc_4_io_pipe_phv_out_data_254; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_255 = proc_4_io_pipe_phv_out_data_255; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_next_processor_id = proc_4_io_pipe_phv_out_next_processor_id; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_next_config_id = proc_4_io_pipe_phv_out_next_config_id; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_is_valid_processor = 4'h5 == proc_4_io_pipe_phv_out_next_processor_id; // @[pisa.scala 36:62]
  assign proc_5_io_mod_mat_mod_en = io_mod_proc_mod_5_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_config_id = io_mod_proc_mod_5_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_5_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_5_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_5_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_5_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_5_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_5_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_5_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_5_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_5_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_5_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_5_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_5_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_5_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_w_en = io_mod_proc_mod_5_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_5_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_w_addr = io_mod_proc_mod_5_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_w_data = io_mod_proc_mod_5_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_5_io_mod_exe_mod_en_0 = io_mod_proc_mod_5_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_5_io_mod_exe_mod_en_1 = io_mod_proc_mod_5_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_5_io_mod_exe_mod_addr = io_mod_proc_mod_5_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_5_io_mod_exe_mod_data_0 = io_mod_proc_mod_5_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_5_io_mod_exe_mod_data_1 = io_mod_proc_mod_5_exe_mod_data_1; // @[pisa.scala 29:20]
  assign proc_6_clock = clock;
  assign proc_6_io_pipe_phv_in_data_0 = proc_5_io_pipe_phv_out_data_0; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_1 = proc_5_io_pipe_phv_out_data_1; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_2 = proc_5_io_pipe_phv_out_data_2; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_3 = proc_5_io_pipe_phv_out_data_3; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_4 = proc_5_io_pipe_phv_out_data_4; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_5 = proc_5_io_pipe_phv_out_data_5; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_6 = proc_5_io_pipe_phv_out_data_6; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_7 = proc_5_io_pipe_phv_out_data_7; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_8 = proc_5_io_pipe_phv_out_data_8; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_9 = proc_5_io_pipe_phv_out_data_9; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_10 = proc_5_io_pipe_phv_out_data_10; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_11 = proc_5_io_pipe_phv_out_data_11; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_12 = proc_5_io_pipe_phv_out_data_12; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_13 = proc_5_io_pipe_phv_out_data_13; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_14 = proc_5_io_pipe_phv_out_data_14; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_15 = proc_5_io_pipe_phv_out_data_15; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_16 = proc_5_io_pipe_phv_out_data_16; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_17 = proc_5_io_pipe_phv_out_data_17; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_18 = proc_5_io_pipe_phv_out_data_18; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_19 = proc_5_io_pipe_phv_out_data_19; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_20 = proc_5_io_pipe_phv_out_data_20; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_21 = proc_5_io_pipe_phv_out_data_21; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_22 = proc_5_io_pipe_phv_out_data_22; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_23 = proc_5_io_pipe_phv_out_data_23; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_24 = proc_5_io_pipe_phv_out_data_24; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_25 = proc_5_io_pipe_phv_out_data_25; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_26 = proc_5_io_pipe_phv_out_data_26; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_27 = proc_5_io_pipe_phv_out_data_27; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_28 = proc_5_io_pipe_phv_out_data_28; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_29 = proc_5_io_pipe_phv_out_data_29; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_30 = proc_5_io_pipe_phv_out_data_30; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_31 = proc_5_io_pipe_phv_out_data_31; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_32 = proc_5_io_pipe_phv_out_data_32; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_33 = proc_5_io_pipe_phv_out_data_33; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_34 = proc_5_io_pipe_phv_out_data_34; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_35 = proc_5_io_pipe_phv_out_data_35; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_36 = proc_5_io_pipe_phv_out_data_36; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_37 = proc_5_io_pipe_phv_out_data_37; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_38 = proc_5_io_pipe_phv_out_data_38; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_39 = proc_5_io_pipe_phv_out_data_39; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_40 = proc_5_io_pipe_phv_out_data_40; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_41 = proc_5_io_pipe_phv_out_data_41; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_42 = proc_5_io_pipe_phv_out_data_42; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_43 = proc_5_io_pipe_phv_out_data_43; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_44 = proc_5_io_pipe_phv_out_data_44; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_45 = proc_5_io_pipe_phv_out_data_45; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_46 = proc_5_io_pipe_phv_out_data_46; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_47 = proc_5_io_pipe_phv_out_data_47; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_48 = proc_5_io_pipe_phv_out_data_48; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_49 = proc_5_io_pipe_phv_out_data_49; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_50 = proc_5_io_pipe_phv_out_data_50; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_51 = proc_5_io_pipe_phv_out_data_51; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_52 = proc_5_io_pipe_phv_out_data_52; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_53 = proc_5_io_pipe_phv_out_data_53; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_54 = proc_5_io_pipe_phv_out_data_54; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_55 = proc_5_io_pipe_phv_out_data_55; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_56 = proc_5_io_pipe_phv_out_data_56; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_57 = proc_5_io_pipe_phv_out_data_57; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_58 = proc_5_io_pipe_phv_out_data_58; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_59 = proc_5_io_pipe_phv_out_data_59; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_60 = proc_5_io_pipe_phv_out_data_60; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_61 = proc_5_io_pipe_phv_out_data_61; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_62 = proc_5_io_pipe_phv_out_data_62; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_63 = proc_5_io_pipe_phv_out_data_63; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_64 = proc_5_io_pipe_phv_out_data_64; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_65 = proc_5_io_pipe_phv_out_data_65; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_66 = proc_5_io_pipe_phv_out_data_66; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_67 = proc_5_io_pipe_phv_out_data_67; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_68 = proc_5_io_pipe_phv_out_data_68; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_69 = proc_5_io_pipe_phv_out_data_69; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_70 = proc_5_io_pipe_phv_out_data_70; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_71 = proc_5_io_pipe_phv_out_data_71; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_72 = proc_5_io_pipe_phv_out_data_72; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_73 = proc_5_io_pipe_phv_out_data_73; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_74 = proc_5_io_pipe_phv_out_data_74; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_75 = proc_5_io_pipe_phv_out_data_75; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_76 = proc_5_io_pipe_phv_out_data_76; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_77 = proc_5_io_pipe_phv_out_data_77; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_78 = proc_5_io_pipe_phv_out_data_78; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_79 = proc_5_io_pipe_phv_out_data_79; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_80 = proc_5_io_pipe_phv_out_data_80; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_81 = proc_5_io_pipe_phv_out_data_81; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_82 = proc_5_io_pipe_phv_out_data_82; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_83 = proc_5_io_pipe_phv_out_data_83; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_84 = proc_5_io_pipe_phv_out_data_84; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_85 = proc_5_io_pipe_phv_out_data_85; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_86 = proc_5_io_pipe_phv_out_data_86; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_87 = proc_5_io_pipe_phv_out_data_87; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_88 = proc_5_io_pipe_phv_out_data_88; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_89 = proc_5_io_pipe_phv_out_data_89; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_90 = proc_5_io_pipe_phv_out_data_90; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_91 = proc_5_io_pipe_phv_out_data_91; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_92 = proc_5_io_pipe_phv_out_data_92; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_93 = proc_5_io_pipe_phv_out_data_93; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_94 = proc_5_io_pipe_phv_out_data_94; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_95 = proc_5_io_pipe_phv_out_data_95; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_96 = proc_5_io_pipe_phv_out_data_96; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_97 = proc_5_io_pipe_phv_out_data_97; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_98 = proc_5_io_pipe_phv_out_data_98; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_99 = proc_5_io_pipe_phv_out_data_99; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_100 = proc_5_io_pipe_phv_out_data_100; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_101 = proc_5_io_pipe_phv_out_data_101; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_102 = proc_5_io_pipe_phv_out_data_102; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_103 = proc_5_io_pipe_phv_out_data_103; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_104 = proc_5_io_pipe_phv_out_data_104; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_105 = proc_5_io_pipe_phv_out_data_105; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_106 = proc_5_io_pipe_phv_out_data_106; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_107 = proc_5_io_pipe_phv_out_data_107; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_108 = proc_5_io_pipe_phv_out_data_108; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_109 = proc_5_io_pipe_phv_out_data_109; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_110 = proc_5_io_pipe_phv_out_data_110; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_111 = proc_5_io_pipe_phv_out_data_111; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_112 = proc_5_io_pipe_phv_out_data_112; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_113 = proc_5_io_pipe_phv_out_data_113; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_114 = proc_5_io_pipe_phv_out_data_114; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_115 = proc_5_io_pipe_phv_out_data_115; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_116 = proc_5_io_pipe_phv_out_data_116; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_117 = proc_5_io_pipe_phv_out_data_117; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_118 = proc_5_io_pipe_phv_out_data_118; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_119 = proc_5_io_pipe_phv_out_data_119; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_120 = proc_5_io_pipe_phv_out_data_120; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_121 = proc_5_io_pipe_phv_out_data_121; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_122 = proc_5_io_pipe_phv_out_data_122; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_123 = proc_5_io_pipe_phv_out_data_123; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_124 = proc_5_io_pipe_phv_out_data_124; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_125 = proc_5_io_pipe_phv_out_data_125; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_126 = proc_5_io_pipe_phv_out_data_126; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_127 = proc_5_io_pipe_phv_out_data_127; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_128 = proc_5_io_pipe_phv_out_data_128; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_129 = proc_5_io_pipe_phv_out_data_129; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_130 = proc_5_io_pipe_phv_out_data_130; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_131 = proc_5_io_pipe_phv_out_data_131; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_132 = proc_5_io_pipe_phv_out_data_132; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_133 = proc_5_io_pipe_phv_out_data_133; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_134 = proc_5_io_pipe_phv_out_data_134; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_135 = proc_5_io_pipe_phv_out_data_135; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_136 = proc_5_io_pipe_phv_out_data_136; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_137 = proc_5_io_pipe_phv_out_data_137; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_138 = proc_5_io_pipe_phv_out_data_138; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_139 = proc_5_io_pipe_phv_out_data_139; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_140 = proc_5_io_pipe_phv_out_data_140; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_141 = proc_5_io_pipe_phv_out_data_141; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_142 = proc_5_io_pipe_phv_out_data_142; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_143 = proc_5_io_pipe_phv_out_data_143; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_144 = proc_5_io_pipe_phv_out_data_144; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_145 = proc_5_io_pipe_phv_out_data_145; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_146 = proc_5_io_pipe_phv_out_data_146; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_147 = proc_5_io_pipe_phv_out_data_147; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_148 = proc_5_io_pipe_phv_out_data_148; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_149 = proc_5_io_pipe_phv_out_data_149; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_150 = proc_5_io_pipe_phv_out_data_150; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_151 = proc_5_io_pipe_phv_out_data_151; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_152 = proc_5_io_pipe_phv_out_data_152; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_153 = proc_5_io_pipe_phv_out_data_153; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_154 = proc_5_io_pipe_phv_out_data_154; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_155 = proc_5_io_pipe_phv_out_data_155; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_156 = proc_5_io_pipe_phv_out_data_156; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_157 = proc_5_io_pipe_phv_out_data_157; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_158 = proc_5_io_pipe_phv_out_data_158; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_159 = proc_5_io_pipe_phv_out_data_159; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_160 = proc_5_io_pipe_phv_out_data_160; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_161 = proc_5_io_pipe_phv_out_data_161; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_162 = proc_5_io_pipe_phv_out_data_162; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_163 = proc_5_io_pipe_phv_out_data_163; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_164 = proc_5_io_pipe_phv_out_data_164; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_165 = proc_5_io_pipe_phv_out_data_165; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_166 = proc_5_io_pipe_phv_out_data_166; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_167 = proc_5_io_pipe_phv_out_data_167; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_168 = proc_5_io_pipe_phv_out_data_168; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_169 = proc_5_io_pipe_phv_out_data_169; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_170 = proc_5_io_pipe_phv_out_data_170; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_171 = proc_5_io_pipe_phv_out_data_171; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_172 = proc_5_io_pipe_phv_out_data_172; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_173 = proc_5_io_pipe_phv_out_data_173; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_174 = proc_5_io_pipe_phv_out_data_174; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_175 = proc_5_io_pipe_phv_out_data_175; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_176 = proc_5_io_pipe_phv_out_data_176; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_177 = proc_5_io_pipe_phv_out_data_177; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_178 = proc_5_io_pipe_phv_out_data_178; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_179 = proc_5_io_pipe_phv_out_data_179; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_180 = proc_5_io_pipe_phv_out_data_180; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_181 = proc_5_io_pipe_phv_out_data_181; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_182 = proc_5_io_pipe_phv_out_data_182; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_183 = proc_5_io_pipe_phv_out_data_183; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_184 = proc_5_io_pipe_phv_out_data_184; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_185 = proc_5_io_pipe_phv_out_data_185; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_186 = proc_5_io_pipe_phv_out_data_186; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_187 = proc_5_io_pipe_phv_out_data_187; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_188 = proc_5_io_pipe_phv_out_data_188; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_189 = proc_5_io_pipe_phv_out_data_189; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_190 = proc_5_io_pipe_phv_out_data_190; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_191 = proc_5_io_pipe_phv_out_data_191; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_192 = proc_5_io_pipe_phv_out_data_192; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_193 = proc_5_io_pipe_phv_out_data_193; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_194 = proc_5_io_pipe_phv_out_data_194; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_195 = proc_5_io_pipe_phv_out_data_195; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_196 = proc_5_io_pipe_phv_out_data_196; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_197 = proc_5_io_pipe_phv_out_data_197; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_198 = proc_5_io_pipe_phv_out_data_198; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_199 = proc_5_io_pipe_phv_out_data_199; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_200 = proc_5_io_pipe_phv_out_data_200; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_201 = proc_5_io_pipe_phv_out_data_201; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_202 = proc_5_io_pipe_phv_out_data_202; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_203 = proc_5_io_pipe_phv_out_data_203; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_204 = proc_5_io_pipe_phv_out_data_204; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_205 = proc_5_io_pipe_phv_out_data_205; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_206 = proc_5_io_pipe_phv_out_data_206; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_207 = proc_5_io_pipe_phv_out_data_207; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_208 = proc_5_io_pipe_phv_out_data_208; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_209 = proc_5_io_pipe_phv_out_data_209; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_210 = proc_5_io_pipe_phv_out_data_210; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_211 = proc_5_io_pipe_phv_out_data_211; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_212 = proc_5_io_pipe_phv_out_data_212; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_213 = proc_5_io_pipe_phv_out_data_213; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_214 = proc_5_io_pipe_phv_out_data_214; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_215 = proc_5_io_pipe_phv_out_data_215; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_216 = proc_5_io_pipe_phv_out_data_216; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_217 = proc_5_io_pipe_phv_out_data_217; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_218 = proc_5_io_pipe_phv_out_data_218; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_219 = proc_5_io_pipe_phv_out_data_219; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_220 = proc_5_io_pipe_phv_out_data_220; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_221 = proc_5_io_pipe_phv_out_data_221; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_222 = proc_5_io_pipe_phv_out_data_222; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_223 = proc_5_io_pipe_phv_out_data_223; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_224 = proc_5_io_pipe_phv_out_data_224; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_225 = proc_5_io_pipe_phv_out_data_225; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_226 = proc_5_io_pipe_phv_out_data_226; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_227 = proc_5_io_pipe_phv_out_data_227; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_228 = proc_5_io_pipe_phv_out_data_228; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_229 = proc_5_io_pipe_phv_out_data_229; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_230 = proc_5_io_pipe_phv_out_data_230; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_231 = proc_5_io_pipe_phv_out_data_231; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_232 = proc_5_io_pipe_phv_out_data_232; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_233 = proc_5_io_pipe_phv_out_data_233; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_234 = proc_5_io_pipe_phv_out_data_234; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_235 = proc_5_io_pipe_phv_out_data_235; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_236 = proc_5_io_pipe_phv_out_data_236; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_237 = proc_5_io_pipe_phv_out_data_237; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_238 = proc_5_io_pipe_phv_out_data_238; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_239 = proc_5_io_pipe_phv_out_data_239; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_240 = proc_5_io_pipe_phv_out_data_240; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_241 = proc_5_io_pipe_phv_out_data_241; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_242 = proc_5_io_pipe_phv_out_data_242; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_243 = proc_5_io_pipe_phv_out_data_243; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_244 = proc_5_io_pipe_phv_out_data_244; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_245 = proc_5_io_pipe_phv_out_data_245; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_246 = proc_5_io_pipe_phv_out_data_246; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_247 = proc_5_io_pipe_phv_out_data_247; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_248 = proc_5_io_pipe_phv_out_data_248; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_249 = proc_5_io_pipe_phv_out_data_249; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_250 = proc_5_io_pipe_phv_out_data_250; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_251 = proc_5_io_pipe_phv_out_data_251; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_252 = proc_5_io_pipe_phv_out_data_252; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_253 = proc_5_io_pipe_phv_out_data_253; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_254 = proc_5_io_pipe_phv_out_data_254; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_255 = proc_5_io_pipe_phv_out_data_255; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_next_processor_id = proc_5_io_pipe_phv_out_next_processor_id; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_next_config_id = proc_5_io_pipe_phv_out_next_config_id; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_is_valid_processor = 4'h6 == proc_5_io_pipe_phv_out_next_processor_id; // @[pisa.scala 36:62]
  assign proc_6_io_mod_mat_mod_en = io_mod_proc_mod_6_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_config_id = io_mod_proc_mod_6_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_6_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_6_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_6_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_6_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_6_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_6_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_6_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_6_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_6_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_6_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_6_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_6_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_6_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_w_en = io_mod_proc_mod_6_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_6_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_w_addr = io_mod_proc_mod_6_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_w_data = io_mod_proc_mod_6_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_6_io_mod_exe_mod_en_0 = io_mod_proc_mod_6_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_6_io_mod_exe_mod_en_1 = io_mod_proc_mod_6_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_6_io_mod_exe_mod_addr = io_mod_proc_mod_6_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_6_io_mod_exe_mod_data_0 = io_mod_proc_mod_6_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_6_io_mod_exe_mod_data_1 = io_mod_proc_mod_6_exe_mod_data_1; // @[pisa.scala 29:20]
  assign proc_7_clock = clock;
  assign proc_7_io_pipe_phv_in_data_0 = proc_6_io_pipe_phv_out_data_0; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_1 = proc_6_io_pipe_phv_out_data_1; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_2 = proc_6_io_pipe_phv_out_data_2; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_3 = proc_6_io_pipe_phv_out_data_3; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_4 = proc_6_io_pipe_phv_out_data_4; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_5 = proc_6_io_pipe_phv_out_data_5; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_6 = proc_6_io_pipe_phv_out_data_6; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_7 = proc_6_io_pipe_phv_out_data_7; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_8 = proc_6_io_pipe_phv_out_data_8; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_9 = proc_6_io_pipe_phv_out_data_9; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_10 = proc_6_io_pipe_phv_out_data_10; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_11 = proc_6_io_pipe_phv_out_data_11; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_12 = proc_6_io_pipe_phv_out_data_12; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_13 = proc_6_io_pipe_phv_out_data_13; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_14 = proc_6_io_pipe_phv_out_data_14; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_15 = proc_6_io_pipe_phv_out_data_15; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_16 = proc_6_io_pipe_phv_out_data_16; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_17 = proc_6_io_pipe_phv_out_data_17; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_18 = proc_6_io_pipe_phv_out_data_18; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_19 = proc_6_io_pipe_phv_out_data_19; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_20 = proc_6_io_pipe_phv_out_data_20; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_21 = proc_6_io_pipe_phv_out_data_21; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_22 = proc_6_io_pipe_phv_out_data_22; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_23 = proc_6_io_pipe_phv_out_data_23; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_24 = proc_6_io_pipe_phv_out_data_24; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_25 = proc_6_io_pipe_phv_out_data_25; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_26 = proc_6_io_pipe_phv_out_data_26; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_27 = proc_6_io_pipe_phv_out_data_27; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_28 = proc_6_io_pipe_phv_out_data_28; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_29 = proc_6_io_pipe_phv_out_data_29; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_30 = proc_6_io_pipe_phv_out_data_30; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_31 = proc_6_io_pipe_phv_out_data_31; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_32 = proc_6_io_pipe_phv_out_data_32; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_33 = proc_6_io_pipe_phv_out_data_33; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_34 = proc_6_io_pipe_phv_out_data_34; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_35 = proc_6_io_pipe_phv_out_data_35; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_36 = proc_6_io_pipe_phv_out_data_36; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_37 = proc_6_io_pipe_phv_out_data_37; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_38 = proc_6_io_pipe_phv_out_data_38; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_39 = proc_6_io_pipe_phv_out_data_39; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_40 = proc_6_io_pipe_phv_out_data_40; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_41 = proc_6_io_pipe_phv_out_data_41; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_42 = proc_6_io_pipe_phv_out_data_42; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_43 = proc_6_io_pipe_phv_out_data_43; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_44 = proc_6_io_pipe_phv_out_data_44; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_45 = proc_6_io_pipe_phv_out_data_45; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_46 = proc_6_io_pipe_phv_out_data_46; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_47 = proc_6_io_pipe_phv_out_data_47; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_48 = proc_6_io_pipe_phv_out_data_48; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_49 = proc_6_io_pipe_phv_out_data_49; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_50 = proc_6_io_pipe_phv_out_data_50; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_51 = proc_6_io_pipe_phv_out_data_51; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_52 = proc_6_io_pipe_phv_out_data_52; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_53 = proc_6_io_pipe_phv_out_data_53; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_54 = proc_6_io_pipe_phv_out_data_54; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_55 = proc_6_io_pipe_phv_out_data_55; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_56 = proc_6_io_pipe_phv_out_data_56; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_57 = proc_6_io_pipe_phv_out_data_57; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_58 = proc_6_io_pipe_phv_out_data_58; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_59 = proc_6_io_pipe_phv_out_data_59; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_60 = proc_6_io_pipe_phv_out_data_60; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_61 = proc_6_io_pipe_phv_out_data_61; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_62 = proc_6_io_pipe_phv_out_data_62; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_63 = proc_6_io_pipe_phv_out_data_63; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_64 = proc_6_io_pipe_phv_out_data_64; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_65 = proc_6_io_pipe_phv_out_data_65; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_66 = proc_6_io_pipe_phv_out_data_66; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_67 = proc_6_io_pipe_phv_out_data_67; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_68 = proc_6_io_pipe_phv_out_data_68; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_69 = proc_6_io_pipe_phv_out_data_69; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_70 = proc_6_io_pipe_phv_out_data_70; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_71 = proc_6_io_pipe_phv_out_data_71; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_72 = proc_6_io_pipe_phv_out_data_72; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_73 = proc_6_io_pipe_phv_out_data_73; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_74 = proc_6_io_pipe_phv_out_data_74; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_75 = proc_6_io_pipe_phv_out_data_75; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_76 = proc_6_io_pipe_phv_out_data_76; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_77 = proc_6_io_pipe_phv_out_data_77; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_78 = proc_6_io_pipe_phv_out_data_78; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_79 = proc_6_io_pipe_phv_out_data_79; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_80 = proc_6_io_pipe_phv_out_data_80; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_81 = proc_6_io_pipe_phv_out_data_81; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_82 = proc_6_io_pipe_phv_out_data_82; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_83 = proc_6_io_pipe_phv_out_data_83; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_84 = proc_6_io_pipe_phv_out_data_84; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_85 = proc_6_io_pipe_phv_out_data_85; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_86 = proc_6_io_pipe_phv_out_data_86; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_87 = proc_6_io_pipe_phv_out_data_87; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_88 = proc_6_io_pipe_phv_out_data_88; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_89 = proc_6_io_pipe_phv_out_data_89; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_90 = proc_6_io_pipe_phv_out_data_90; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_91 = proc_6_io_pipe_phv_out_data_91; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_92 = proc_6_io_pipe_phv_out_data_92; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_93 = proc_6_io_pipe_phv_out_data_93; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_94 = proc_6_io_pipe_phv_out_data_94; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_95 = proc_6_io_pipe_phv_out_data_95; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_96 = proc_6_io_pipe_phv_out_data_96; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_97 = proc_6_io_pipe_phv_out_data_97; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_98 = proc_6_io_pipe_phv_out_data_98; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_99 = proc_6_io_pipe_phv_out_data_99; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_100 = proc_6_io_pipe_phv_out_data_100; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_101 = proc_6_io_pipe_phv_out_data_101; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_102 = proc_6_io_pipe_phv_out_data_102; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_103 = proc_6_io_pipe_phv_out_data_103; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_104 = proc_6_io_pipe_phv_out_data_104; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_105 = proc_6_io_pipe_phv_out_data_105; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_106 = proc_6_io_pipe_phv_out_data_106; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_107 = proc_6_io_pipe_phv_out_data_107; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_108 = proc_6_io_pipe_phv_out_data_108; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_109 = proc_6_io_pipe_phv_out_data_109; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_110 = proc_6_io_pipe_phv_out_data_110; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_111 = proc_6_io_pipe_phv_out_data_111; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_112 = proc_6_io_pipe_phv_out_data_112; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_113 = proc_6_io_pipe_phv_out_data_113; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_114 = proc_6_io_pipe_phv_out_data_114; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_115 = proc_6_io_pipe_phv_out_data_115; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_116 = proc_6_io_pipe_phv_out_data_116; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_117 = proc_6_io_pipe_phv_out_data_117; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_118 = proc_6_io_pipe_phv_out_data_118; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_119 = proc_6_io_pipe_phv_out_data_119; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_120 = proc_6_io_pipe_phv_out_data_120; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_121 = proc_6_io_pipe_phv_out_data_121; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_122 = proc_6_io_pipe_phv_out_data_122; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_123 = proc_6_io_pipe_phv_out_data_123; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_124 = proc_6_io_pipe_phv_out_data_124; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_125 = proc_6_io_pipe_phv_out_data_125; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_126 = proc_6_io_pipe_phv_out_data_126; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_127 = proc_6_io_pipe_phv_out_data_127; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_128 = proc_6_io_pipe_phv_out_data_128; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_129 = proc_6_io_pipe_phv_out_data_129; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_130 = proc_6_io_pipe_phv_out_data_130; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_131 = proc_6_io_pipe_phv_out_data_131; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_132 = proc_6_io_pipe_phv_out_data_132; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_133 = proc_6_io_pipe_phv_out_data_133; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_134 = proc_6_io_pipe_phv_out_data_134; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_135 = proc_6_io_pipe_phv_out_data_135; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_136 = proc_6_io_pipe_phv_out_data_136; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_137 = proc_6_io_pipe_phv_out_data_137; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_138 = proc_6_io_pipe_phv_out_data_138; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_139 = proc_6_io_pipe_phv_out_data_139; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_140 = proc_6_io_pipe_phv_out_data_140; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_141 = proc_6_io_pipe_phv_out_data_141; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_142 = proc_6_io_pipe_phv_out_data_142; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_143 = proc_6_io_pipe_phv_out_data_143; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_144 = proc_6_io_pipe_phv_out_data_144; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_145 = proc_6_io_pipe_phv_out_data_145; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_146 = proc_6_io_pipe_phv_out_data_146; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_147 = proc_6_io_pipe_phv_out_data_147; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_148 = proc_6_io_pipe_phv_out_data_148; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_149 = proc_6_io_pipe_phv_out_data_149; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_150 = proc_6_io_pipe_phv_out_data_150; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_151 = proc_6_io_pipe_phv_out_data_151; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_152 = proc_6_io_pipe_phv_out_data_152; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_153 = proc_6_io_pipe_phv_out_data_153; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_154 = proc_6_io_pipe_phv_out_data_154; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_155 = proc_6_io_pipe_phv_out_data_155; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_156 = proc_6_io_pipe_phv_out_data_156; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_157 = proc_6_io_pipe_phv_out_data_157; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_158 = proc_6_io_pipe_phv_out_data_158; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_159 = proc_6_io_pipe_phv_out_data_159; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_160 = proc_6_io_pipe_phv_out_data_160; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_161 = proc_6_io_pipe_phv_out_data_161; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_162 = proc_6_io_pipe_phv_out_data_162; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_163 = proc_6_io_pipe_phv_out_data_163; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_164 = proc_6_io_pipe_phv_out_data_164; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_165 = proc_6_io_pipe_phv_out_data_165; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_166 = proc_6_io_pipe_phv_out_data_166; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_167 = proc_6_io_pipe_phv_out_data_167; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_168 = proc_6_io_pipe_phv_out_data_168; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_169 = proc_6_io_pipe_phv_out_data_169; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_170 = proc_6_io_pipe_phv_out_data_170; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_171 = proc_6_io_pipe_phv_out_data_171; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_172 = proc_6_io_pipe_phv_out_data_172; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_173 = proc_6_io_pipe_phv_out_data_173; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_174 = proc_6_io_pipe_phv_out_data_174; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_175 = proc_6_io_pipe_phv_out_data_175; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_176 = proc_6_io_pipe_phv_out_data_176; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_177 = proc_6_io_pipe_phv_out_data_177; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_178 = proc_6_io_pipe_phv_out_data_178; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_179 = proc_6_io_pipe_phv_out_data_179; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_180 = proc_6_io_pipe_phv_out_data_180; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_181 = proc_6_io_pipe_phv_out_data_181; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_182 = proc_6_io_pipe_phv_out_data_182; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_183 = proc_6_io_pipe_phv_out_data_183; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_184 = proc_6_io_pipe_phv_out_data_184; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_185 = proc_6_io_pipe_phv_out_data_185; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_186 = proc_6_io_pipe_phv_out_data_186; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_187 = proc_6_io_pipe_phv_out_data_187; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_188 = proc_6_io_pipe_phv_out_data_188; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_189 = proc_6_io_pipe_phv_out_data_189; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_190 = proc_6_io_pipe_phv_out_data_190; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_191 = proc_6_io_pipe_phv_out_data_191; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_192 = proc_6_io_pipe_phv_out_data_192; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_193 = proc_6_io_pipe_phv_out_data_193; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_194 = proc_6_io_pipe_phv_out_data_194; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_195 = proc_6_io_pipe_phv_out_data_195; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_196 = proc_6_io_pipe_phv_out_data_196; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_197 = proc_6_io_pipe_phv_out_data_197; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_198 = proc_6_io_pipe_phv_out_data_198; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_199 = proc_6_io_pipe_phv_out_data_199; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_200 = proc_6_io_pipe_phv_out_data_200; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_201 = proc_6_io_pipe_phv_out_data_201; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_202 = proc_6_io_pipe_phv_out_data_202; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_203 = proc_6_io_pipe_phv_out_data_203; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_204 = proc_6_io_pipe_phv_out_data_204; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_205 = proc_6_io_pipe_phv_out_data_205; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_206 = proc_6_io_pipe_phv_out_data_206; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_207 = proc_6_io_pipe_phv_out_data_207; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_208 = proc_6_io_pipe_phv_out_data_208; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_209 = proc_6_io_pipe_phv_out_data_209; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_210 = proc_6_io_pipe_phv_out_data_210; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_211 = proc_6_io_pipe_phv_out_data_211; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_212 = proc_6_io_pipe_phv_out_data_212; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_213 = proc_6_io_pipe_phv_out_data_213; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_214 = proc_6_io_pipe_phv_out_data_214; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_215 = proc_6_io_pipe_phv_out_data_215; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_216 = proc_6_io_pipe_phv_out_data_216; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_217 = proc_6_io_pipe_phv_out_data_217; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_218 = proc_6_io_pipe_phv_out_data_218; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_219 = proc_6_io_pipe_phv_out_data_219; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_220 = proc_6_io_pipe_phv_out_data_220; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_221 = proc_6_io_pipe_phv_out_data_221; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_222 = proc_6_io_pipe_phv_out_data_222; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_223 = proc_6_io_pipe_phv_out_data_223; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_224 = proc_6_io_pipe_phv_out_data_224; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_225 = proc_6_io_pipe_phv_out_data_225; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_226 = proc_6_io_pipe_phv_out_data_226; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_227 = proc_6_io_pipe_phv_out_data_227; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_228 = proc_6_io_pipe_phv_out_data_228; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_229 = proc_6_io_pipe_phv_out_data_229; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_230 = proc_6_io_pipe_phv_out_data_230; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_231 = proc_6_io_pipe_phv_out_data_231; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_232 = proc_6_io_pipe_phv_out_data_232; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_233 = proc_6_io_pipe_phv_out_data_233; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_234 = proc_6_io_pipe_phv_out_data_234; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_235 = proc_6_io_pipe_phv_out_data_235; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_236 = proc_6_io_pipe_phv_out_data_236; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_237 = proc_6_io_pipe_phv_out_data_237; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_238 = proc_6_io_pipe_phv_out_data_238; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_239 = proc_6_io_pipe_phv_out_data_239; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_240 = proc_6_io_pipe_phv_out_data_240; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_241 = proc_6_io_pipe_phv_out_data_241; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_242 = proc_6_io_pipe_phv_out_data_242; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_243 = proc_6_io_pipe_phv_out_data_243; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_244 = proc_6_io_pipe_phv_out_data_244; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_245 = proc_6_io_pipe_phv_out_data_245; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_246 = proc_6_io_pipe_phv_out_data_246; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_247 = proc_6_io_pipe_phv_out_data_247; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_248 = proc_6_io_pipe_phv_out_data_248; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_249 = proc_6_io_pipe_phv_out_data_249; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_250 = proc_6_io_pipe_phv_out_data_250; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_251 = proc_6_io_pipe_phv_out_data_251; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_252 = proc_6_io_pipe_phv_out_data_252; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_253 = proc_6_io_pipe_phv_out_data_253; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_254 = proc_6_io_pipe_phv_out_data_254; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_255 = proc_6_io_pipe_phv_out_data_255; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_next_processor_id = proc_6_io_pipe_phv_out_next_processor_id; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_next_config_id = proc_6_io_pipe_phv_out_next_config_id; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_is_valid_processor = 4'h7 == proc_6_io_pipe_phv_out_next_processor_id; // @[pisa.scala 36:62]
  assign proc_7_io_mod_mat_mod_en = io_mod_proc_mod_7_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_config_id = io_mod_proc_mod_7_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_7_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_7_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_7_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_7_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_7_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_7_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_7_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_7_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_7_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_7_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_7_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_7_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_7_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_w_en = io_mod_proc_mod_7_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_7_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_w_addr = io_mod_proc_mod_7_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_w_data = io_mod_proc_mod_7_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_7_io_mod_exe_mod_en_0 = io_mod_proc_mod_7_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_7_io_mod_exe_mod_en_1 = io_mod_proc_mod_7_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_7_io_mod_exe_mod_addr = io_mod_proc_mod_7_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_7_io_mod_exe_mod_data_0 = io_mod_proc_mod_7_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_7_io_mod_exe_mod_data_1 = io_mod_proc_mod_7_exe_mod_data_1; // @[pisa.scala 29:20]
  assign proc_8_clock = clock;
  assign proc_8_io_pipe_phv_in_data_0 = proc_7_io_pipe_phv_out_data_0; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_1 = proc_7_io_pipe_phv_out_data_1; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_2 = proc_7_io_pipe_phv_out_data_2; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_3 = proc_7_io_pipe_phv_out_data_3; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_4 = proc_7_io_pipe_phv_out_data_4; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_5 = proc_7_io_pipe_phv_out_data_5; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_6 = proc_7_io_pipe_phv_out_data_6; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_7 = proc_7_io_pipe_phv_out_data_7; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_8 = proc_7_io_pipe_phv_out_data_8; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_9 = proc_7_io_pipe_phv_out_data_9; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_10 = proc_7_io_pipe_phv_out_data_10; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_11 = proc_7_io_pipe_phv_out_data_11; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_12 = proc_7_io_pipe_phv_out_data_12; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_13 = proc_7_io_pipe_phv_out_data_13; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_14 = proc_7_io_pipe_phv_out_data_14; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_15 = proc_7_io_pipe_phv_out_data_15; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_16 = proc_7_io_pipe_phv_out_data_16; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_17 = proc_7_io_pipe_phv_out_data_17; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_18 = proc_7_io_pipe_phv_out_data_18; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_19 = proc_7_io_pipe_phv_out_data_19; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_20 = proc_7_io_pipe_phv_out_data_20; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_21 = proc_7_io_pipe_phv_out_data_21; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_22 = proc_7_io_pipe_phv_out_data_22; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_23 = proc_7_io_pipe_phv_out_data_23; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_24 = proc_7_io_pipe_phv_out_data_24; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_25 = proc_7_io_pipe_phv_out_data_25; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_26 = proc_7_io_pipe_phv_out_data_26; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_27 = proc_7_io_pipe_phv_out_data_27; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_28 = proc_7_io_pipe_phv_out_data_28; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_29 = proc_7_io_pipe_phv_out_data_29; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_30 = proc_7_io_pipe_phv_out_data_30; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_31 = proc_7_io_pipe_phv_out_data_31; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_32 = proc_7_io_pipe_phv_out_data_32; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_33 = proc_7_io_pipe_phv_out_data_33; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_34 = proc_7_io_pipe_phv_out_data_34; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_35 = proc_7_io_pipe_phv_out_data_35; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_36 = proc_7_io_pipe_phv_out_data_36; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_37 = proc_7_io_pipe_phv_out_data_37; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_38 = proc_7_io_pipe_phv_out_data_38; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_39 = proc_7_io_pipe_phv_out_data_39; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_40 = proc_7_io_pipe_phv_out_data_40; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_41 = proc_7_io_pipe_phv_out_data_41; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_42 = proc_7_io_pipe_phv_out_data_42; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_43 = proc_7_io_pipe_phv_out_data_43; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_44 = proc_7_io_pipe_phv_out_data_44; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_45 = proc_7_io_pipe_phv_out_data_45; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_46 = proc_7_io_pipe_phv_out_data_46; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_47 = proc_7_io_pipe_phv_out_data_47; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_48 = proc_7_io_pipe_phv_out_data_48; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_49 = proc_7_io_pipe_phv_out_data_49; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_50 = proc_7_io_pipe_phv_out_data_50; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_51 = proc_7_io_pipe_phv_out_data_51; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_52 = proc_7_io_pipe_phv_out_data_52; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_53 = proc_7_io_pipe_phv_out_data_53; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_54 = proc_7_io_pipe_phv_out_data_54; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_55 = proc_7_io_pipe_phv_out_data_55; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_56 = proc_7_io_pipe_phv_out_data_56; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_57 = proc_7_io_pipe_phv_out_data_57; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_58 = proc_7_io_pipe_phv_out_data_58; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_59 = proc_7_io_pipe_phv_out_data_59; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_60 = proc_7_io_pipe_phv_out_data_60; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_61 = proc_7_io_pipe_phv_out_data_61; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_62 = proc_7_io_pipe_phv_out_data_62; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_63 = proc_7_io_pipe_phv_out_data_63; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_64 = proc_7_io_pipe_phv_out_data_64; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_65 = proc_7_io_pipe_phv_out_data_65; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_66 = proc_7_io_pipe_phv_out_data_66; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_67 = proc_7_io_pipe_phv_out_data_67; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_68 = proc_7_io_pipe_phv_out_data_68; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_69 = proc_7_io_pipe_phv_out_data_69; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_70 = proc_7_io_pipe_phv_out_data_70; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_71 = proc_7_io_pipe_phv_out_data_71; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_72 = proc_7_io_pipe_phv_out_data_72; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_73 = proc_7_io_pipe_phv_out_data_73; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_74 = proc_7_io_pipe_phv_out_data_74; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_75 = proc_7_io_pipe_phv_out_data_75; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_76 = proc_7_io_pipe_phv_out_data_76; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_77 = proc_7_io_pipe_phv_out_data_77; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_78 = proc_7_io_pipe_phv_out_data_78; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_79 = proc_7_io_pipe_phv_out_data_79; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_80 = proc_7_io_pipe_phv_out_data_80; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_81 = proc_7_io_pipe_phv_out_data_81; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_82 = proc_7_io_pipe_phv_out_data_82; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_83 = proc_7_io_pipe_phv_out_data_83; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_84 = proc_7_io_pipe_phv_out_data_84; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_85 = proc_7_io_pipe_phv_out_data_85; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_86 = proc_7_io_pipe_phv_out_data_86; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_87 = proc_7_io_pipe_phv_out_data_87; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_88 = proc_7_io_pipe_phv_out_data_88; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_89 = proc_7_io_pipe_phv_out_data_89; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_90 = proc_7_io_pipe_phv_out_data_90; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_91 = proc_7_io_pipe_phv_out_data_91; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_92 = proc_7_io_pipe_phv_out_data_92; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_93 = proc_7_io_pipe_phv_out_data_93; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_94 = proc_7_io_pipe_phv_out_data_94; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_95 = proc_7_io_pipe_phv_out_data_95; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_96 = proc_7_io_pipe_phv_out_data_96; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_97 = proc_7_io_pipe_phv_out_data_97; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_98 = proc_7_io_pipe_phv_out_data_98; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_99 = proc_7_io_pipe_phv_out_data_99; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_100 = proc_7_io_pipe_phv_out_data_100; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_101 = proc_7_io_pipe_phv_out_data_101; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_102 = proc_7_io_pipe_phv_out_data_102; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_103 = proc_7_io_pipe_phv_out_data_103; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_104 = proc_7_io_pipe_phv_out_data_104; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_105 = proc_7_io_pipe_phv_out_data_105; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_106 = proc_7_io_pipe_phv_out_data_106; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_107 = proc_7_io_pipe_phv_out_data_107; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_108 = proc_7_io_pipe_phv_out_data_108; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_109 = proc_7_io_pipe_phv_out_data_109; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_110 = proc_7_io_pipe_phv_out_data_110; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_111 = proc_7_io_pipe_phv_out_data_111; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_112 = proc_7_io_pipe_phv_out_data_112; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_113 = proc_7_io_pipe_phv_out_data_113; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_114 = proc_7_io_pipe_phv_out_data_114; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_115 = proc_7_io_pipe_phv_out_data_115; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_116 = proc_7_io_pipe_phv_out_data_116; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_117 = proc_7_io_pipe_phv_out_data_117; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_118 = proc_7_io_pipe_phv_out_data_118; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_119 = proc_7_io_pipe_phv_out_data_119; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_120 = proc_7_io_pipe_phv_out_data_120; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_121 = proc_7_io_pipe_phv_out_data_121; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_122 = proc_7_io_pipe_phv_out_data_122; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_123 = proc_7_io_pipe_phv_out_data_123; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_124 = proc_7_io_pipe_phv_out_data_124; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_125 = proc_7_io_pipe_phv_out_data_125; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_126 = proc_7_io_pipe_phv_out_data_126; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_127 = proc_7_io_pipe_phv_out_data_127; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_128 = proc_7_io_pipe_phv_out_data_128; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_129 = proc_7_io_pipe_phv_out_data_129; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_130 = proc_7_io_pipe_phv_out_data_130; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_131 = proc_7_io_pipe_phv_out_data_131; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_132 = proc_7_io_pipe_phv_out_data_132; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_133 = proc_7_io_pipe_phv_out_data_133; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_134 = proc_7_io_pipe_phv_out_data_134; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_135 = proc_7_io_pipe_phv_out_data_135; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_136 = proc_7_io_pipe_phv_out_data_136; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_137 = proc_7_io_pipe_phv_out_data_137; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_138 = proc_7_io_pipe_phv_out_data_138; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_139 = proc_7_io_pipe_phv_out_data_139; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_140 = proc_7_io_pipe_phv_out_data_140; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_141 = proc_7_io_pipe_phv_out_data_141; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_142 = proc_7_io_pipe_phv_out_data_142; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_143 = proc_7_io_pipe_phv_out_data_143; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_144 = proc_7_io_pipe_phv_out_data_144; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_145 = proc_7_io_pipe_phv_out_data_145; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_146 = proc_7_io_pipe_phv_out_data_146; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_147 = proc_7_io_pipe_phv_out_data_147; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_148 = proc_7_io_pipe_phv_out_data_148; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_149 = proc_7_io_pipe_phv_out_data_149; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_150 = proc_7_io_pipe_phv_out_data_150; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_151 = proc_7_io_pipe_phv_out_data_151; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_152 = proc_7_io_pipe_phv_out_data_152; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_153 = proc_7_io_pipe_phv_out_data_153; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_154 = proc_7_io_pipe_phv_out_data_154; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_155 = proc_7_io_pipe_phv_out_data_155; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_156 = proc_7_io_pipe_phv_out_data_156; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_157 = proc_7_io_pipe_phv_out_data_157; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_158 = proc_7_io_pipe_phv_out_data_158; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_159 = proc_7_io_pipe_phv_out_data_159; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_160 = proc_7_io_pipe_phv_out_data_160; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_161 = proc_7_io_pipe_phv_out_data_161; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_162 = proc_7_io_pipe_phv_out_data_162; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_163 = proc_7_io_pipe_phv_out_data_163; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_164 = proc_7_io_pipe_phv_out_data_164; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_165 = proc_7_io_pipe_phv_out_data_165; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_166 = proc_7_io_pipe_phv_out_data_166; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_167 = proc_7_io_pipe_phv_out_data_167; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_168 = proc_7_io_pipe_phv_out_data_168; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_169 = proc_7_io_pipe_phv_out_data_169; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_170 = proc_7_io_pipe_phv_out_data_170; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_171 = proc_7_io_pipe_phv_out_data_171; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_172 = proc_7_io_pipe_phv_out_data_172; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_173 = proc_7_io_pipe_phv_out_data_173; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_174 = proc_7_io_pipe_phv_out_data_174; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_175 = proc_7_io_pipe_phv_out_data_175; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_176 = proc_7_io_pipe_phv_out_data_176; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_177 = proc_7_io_pipe_phv_out_data_177; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_178 = proc_7_io_pipe_phv_out_data_178; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_179 = proc_7_io_pipe_phv_out_data_179; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_180 = proc_7_io_pipe_phv_out_data_180; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_181 = proc_7_io_pipe_phv_out_data_181; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_182 = proc_7_io_pipe_phv_out_data_182; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_183 = proc_7_io_pipe_phv_out_data_183; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_184 = proc_7_io_pipe_phv_out_data_184; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_185 = proc_7_io_pipe_phv_out_data_185; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_186 = proc_7_io_pipe_phv_out_data_186; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_187 = proc_7_io_pipe_phv_out_data_187; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_188 = proc_7_io_pipe_phv_out_data_188; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_189 = proc_7_io_pipe_phv_out_data_189; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_190 = proc_7_io_pipe_phv_out_data_190; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_191 = proc_7_io_pipe_phv_out_data_191; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_192 = proc_7_io_pipe_phv_out_data_192; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_193 = proc_7_io_pipe_phv_out_data_193; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_194 = proc_7_io_pipe_phv_out_data_194; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_195 = proc_7_io_pipe_phv_out_data_195; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_196 = proc_7_io_pipe_phv_out_data_196; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_197 = proc_7_io_pipe_phv_out_data_197; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_198 = proc_7_io_pipe_phv_out_data_198; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_199 = proc_7_io_pipe_phv_out_data_199; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_200 = proc_7_io_pipe_phv_out_data_200; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_201 = proc_7_io_pipe_phv_out_data_201; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_202 = proc_7_io_pipe_phv_out_data_202; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_203 = proc_7_io_pipe_phv_out_data_203; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_204 = proc_7_io_pipe_phv_out_data_204; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_205 = proc_7_io_pipe_phv_out_data_205; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_206 = proc_7_io_pipe_phv_out_data_206; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_207 = proc_7_io_pipe_phv_out_data_207; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_208 = proc_7_io_pipe_phv_out_data_208; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_209 = proc_7_io_pipe_phv_out_data_209; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_210 = proc_7_io_pipe_phv_out_data_210; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_211 = proc_7_io_pipe_phv_out_data_211; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_212 = proc_7_io_pipe_phv_out_data_212; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_213 = proc_7_io_pipe_phv_out_data_213; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_214 = proc_7_io_pipe_phv_out_data_214; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_215 = proc_7_io_pipe_phv_out_data_215; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_216 = proc_7_io_pipe_phv_out_data_216; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_217 = proc_7_io_pipe_phv_out_data_217; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_218 = proc_7_io_pipe_phv_out_data_218; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_219 = proc_7_io_pipe_phv_out_data_219; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_220 = proc_7_io_pipe_phv_out_data_220; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_221 = proc_7_io_pipe_phv_out_data_221; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_222 = proc_7_io_pipe_phv_out_data_222; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_223 = proc_7_io_pipe_phv_out_data_223; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_224 = proc_7_io_pipe_phv_out_data_224; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_225 = proc_7_io_pipe_phv_out_data_225; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_226 = proc_7_io_pipe_phv_out_data_226; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_227 = proc_7_io_pipe_phv_out_data_227; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_228 = proc_7_io_pipe_phv_out_data_228; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_229 = proc_7_io_pipe_phv_out_data_229; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_230 = proc_7_io_pipe_phv_out_data_230; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_231 = proc_7_io_pipe_phv_out_data_231; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_232 = proc_7_io_pipe_phv_out_data_232; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_233 = proc_7_io_pipe_phv_out_data_233; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_234 = proc_7_io_pipe_phv_out_data_234; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_235 = proc_7_io_pipe_phv_out_data_235; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_236 = proc_7_io_pipe_phv_out_data_236; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_237 = proc_7_io_pipe_phv_out_data_237; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_238 = proc_7_io_pipe_phv_out_data_238; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_239 = proc_7_io_pipe_phv_out_data_239; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_240 = proc_7_io_pipe_phv_out_data_240; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_241 = proc_7_io_pipe_phv_out_data_241; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_242 = proc_7_io_pipe_phv_out_data_242; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_243 = proc_7_io_pipe_phv_out_data_243; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_244 = proc_7_io_pipe_phv_out_data_244; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_245 = proc_7_io_pipe_phv_out_data_245; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_246 = proc_7_io_pipe_phv_out_data_246; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_247 = proc_7_io_pipe_phv_out_data_247; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_248 = proc_7_io_pipe_phv_out_data_248; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_249 = proc_7_io_pipe_phv_out_data_249; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_250 = proc_7_io_pipe_phv_out_data_250; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_251 = proc_7_io_pipe_phv_out_data_251; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_252 = proc_7_io_pipe_phv_out_data_252; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_253 = proc_7_io_pipe_phv_out_data_253; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_254 = proc_7_io_pipe_phv_out_data_254; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_255 = proc_7_io_pipe_phv_out_data_255; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_next_processor_id = proc_7_io_pipe_phv_out_next_processor_id; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_next_config_id = proc_7_io_pipe_phv_out_next_config_id; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_is_valid_processor = 4'h8 == proc_7_io_pipe_phv_out_next_processor_id; // @[pisa.scala 36:62]
  assign proc_8_io_mod_mat_mod_en = io_mod_proc_mod_8_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_config_id = io_mod_proc_mod_8_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_8_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_8_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_8_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_8_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_8_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_8_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_8_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_8_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_8_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_8_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_8_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_8_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_8_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_w_en = io_mod_proc_mod_8_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_8_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_w_addr = io_mod_proc_mod_8_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_w_data = io_mod_proc_mod_8_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_8_io_mod_exe_mod_en_0 = io_mod_proc_mod_8_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_8_io_mod_exe_mod_en_1 = io_mod_proc_mod_8_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_8_io_mod_exe_mod_addr = io_mod_proc_mod_8_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_8_io_mod_exe_mod_data_0 = io_mod_proc_mod_8_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_8_io_mod_exe_mod_data_1 = io_mod_proc_mod_8_exe_mod_data_1; // @[pisa.scala 29:20]
  assign proc_9_clock = clock;
  assign proc_9_io_pipe_phv_in_data_0 = proc_8_io_pipe_phv_out_data_0; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_1 = proc_8_io_pipe_phv_out_data_1; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_2 = proc_8_io_pipe_phv_out_data_2; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_3 = proc_8_io_pipe_phv_out_data_3; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_4 = proc_8_io_pipe_phv_out_data_4; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_5 = proc_8_io_pipe_phv_out_data_5; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_6 = proc_8_io_pipe_phv_out_data_6; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_7 = proc_8_io_pipe_phv_out_data_7; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_8 = proc_8_io_pipe_phv_out_data_8; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_9 = proc_8_io_pipe_phv_out_data_9; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_10 = proc_8_io_pipe_phv_out_data_10; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_11 = proc_8_io_pipe_phv_out_data_11; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_12 = proc_8_io_pipe_phv_out_data_12; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_13 = proc_8_io_pipe_phv_out_data_13; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_14 = proc_8_io_pipe_phv_out_data_14; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_15 = proc_8_io_pipe_phv_out_data_15; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_16 = proc_8_io_pipe_phv_out_data_16; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_17 = proc_8_io_pipe_phv_out_data_17; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_18 = proc_8_io_pipe_phv_out_data_18; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_19 = proc_8_io_pipe_phv_out_data_19; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_20 = proc_8_io_pipe_phv_out_data_20; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_21 = proc_8_io_pipe_phv_out_data_21; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_22 = proc_8_io_pipe_phv_out_data_22; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_23 = proc_8_io_pipe_phv_out_data_23; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_24 = proc_8_io_pipe_phv_out_data_24; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_25 = proc_8_io_pipe_phv_out_data_25; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_26 = proc_8_io_pipe_phv_out_data_26; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_27 = proc_8_io_pipe_phv_out_data_27; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_28 = proc_8_io_pipe_phv_out_data_28; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_29 = proc_8_io_pipe_phv_out_data_29; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_30 = proc_8_io_pipe_phv_out_data_30; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_31 = proc_8_io_pipe_phv_out_data_31; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_32 = proc_8_io_pipe_phv_out_data_32; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_33 = proc_8_io_pipe_phv_out_data_33; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_34 = proc_8_io_pipe_phv_out_data_34; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_35 = proc_8_io_pipe_phv_out_data_35; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_36 = proc_8_io_pipe_phv_out_data_36; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_37 = proc_8_io_pipe_phv_out_data_37; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_38 = proc_8_io_pipe_phv_out_data_38; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_39 = proc_8_io_pipe_phv_out_data_39; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_40 = proc_8_io_pipe_phv_out_data_40; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_41 = proc_8_io_pipe_phv_out_data_41; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_42 = proc_8_io_pipe_phv_out_data_42; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_43 = proc_8_io_pipe_phv_out_data_43; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_44 = proc_8_io_pipe_phv_out_data_44; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_45 = proc_8_io_pipe_phv_out_data_45; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_46 = proc_8_io_pipe_phv_out_data_46; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_47 = proc_8_io_pipe_phv_out_data_47; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_48 = proc_8_io_pipe_phv_out_data_48; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_49 = proc_8_io_pipe_phv_out_data_49; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_50 = proc_8_io_pipe_phv_out_data_50; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_51 = proc_8_io_pipe_phv_out_data_51; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_52 = proc_8_io_pipe_phv_out_data_52; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_53 = proc_8_io_pipe_phv_out_data_53; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_54 = proc_8_io_pipe_phv_out_data_54; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_55 = proc_8_io_pipe_phv_out_data_55; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_56 = proc_8_io_pipe_phv_out_data_56; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_57 = proc_8_io_pipe_phv_out_data_57; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_58 = proc_8_io_pipe_phv_out_data_58; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_59 = proc_8_io_pipe_phv_out_data_59; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_60 = proc_8_io_pipe_phv_out_data_60; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_61 = proc_8_io_pipe_phv_out_data_61; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_62 = proc_8_io_pipe_phv_out_data_62; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_63 = proc_8_io_pipe_phv_out_data_63; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_64 = proc_8_io_pipe_phv_out_data_64; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_65 = proc_8_io_pipe_phv_out_data_65; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_66 = proc_8_io_pipe_phv_out_data_66; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_67 = proc_8_io_pipe_phv_out_data_67; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_68 = proc_8_io_pipe_phv_out_data_68; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_69 = proc_8_io_pipe_phv_out_data_69; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_70 = proc_8_io_pipe_phv_out_data_70; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_71 = proc_8_io_pipe_phv_out_data_71; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_72 = proc_8_io_pipe_phv_out_data_72; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_73 = proc_8_io_pipe_phv_out_data_73; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_74 = proc_8_io_pipe_phv_out_data_74; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_75 = proc_8_io_pipe_phv_out_data_75; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_76 = proc_8_io_pipe_phv_out_data_76; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_77 = proc_8_io_pipe_phv_out_data_77; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_78 = proc_8_io_pipe_phv_out_data_78; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_79 = proc_8_io_pipe_phv_out_data_79; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_80 = proc_8_io_pipe_phv_out_data_80; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_81 = proc_8_io_pipe_phv_out_data_81; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_82 = proc_8_io_pipe_phv_out_data_82; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_83 = proc_8_io_pipe_phv_out_data_83; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_84 = proc_8_io_pipe_phv_out_data_84; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_85 = proc_8_io_pipe_phv_out_data_85; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_86 = proc_8_io_pipe_phv_out_data_86; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_87 = proc_8_io_pipe_phv_out_data_87; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_88 = proc_8_io_pipe_phv_out_data_88; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_89 = proc_8_io_pipe_phv_out_data_89; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_90 = proc_8_io_pipe_phv_out_data_90; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_91 = proc_8_io_pipe_phv_out_data_91; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_92 = proc_8_io_pipe_phv_out_data_92; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_93 = proc_8_io_pipe_phv_out_data_93; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_94 = proc_8_io_pipe_phv_out_data_94; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_95 = proc_8_io_pipe_phv_out_data_95; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_96 = proc_8_io_pipe_phv_out_data_96; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_97 = proc_8_io_pipe_phv_out_data_97; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_98 = proc_8_io_pipe_phv_out_data_98; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_99 = proc_8_io_pipe_phv_out_data_99; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_100 = proc_8_io_pipe_phv_out_data_100; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_101 = proc_8_io_pipe_phv_out_data_101; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_102 = proc_8_io_pipe_phv_out_data_102; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_103 = proc_8_io_pipe_phv_out_data_103; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_104 = proc_8_io_pipe_phv_out_data_104; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_105 = proc_8_io_pipe_phv_out_data_105; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_106 = proc_8_io_pipe_phv_out_data_106; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_107 = proc_8_io_pipe_phv_out_data_107; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_108 = proc_8_io_pipe_phv_out_data_108; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_109 = proc_8_io_pipe_phv_out_data_109; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_110 = proc_8_io_pipe_phv_out_data_110; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_111 = proc_8_io_pipe_phv_out_data_111; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_112 = proc_8_io_pipe_phv_out_data_112; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_113 = proc_8_io_pipe_phv_out_data_113; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_114 = proc_8_io_pipe_phv_out_data_114; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_115 = proc_8_io_pipe_phv_out_data_115; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_116 = proc_8_io_pipe_phv_out_data_116; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_117 = proc_8_io_pipe_phv_out_data_117; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_118 = proc_8_io_pipe_phv_out_data_118; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_119 = proc_8_io_pipe_phv_out_data_119; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_120 = proc_8_io_pipe_phv_out_data_120; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_121 = proc_8_io_pipe_phv_out_data_121; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_122 = proc_8_io_pipe_phv_out_data_122; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_123 = proc_8_io_pipe_phv_out_data_123; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_124 = proc_8_io_pipe_phv_out_data_124; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_125 = proc_8_io_pipe_phv_out_data_125; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_126 = proc_8_io_pipe_phv_out_data_126; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_127 = proc_8_io_pipe_phv_out_data_127; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_128 = proc_8_io_pipe_phv_out_data_128; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_129 = proc_8_io_pipe_phv_out_data_129; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_130 = proc_8_io_pipe_phv_out_data_130; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_131 = proc_8_io_pipe_phv_out_data_131; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_132 = proc_8_io_pipe_phv_out_data_132; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_133 = proc_8_io_pipe_phv_out_data_133; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_134 = proc_8_io_pipe_phv_out_data_134; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_135 = proc_8_io_pipe_phv_out_data_135; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_136 = proc_8_io_pipe_phv_out_data_136; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_137 = proc_8_io_pipe_phv_out_data_137; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_138 = proc_8_io_pipe_phv_out_data_138; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_139 = proc_8_io_pipe_phv_out_data_139; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_140 = proc_8_io_pipe_phv_out_data_140; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_141 = proc_8_io_pipe_phv_out_data_141; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_142 = proc_8_io_pipe_phv_out_data_142; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_143 = proc_8_io_pipe_phv_out_data_143; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_144 = proc_8_io_pipe_phv_out_data_144; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_145 = proc_8_io_pipe_phv_out_data_145; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_146 = proc_8_io_pipe_phv_out_data_146; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_147 = proc_8_io_pipe_phv_out_data_147; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_148 = proc_8_io_pipe_phv_out_data_148; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_149 = proc_8_io_pipe_phv_out_data_149; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_150 = proc_8_io_pipe_phv_out_data_150; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_151 = proc_8_io_pipe_phv_out_data_151; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_152 = proc_8_io_pipe_phv_out_data_152; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_153 = proc_8_io_pipe_phv_out_data_153; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_154 = proc_8_io_pipe_phv_out_data_154; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_155 = proc_8_io_pipe_phv_out_data_155; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_156 = proc_8_io_pipe_phv_out_data_156; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_157 = proc_8_io_pipe_phv_out_data_157; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_158 = proc_8_io_pipe_phv_out_data_158; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_159 = proc_8_io_pipe_phv_out_data_159; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_160 = proc_8_io_pipe_phv_out_data_160; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_161 = proc_8_io_pipe_phv_out_data_161; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_162 = proc_8_io_pipe_phv_out_data_162; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_163 = proc_8_io_pipe_phv_out_data_163; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_164 = proc_8_io_pipe_phv_out_data_164; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_165 = proc_8_io_pipe_phv_out_data_165; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_166 = proc_8_io_pipe_phv_out_data_166; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_167 = proc_8_io_pipe_phv_out_data_167; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_168 = proc_8_io_pipe_phv_out_data_168; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_169 = proc_8_io_pipe_phv_out_data_169; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_170 = proc_8_io_pipe_phv_out_data_170; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_171 = proc_8_io_pipe_phv_out_data_171; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_172 = proc_8_io_pipe_phv_out_data_172; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_173 = proc_8_io_pipe_phv_out_data_173; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_174 = proc_8_io_pipe_phv_out_data_174; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_175 = proc_8_io_pipe_phv_out_data_175; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_176 = proc_8_io_pipe_phv_out_data_176; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_177 = proc_8_io_pipe_phv_out_data_177; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_178 = proc_8_io_pipe_phv_out_data_178; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_179 = proc_8_io_pipe_phv_out_data_179; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_180 = proc_8_io_pipe_phv_out_data_180; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_181 = proc_8_io_pipe_phv_out_data_181; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_182 = proc_8_io_pipe_phv_out_data_182; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_183 = proc_8_io_pipe_phv_out_data_183; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_184 = proc_8_io_pipe_phv_out_data_184; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_185 = proc_8_io_pipe_phv_out_data_185; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_186 = proc_8_io_pipe_phv_out_data_186; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_187 = proc_8_io_pipe_phv_out_data_187; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_188 = proc_8_io_pipe_phv_out_data_188; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_189 = proc_8_io_pipe_phv_out_data_189; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_190 = proc_8_io_pipe_phv_out_data_190; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_191 = proc_8_io_pipe_phv_out_data_191; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_192 = proc_8_io_pipe_phv_out_data_192; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_193 = proc_8_io_pipe_phv_out_data_193; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_194 = proc_8_io_pipe_phv_out_data_194; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_195 = proc_8_io_pipe_phv_out_data_195; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_196 = proc_8_io_pipe_phv_out_data_196; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_197 = proc_8_io_pipe_phv_out_data_197; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_198 = proc_8_io_pipe_phv_out_data_198; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_199 = proc_8_io_pipe_phv_out_data_199; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_200 = proc_8_io_pipe_phv_out_data_200; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_201 = proc_8_io_pipe_phv_out_data_201; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_202 = proc_8_io_pipe_phv_out_data_202; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_203 = proc_8_io_pipe_phv_out_data_203; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_204 = proc_8_io_pipe_phv_out_data_204; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_205 = proc_8_io_pipe_phv_out_data_205; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_206 = proc_8_io_pipe_phv_out_data_206; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_207 = proc_8_io_pipe_phv_out_data_207; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_208 = proc_8_io_pipe_phv_out_data_208; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_209 = proc_8_io_pipe_phv_out_data_209; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_210 = proc_8_io_pipe_phv_out_data_210; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_211 = proc_8_io_pipe_phv_out_data_211; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_212 = proc_8_io_pipe_phv_out_data_212; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_213 = proc_8_io_pipe_phv_out_data_213; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_214 = proc_8_io_pipe_phv_out_data_214; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_215 = proc_8_io_pipe_phv_out_data_215; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_216 = proc_8_io_pipe_phv_out_data_216; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_217 = proc_8_io_pipe_phv_out_data_217; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_218 = proc_8_io_pipe_phv_out_data_218; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_219 = proc_8_io_pipe_phv_out_data_219; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_220 = proc_8_io_pipe_phv_out_data_220; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_221 = proc_8_io_pipe_phv_out_data_221; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_222 = proc_8_io_pipe_phv_out_data_222; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_223 = proc_8_io_pipe_phv_out_data_223; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_224 = proc_8_io_pipe_phv_out_data_224; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_225 = proc_8_io_pipe_phv_out_data_225; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_226 = proc_8_io_pipe_phv_out_data_226; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_227 = proc_8_io_pipe_phv_out_data_227; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_228 = proc_8_io_pipe_phv_out_data_228; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_229 = proc_8_io_pipe_phv_out_data_229; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_230 = proc_8_io_pipe_phv_out_data_230; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_231 = proc_8_io_pipe_phv_out_data_231; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_232 = proc_8_io_pipe_phv_out_data_232; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_233 = proc_8_io_pipe_phv_out_data_233; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_234 = proc_8_io_pipe_phv_out_data_234; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_235 = proc_8_io_pipe_phv_out_data_235; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_236 = proc_8_io_pipe_phv_out_data_236; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_237 = proc_8_io_pipe_phv_out_data_237; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_238 = proc_8_io_pipe_phv_out_data_238; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_239 = proc_8_io_pipe_phv_out_data_239; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_240 = proc_8_io_pipe_phv_out_data_240; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_241 = proc_8_io_pipe_phv_out_data_241; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_242 = proc_8_io_pipe_phv_out_data_242; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_243 = proc_8_io_pipe_phv_out_data_243; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_244 = proc_8_io_pipe_phv_out_data_244; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_245 = proc_8_io_pipe_phv_out_data_245; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_246 = proc_8_io_pipe_phv_out_data_246; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_247 = proc_8_io_pipe_phv_out_data_247; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_248 = proc_8_io_pipe_phv_out_data_248; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_249 = proc_8_io_pipe_phv_out_data_249; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_250 = proc_8_io_pipe_phv_out_data_250; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_251 = proc_8_io_pipe_phv_out_data_251; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_252 = proc_8_io_pipe_phv_out_data_252; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_253 = proc_8_io_pipe_phv_out_data_253; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_254 = proc_8_io_pipe_phv_out_data_254; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_255 = proc_8_io_pipe_phv_out_data_255; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_next_processor_id = proc_8_io_pipe_phv_out_next_processor_id; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_next_config_id = proc_8_io_pipe_phv_out_next_config_id; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_is_valid_processor = 4'h9 == proc_8_io_pipe_phv_out_next_processor_id; // @[pisa.scala 36:62]
  assign proc_9_io_mod_mat_mod_en = io_mod_proc_mod_9_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_config_id = io_mod_proc_mod_9_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_9_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_9_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_9_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_9_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_9_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_9_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_9_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_9_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_9_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_9_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_9_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_9_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_9_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_w_en = io_mod_proc_mod_9_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_9_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_w_addr = io_mod_proc_mod_9_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_w_data = io_mod_proc_mod_9_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_9_io_mod_exe_mod_en_0 = io_mod_proc_mod_9_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_9_io_mod_exe_mod_en_1 = io_mod_proc_mod_9_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_9_io_mod_exe_mod_addr = io_mod_proc_mod_9_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_9_io_mod_exe_mod_data_0 = io_mod_proc_mod_9_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_9_io_mod_exe_mod_data_1 = io_mod_proc_mod_9_exe_mod_data_1; // @[pisa.scala 29:20]
  assign proc_10_clock = clock;
  assign proc_10_io_pipe_phv_in_data_0 = proc_9_io_pipe_phv_out_data_0; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_1 = proc_9_io_pipe_phv_out_data_1; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_2 = proc_9_io_pipe_phv_out_data_2; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_3 = proc_9_io_pipe_phv_out_data_3; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_4 = proc_9_io_pipe_phv_out_data_4; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_5 = proc_9_io_pipe_phv_out_data_5; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_6 = proc_9_io_pipe_phv_out_data_6; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_7 = proc_9_io_pipe_phv_out_data_7; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_8 = proc_9_io_pipe_phv_out_data_8; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_9 = proc_9_io_pipe_phv_out_data_9; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_10 = proc_9_io_pipe_phv_out_data_10; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_11 = proc_9_io_pipe_phv_out_data_11; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_12 = proc_9_io_pipe_phv_out_data_12; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_13 = proc_9_io_pipe_phv_out_data_13; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_14 = proc_9_io_pipe_phv_out_data_14; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_15 = proc_9_io_pipe_phv_out_data_15; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_16 = proc_9_io_pipe_phv_out_data_16; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_17 = proc_9_io_pipe_phv_out_data_17; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_18 = proc_9_io_pipe_phv_out_data_18; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_19 = proc_9_io_pipe_phv_out_data_19; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_20 = proc_9_io_pipe_phv_out_data_20; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_21 = proc_9_io_pipe_phv_out_data_21; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_22 = proc_9_io_pipe_phv_out_data_22; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_23 = proc_9_io_pipe_phv_out_data_23; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_24 = proc_9_io_pipe_phv_out_data_24; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_25 = proc_9_io_pipe_phv_out_data_25; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_26 = proc_9_io_pipe_phv_out_data_26; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_27 = proc_9_io_pipe_phv_out_data_27; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_28 = proc_9_io_pipe_phv_out_data_28; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_29 = proc_9_io_pipe_phv_out_data_29; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_30 = proc_9_io_pipe_phv_out_data_30; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_31 = proc_9_io_pipe_phv_out_data_31; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_32 = proc_9_io_pipe_phv_out_data_32; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_33 = proc_9_io_pipe_phv_out_data_33; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_34 = proc_9_io_pipe_phv_out_data_34; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_35 = proc_9_io_pipe_phv_out_data_35; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_36 = proc_9_io_pipe_phv_out_data_36; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_37 = proc_9_io_pipe_phv_out_data_37; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_38 = proc_9_io_pipe_phv_out_data_38; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_39 = proc_9_io_pipe_phv_out_data_39; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_40 = proc_9_io_pipe_phv_out_data_40; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_41 = proc_9_io_pipe_phv_out_data_41; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_42 = proc_9_io_pipe_phv_out_data_42; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_43 = proc_9_io_pipe_phv_out_data_43; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_44 = proc_9_io_pipe_phv_out_data_44; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_45 = proc_9_io_pipe_phv_out_data_45; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_46 = proc_9_io_pipe_phv_out_data_46; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_47 = proc_9_io_pipe_phv_out_data_47; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_48 = proc_9_io_pipe_phv_out_data_48; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_49 = proc_9_io_pipe_phv_out_data_49; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_50 = proc_9_io_pipe_phv_out_data_50; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_51 = proc_9_io_pipe_phv_out_data_51; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_52 = proc_9_io_pipe_phv_out_data_52; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_53 = proc_9_io_pipe_phv_out_data_53; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_54 = proc_9_io_pipe_phv_out_data_54; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_55 = proc_9_io_pipe_phv_out_data_55; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_56 = proc_9_io_pipe_phv_out_data_56; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_57 = proc_9_io_pipe_phv_out_data_57; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_58 = proc_9_io_pipe_phv_out_data_58; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_59 = proc_9_io_pipe_phv_out_data_59; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_60 = proc_9_io_pipe_phv_out_data_60; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_61 = proc_9_io_pipe_phv_out_data_61; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_62 = proc_9_io_pipe_phv_out_data_62; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_63 = proc_9_io_pipe_phv_out_data_63; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_64 = proc_9_io_pipe_phv_out_data_64; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_65 = proc_9_io_pipe_phv_out_data_65; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_66 = proc_9_io_pipe_phv_out_data_66; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_67 = proc_9_io_pipe_phv_out_data_67; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_68 = proc_9_io_pipe_phv_out_data_68; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_69 = proc_9_io_pipe_phv_out_data_69; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_70 = proc_9_io_pipe_phv_out_data_70; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_71 = proc_9_io_pipe_phv_out_data_71; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_72 = proc_9_io_pipe_phv_out_data_72; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_73 = proc_9_io_pipe_phv_out_data_73; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_74 = proc_9_io_pipe_phv_out_data_74; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_75 = proc_9_io_pipe_phv_out_data_75; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_76 = proc_9_io_pipe_phv_out_data_76; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_77 = proc_9_io_pipe_phv_out_data_77; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_78 = proc_9_io_pipe_phv_out_data_78; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_79 = proc_9_io_pipe_phv_out_data_79; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_80 = proc_9_io_pipe_phv_out_data_80; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_81 = proc_9_io_pipe_phv_out_data_81; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_82 = proc_9_io_pipe_phv_out_data_82; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_83 = proc_9_io_pipe_phv_out_data_83; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_84 = proc_9_io_pipe_phv_out_data_84; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_85 = proc_9_io_pipe_phv_out_data_85; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_86 = proc_9_io_pipe_phv_out_data_86; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_87 = proc_9_io_pipe_phv_out_data_87; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_88 = proc_9_io_pipe_phv_out_data_88; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_89 = proc_9_io_pipe_phv_out_data_89; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_90 = proc_9_io_pipe_phv_out_data_90; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_91 = proc_9_io_pipe_phv_out_data_91; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_92 = proc_9_io_pipe_phv_out_data_92; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_93 = proc_9_io_pipe_phv_out_data_93; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_94 = proc_9_io_pipe_phv_out_data_94; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_95 = proc_9_io_pipe_phv_out_data_95; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_96 = proc_9_io_pipe_phv_out_data_96; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_97 = proc_9_io_pipe_phv_out_data_97; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_98 = proc_9_io_pipe_phv_out_data_98; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_99 = proc_9_io_pipe_phv_out_data_99; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_100 = proc_9_io_pipe_phv_out_data_100; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_101 = proc_9_io_pipe_phv_out_data_101; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_102 = proc_9_io_pipe_phv_out_data_102; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_103 = proc_9_io_pipe_phv_out_data_103; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_104 = proc_9_io_pipe_phv_out_data_104; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_105 = proc_9_io_pipe_phv_out_data_105; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_106 = proc_9_io_pipe_phv_out_data_106; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_107 = proc_9_io_pipe_phv_out_data_107; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_108 = proc_9_io_pipe_phv_out_data_108; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_109 = proc_9_io_pipe_phv_out_data_109; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_110 = proc_9_io_pipe_phv_out_data_110; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_111 = proc_9_io_pipe_phv_out_data_111; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_112 = proc_9_io_pipe_phv_out_data_112; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_113 = proc_9_io_pipe_phv_out_data_113; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_114 = proc_9_io_pipe_phv_out_data_114; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_115 = proc_9_io_pipe_phv_out_data_115; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_116 = proc_9_io_pipe_phv_out_data_116; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_117 = proc_9_io_pipe_phv_out_data_117; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_118 = proc_9_io_pipe_phv_out_data_118; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_119 = proc_9_io_pipe_phv_out_data_119; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_120 = proc_9_io_pipe_phv_out_data_120; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_121 = proc_9_io_pipe_phv_out_data_121; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_122 = proc_9_io_pipe_phv_out_data_122; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_123 = proc_9_io_pipe_phv_out_data_123; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_124 = proc_9_io_pipe_phv_out_data_124; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_125 = proc_9_io_pipe_phv_out_data_125; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_126 = proc_9_io_pipe_phv_out_data_126; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_127 = proc_9_io_pipe_phv_out_data_127; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_128 = proc_9_io_pipe_phv_out_data_128; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_129 = proc_9_io_pipe_phv_out_data_129; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_130 = proc_9_io_pipe_phv_out_data_130; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_131 = proc_9_io_pipe_phv_out_data_131; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_132 = proc_9_io_pipe_phv_out_data_132; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_133 = proc_9_io_pipe_phv_out_data_133; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_134 = proc_9_io_pipe_phv_out_data_134; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_135 = proc_9_io_pipe_phv_out_data_135; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_136 = proc_9_io_pipe_phv_out_data_136; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_137 = proc_9_io_pipe_phv_out_data_137; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_138 = proc_9_io_pipe_phv_out_data_138; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_139 = proc_9_io_pipe_phv_out_data_139; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_140 = proc_9_io_pipe_phv_out_data_140; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_141 = proc_9_io_pipe_phv_out_data_141; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_142 = proc_9_io_pipe_phv_out_data_142; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_143 = proc_9_io_pipe_phv_out_data_143; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_144 = proc_9_io_pipe_phv_out_data_144; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_145 = proc_9_io_pipe_phv_out_data_145; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_146 = proc_9_io_pipe_phv_out_data_146; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_147 = proc_9_io_pipe_phv_out_data_147; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_148 = proc_9_io_pipe_phv_out_data_148; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_149 = proc_9_io_pipe_phv_out_data_149; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_150 = proc_9_io_pipe_phv_out_data_150; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_151 = proc_9_io_pipe_phv_out_data_151; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_152 = proc_9_io_pipe_phv_out_data_152; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_153 = proc_9_io_pipe_phv_out_data_153; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_154 = proc_9_io_pipe_phv_out_data_154; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_155 = proc_9_io_pipe_phv_out_data_155; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_156 = proc_9_io_pipe_phv_out_data_156; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_157 = proc_9_io_pipe_phv_out_data_157; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_158 = proc_9_io_pipe_phv_out_data_158; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_159 = proc_9_io_pipe_phv_out_data_159; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_160 = proc_9_io_pipe_phv_out_data_160; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_161 = proc_9_io_pipe_phv_out_data_161; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_162 = proc_9_io_pipe_phv_out_data_162; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_163 = proc_9_io_pipe_phv_out_data_163; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_164 = proc_9_io_pipe_phv_out_data_164; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_165 = proc_9_io_pipe_phv_out_data_165; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_166 = proc_9_io_pipe_phv_out_data_166; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_167 = proc_9_io_pipe_phv_out_data_167; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_168 = proc_9_io_pipe_phv_out_data_168; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_169 = proc_9_io_pipe_phv_out_data_169; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_170 = proc_9_io_pipe_phv_out_data_170; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_171 = proc_9_io_pipe_phv_out_data_171; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_172 = proc_9_io_pipe_phv_out_data_172; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_173 = proc_9_io_pipe_phv_out_data_173; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_174 = proc_9_io_pipe_phv_out_data_174; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_175 = proc_9_io_pipe_phv_out_data_175; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_176 = proc_9_io_pipe_phv_out_data_176; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_177 = proc_9_io_pipe_phv_out_data_177; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_178 = proc_9_io_pipe_phv_out_data_178; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_179 = proc_9_io_pipe_phv_out_data_179; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_180 = proc_9_io_pipe_phv_out_data_180; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_181 = proc_9_io_pipe_phv_out_data_181; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_182 = proc_9_io_pipe_phv_out_data_182; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_183 = proc_9_io_pipe_phv_out_data_183; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_184 = proc_9_io_pipe_phv_out_data_184; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_185 = proc_9_io_pipe_phv_out_data_185; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_186 = proc_9_io_pipe_phv_out_data_186; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_187 = proc_9_io_pipe_phv_out_data_187; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_188 = proc_9_io_pipe_phv_out_data_188; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_189 = proc_9_io_pipe_phv_out_data_189; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_190 = proc_9_io_pipe_phv_out_data_190; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_191 = proc_9_io_pipe_phv_out_data_191; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_192 = proc_9_io_pipe_phv_out_data_192; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_193 = proc_9_io_pipe_phv_out_data_193; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_194 = proc_9_io_pipe_phv_out_data_194; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_195 = proc_9_io_pipe_phv_out_data_195; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_196 = proc_9_io_pipe_phv_out_data_196; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_197 = proc_9_io_pipe_phv_out_data_197; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_198 = proc_9_io_pipe_phv_out_data_198; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_199 = proc_9_io_pipe_phv_out_data_199; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_200 = proc_9_io_pipe_phv_out_data_200; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_201 = proc_9_io_pipe_phv_out_data_201; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_202 = proc_9_io_pipe_phv_out_data_202; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_203 = proc_9_io_pipe_phv_out_data_203; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_204 = proc_9_io_pipe_phv_out_data_204; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_205 = proc_9_io_pipe_phv_out_data_205; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_206 = proc_9_io_pipe_phv_out_data_206; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_207 = proc_9_io_pipe_phv_out_data_207; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_208 = proc_9_io_pipe_phv_out_data_208; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_209 = proc_9_io_pipe_phv_out_data_209; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_210 = proc_9_io_pipe_phv_out_data_210; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_211 = proc_9_io_pipe_phv_out_data_211; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_212 = proc_9_io_pipe_phv_out_data_212; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_213 = proc_9_io_pipe_phv_out_data_213; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_214 = proc_9_io_pipe_phv_out_data_214; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_215 = proc_9_io_pipe_phv_out_data_215; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_216 = proc_9_io_pipe_phv_out_data_216; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_217 = proc_9_io_pipe_phv_out_data_217; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_218 = proc_9_io_pipe_phv_out_data_218; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_219 = proc_9_io_pipe_phv_out_data_219; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_220 = proc_9_io_pipe_phv_out_data_220; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_221 = proc_9_io_pipe_phv_out_data_221; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_222 = proc_9_io_pipe_phv_out_data_222; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_223 = proc_9_io_pipe_phv_out_data_223; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_224 = proc_9_io_pipe_phv_out_data_224; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_225 = proc_9_io_pipe_phv_out_data_225; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_226 = proc_9_io_pipe_phv_out_data_226; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_227 = proc_9_io_pipe_phv_out_data_227; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_228 = proc_9_io_pipe_phv_out_data_228; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_229 = proc_9_io_pipe_phv_out_data_229; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_230 = proc_9_io_pipe_phv_out_data_230; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_231 = proc_9_io_pipe_phv_out_data_231; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_232 = proc_9_io_pipe_phv_out_data_232; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_233 = proc_9_io_pipe_phv_out_data_233; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_234 = proc_9_io_pipe_phv_out_data_234; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_235 = proc_9_io_pipe_phv_out_data_235; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_236 = proc_9_io_pipe_phv_out_data_236; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_237 = proc_9_io_pipe_phv_out_data_237; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_238 = proc_9_io_pipe_phv_out_data_238; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_239 = proc_9_io_pipe_phv_out_data_239; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_240 = proc_9_io_pipe_phv_out_data_240; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_241 = proc_9_io_pipe_phv_out_data_241; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_242 = proc_9_io_pipe_phv_out_data_242; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_243 = proc_9_io_pipe_phv_out_data_243; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_244 = proc_9_io_pipe_phv_out_data_244; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_245 = proc_9_io_pipe_phv_out_data_245; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_246 = proc_9_io_pipe_phv_out_data_246; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_247 = proc_9_io_pipe_phv_out_data_247; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_248 = proc_9_io_pipe_phv_out_data_248; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_249 = proc_9_io_pipe_phv_out_data_249; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_250 = proc_9_io_pipe_phv_out_data_250; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_251 = proc_9_io_pipe_phv_out_data_251; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_252 = proc_9_io_pipe_phv_out_data_252; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_253 = proc_9_io_pipe_phv_out_data_253; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_254 = proc_9_io_pipe_phv_out_data_254; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_255 = proc_9_io_pipe_phv_out_data_255; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_next_processor_id = proc_9_io_pipe_phv_out_next_processor_id; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_next_config_id = proc_9_io_pipe_phv_out_next_config_id; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_is_valid_processor = 4'ha == proc_9_io_pipe_phv_out_next_processor_id; // @[pisa.scala 36:62]
  assign proc_10_io_mod_mat_mod_en = io_mod_proc_mod_10_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_config_id = io_mod_proc_mod_10_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_10_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_10_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_10_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_10_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_10_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_10_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_10_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_10_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_10_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_10_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_10_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_10_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_10_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_w_en = io_mod_proc_mod_10_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_10_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_w_addr = io_mod_proc_mod_10_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_w_data = io_mod_proc_mod_10_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_10_io_mod_exe_mod_en_0 = io_mod_proc_mod_10_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_10_io_mod_exe_mod_en_1 = io_mod_proc_mod_10_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_10_io_mod_exe_mod_addr = io_mod_proc_mod_10_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_10_io_mod_exe_mod_data_0 = io_mod_proc_mod_10_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_10_io_mod_exe_mod_data_1 = io_mod_proc_mod_10_exe_mod_data_1; // @[pisa.scala 29:20]
  assign proc_11_clock = clock;
  assign proc_11_io_pipe_phv_in_data_0 = proc_10_io_pipe_phv_out_data_0; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_1 = proc_10_io_pipe_phv_out_data_1; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_2 = proc_10_io_pipe_phv_out_data_2; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_3 = proc_10_io_pipe_phv_out_data_3; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_4 = proc_10_io_pipe_phv_out_data_4; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_5 = proc_10_io_pipe_phv_out_data_5; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_6 = proc_10_io_pipe_phv_out_data_6; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_7 = proc_10_io_pipe_phv_out_data_7; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_8 = proc_10_io_pipe_phv_out_data_8; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_9 = proc_10_io_pipe_phv_out_data_9; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_10 = proc_10_io_pipe_phv_out_data_10; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_11 = proc_10_io_pipe_phv_out_data_11; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_12 = proc_10_io_pipe_phv_out_data_12; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_13 = proc_10_io_pipe_phv_out_data_13; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_14 = proc_10_io_pipe_phv_out_data_14; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_15 = proc_10_io_pipe_phv_out_data_15; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_16 = proc_10_io_pipe_phv_out_data_16; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_17 = proc_10_io_pipe_phv_out_data_17; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_18 = proc_10_io_pipe_phv_out_data_18; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_19 = proc_10_io_pipe_phv_out_data_19; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_20 = proc_10_io_pipe_phv_out_data_20; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_21 = proc_10_io_pipe_phv_out_data_21; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_22 = proc_10_io_pipe_phv_out_data_22; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_23 = proc_10_io_pipe_phv_out_data_23; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_24 = proc_10_io_pipe_phv_out_data_24; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_25 = proc_10_io_pipe_phv_out_data_25; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_26 = proc_10_io_pipe_phv_out_data_26; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_27 = proc_10_io_pipe_phv_out_data_27; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_28 = proc_10_io_pipe_phv_out_data_28; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_29 = proc_10_io_pipe_phv_out_data_29; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_30 = proc_10_io_pipe_phv_out_data_30; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_31 = proc_10_io_pipe_phv_out_data_31; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_32 = proc_10_io_pipe_phv_out_data_32; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_33 = proc_10_io_pipe_phv_out_data_33; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_34 = proc_10_io_pipe_phv_out_data_34; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_35 = proc_10_io_pipe_phv_out_data_35; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_36 = proc_10_io_pipe_phv_out_data_36; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_37 = proc_10_io_pipe_phv_out_data_37; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_38 = proc_10_io_pipe_phv_out_data_38; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_39 = proc_10_io_pipe_phv_out_data_39; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_40 = proc_10_io_pipe_phv_out_data_40; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_41 = proc_10_io_pipe_phv_out_data_41; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_42 = proc_10_io_pipe_phv_out_data_42; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_43 = proc_10_io_pipe_phv_out_data_43; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_44 = proc_10_io_pipe_phv_out_data_44; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_45 = proc_10_io_pipe_phv_out_data_45; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_46 = proc_10_io_pipe_phv_out_data_46; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_47 = proc_10_io_pipe_phv_out_data_47; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_48 = proc_10_io_pipe_phv_out_data_48; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_49 = proc_10_io_pipe_phv_out_data_49; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_50 = proc_10_io_pipe_phv_out_data_50; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_51 = proc_10_io_pipe_phv_out_data_51; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_52 = proc_10_io_pipe_phv_out_data_52; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_53 = proc_10_io_pipe_phv_out_data_53; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_54 = proc_10_io_pipe_phv_out_data_54; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_55 = proc_10_io_pipe_phv_out_data_55; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_56 = proc_10_io_pipe_phv_out_data_56; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_57 = proc_10_io_pipe_phv_out_data_57; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_58 = proc_10_io_pipe_phv_out_data_58; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_59 = proc_10_io_pipe_phv_out_data_59; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_60 = proc_10_io_pipe_phv_out_data_60; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_61 = proc_10_io_pipe_phv_out_data_61; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_62 = proc_10_io_pipe_phv_out_data_62; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_63 = proc_10_io_pipe_phv_out_data_63; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_64 = proc_10_io_pipe_phv_out_data_64; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_65 = proc_10_io_pipe_phv_out_data_65; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_66 = proc_10_io_pipe_phv_out_data_66; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_67 = proc_10_io_pipe_phv_out_data_67; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_68 = proc_10_io_pipe_phv_out_data_68; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_69 = proc_10_io_pipe_phv_out_data_69; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_70 = proc_10_io_pipe_phv_out_data_70; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_71 = proc_10_io_pipe_phv_out_data_71; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_72 = proc_10_io_pipe_phv_out_data_72; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_73 = proc_10_io_pipe_phv_out_data_73; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_74 = proc_10_io_pipe_phv_out_data_74; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_75 = proc_10_io_pipe_phv_out_data_75; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_76 = proc_10_io_pipe_phv_out_data_76; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_77 = proc_10_io_pipe_phv_out_data_77; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_78 = proc_10_io_pipe_phv_out_data_78; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_79 = proc_10_io_pipe_phv_out_data_79; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_80 = proc_10_io_pipe_phv_out_data_80; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_81 = proc_10_io_pipe_phv_out_data_81; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_82 = proc_10_io_pipe_phv_out_data_82; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_83 = proc_10_io_pipe_phv_out_data_83; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_84 = proc_10_io_pipe_phv_out_data_84; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_85 = proc_10_io_pipe_phv_out_data_85; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_86 = proc_10_io_pipe_phv_out_data_86; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_87 = proc_10_io_pipe_phv_out_data_87; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_88 = proc_10_io_pipe_phv_out_data_88; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_89 = proc_10_io_pipe_phv_out_data_89; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_90 = proc_10_io_pipe_phv_out_data_90; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_91 = proc_10_io_pipe_phv_out_data_91; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_92 = proc_10_io_pipe_phv_out_data_92; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_93 = proc_10_io_pipe_phv_out_data_93; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_94 = proc_10_io_pipe_phv_out_data_94; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_95 = proc_10_io_pipe_phv_out_data_95; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_96 = proc_10_io_pipe_phv_out_data_96; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_97 = proc_10_io_pipe_phv_out_data_97; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_98 = proc_10_io_pipe_phv_out_data_98; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_99 = proc_10_io_pipe_phv_out_data_99; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_100 = proc_10_io_pipe_phv_out_data_100; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_101 = proc_10_io_pipe_phv_out_data_101; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_102 = proc_10_io_pipe_phv_out_data_102; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_103 = proc_10_io_pipe_phv_out_data_103; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_104 = proc_10_io_pipe_phv_out_data_104; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_105 = proc_10_io_pipe_phv_out_data_105; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_106 = proc_10_io_pipe_phv_out_data_106; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_107 = proc_10_io_pipe_phv_out_data_107; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_108 = proc_10_io_pipe_phv_out_data_108; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_109 = proc_10_io_pipe_phv_out_data_109; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_110 = proc_10_io_pipe_phv_out_data_110; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_111 = proc_10_io_pipe_phv_out_data_111; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_112 = proc_10_io_pipe_phv_out_data_112; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_113 = proc_10_io_pipe_phv_out_data_113; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_114 = proc_10_io_pipe_phv_out_data_114; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_115 = proc_10_io_pipe_phv_out_data_115; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_116 = proc_10_io_pipe_phv_out_data_116; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_117 = proc_10_io_pipe_phv_out_data_117; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_118 = proc_10_io_pipe_phv_out_data_118; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_119 = proc_10_io_pipe_phv_out_data_119; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_120 = proc_10_io_pipe_phv_out_data_120; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_121 = proc_10_io_pipe_phv_out_data_121; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_122 = proc_10_io_pipe_phv_out_data_122; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_123 = proc_10_io_pipe_phv_out_data_123; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_124 = proc_10_io_pipe_phv_out_data_124; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_125 = proc_10_io_pipe_phv_out_data_125; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_126 = proc_10_io_pipe_phv_out_data_126; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_127 = proc_10_io_pipe_phv_out_data_127; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_128 = proc_10_io_pipe_phv_out_data_128; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_129 = proc_10_io_pipe_phv_out_data_129; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_130 = proc_10_io_pipe_phv_out_data_130; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_131 = proc_10_io_pipe_phv_out_data_131; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_132 = proc_10_io_pipe_phv_out_data_132; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_133 = proc_10_io_pipe_phv_out_data_133; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_134 = proc_10_io_pipe_phv_out_data_134; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_135 = proc_10_io_pipe_phv_out_data_135; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_136 = proc_10_io_pipe_phv_out_data_136; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_137 = proc_10_io_pipe_phv_out_data_137; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_138 = proc_10_io_pipe_phv_out_data_138; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_139 = proc_10_io_pipe_phv_out_data_139; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_140 = proc_10_io_pipe_phv_out_data_140; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_141 = proc_10_io_pipe_phv_out_data_141; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_142 = proc_10_io_pipe_phv_out_data_142; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_143 = proc_10_io_pipe_phv_out_data_143; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_144 = proc_10_io_pipe_phv_out_data_144; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_145 = proc_10_io_pipe_phv_out_data_145; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_146 = proc_10_io_pipe_phv_out_data_146; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_147 = proc_10_io_pipe_phv_out_data_147; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_148 = proc_10_io_pipe_phv_out_data_148; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_149 = proc_10_io_pipe_phv_out_data_149; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_150 = proc_10_io_pipe_phv_out_data_150; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_151 = proc_10_io_pipe_phv_out_data_151; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_152 = proc_10_io_pipe_phv_out_data_152; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_153 = proc_10_io_pipe_phv_out_data_153; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_154 = proc_10_io_pipe_phv_out_data_154; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_155 = proc_10_io_pipe_phv_out_data_155; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_156 = proc_10_io_pipe_phv_out_data_156; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_157 = proc_10_io_pipe_phv_out_data_157; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_158 = proc_10_io_pipe_phv_out_data_158; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_159 = proc_10_io_pipe_phv_out_data_159; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_160 = proc_10_io_pipe_phv_out_data_160; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_161 = proc_10_io_pipe_phv_out_data_161; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_162 = proc_10_io_pipe_phv_out_data_162; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_163 = proc_10_io_pipe_phv_out_data_163; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_164 = proc_10_io_pipe_phv_out_data_164; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_165 = proc_10_io_pipe_phv_out_data_165; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_166 = proc_10_io_pipe_phv_out_data_166; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_167 = proc_10_io_pipe_phv_out_data_167; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_168 = proc_10_io_pipe_phv_out_data_168; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_169 = proc_10_io_pipe_phv_out_data_169; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_170 = proc_10_io_pipe_phv_out_data_170; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_171 = proc_10_io_pipe_phv_out_data_171; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_172 = proc_10_io_pipe_phv_out_data_172; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_173 = proc_10_io_pipe_phv_out_data_173; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_174 = proc_10_io_pipe_phv_out_data_174; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_175 = proc_10_io_pipe_phv_out_data_175; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_176 = proc_10_io_pipe_phv_out_data_176; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_177 = proc_10_io_pipe_phv_out_data_177; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_178 = proc_10_io_pipe_phv_out_data_178; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_179 = proc_10_io_pipe_phv_out_data_179; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_180 = proc_10_io_pipe_phv_out_data_180; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_181 = proc_10_io_pipe_phv_out_data_181; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_182 = proc_10_io_pipe_phv_out_data_182; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_183 = proc_10_io_pipe_phv_out_data_183; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_184 = proc_10_io_pipe_phv_out_data_184; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_185 = proc_10_io_pipe_phv_out_data_185; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_186 = proc_10_io_pipe_phv_out_data_186; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_187 = proc_10_io_pipe_phv_out_data_187; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_188 = proc_10_io_pipe_phv_out_data_188; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_189 = proc_10_io_pipe_phv_out_data_189; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_190 = proc_10_io_pipe_phv_out_data_190; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_191 = proc_10_io_pipe_phv_out_data_191; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_192 = proc_10_io_pipe_phv_out_data_192; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_193 = proc_10_io_pipe_phv_out_data_193; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_194 = proc_10_io_pipe_phv_out_data_194; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_195 = proc_10_io_pipe_phv_out_data_195; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_196 = proc_10_io_pipe_phv_out_data_196; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_197 = proc_10_io_pipe_phv_out_data_197; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_198 = proc_10_io_pipe_phv_out_data_198; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_199 = proc_10_io_pipe_phv_out_data_199; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_200 = proc_10_io_pipe_phv_out_data_200; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_201 = proc_10_io_pipe_phv_out_data_201; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_202 = proc_10_io_pipe_phv_out_data_202; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_203 = proc_10_io_pipe_phv_out_data_203; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_204 = proc_10_io_pipe_phv_out_data_204; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_205 = proc_10_io_pipe_phv_out_data_205; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_206 = proc_10_io_pipe_phv_out_data_206; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_207 = proc_10_io_pipe_phv_out_data_207; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_208 = proc_10_io_pipe_phv_out_data_208; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_209 = proc_10_io_pipe_phv_out_data_209; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_210 = proc_10_io_pipe_phv_out_data_210; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_211 = proc_10_io_pipe_phv_out_data_211; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_212 = proc_10_io_pipe_phv_out_data_212; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_213 = proc_10_io_pipe_phv_out_data_213; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_214 = proc_10_io_pipe_phv_out_data_214; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_215 = proc_10_io_pipe_phv_out_data_215; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_216 = proc_10_io_pipe_phv_out_data_216; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_217 = proc_10_io_pipe_phv_out_data_217; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_218 = proc_10_io_pipe_phv_out_data_218; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_219 = proc_10_io_pipe_phv_out_data_219; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_220 = proc_10_io_pipe_phv_out_data_220; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_221 = proc_10_io_pipe_phv_out_data_221; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_222 = proc_10_io_pipe_phv_out_data_222; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_223 = proc_10_io_pipe_phv_out_data_223; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_224 = proc_10_io_pipe_phv_out_data_224; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_225 = proc_10_io_pipe_phv_out_data_225; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_226 = proc_10_io_pipe_phv_out_data_226; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_227 = proc_10_io_pipe_phv_out_data_227; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_228 = proc_10_io_pipe_phv_out_data_228; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_229 = proc_10_io_pipe_phv_out_data_229; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_230 = proc_10_io_pipe_phv_out_data_230; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_231 = proc_10_io_pipe_phv_out_data_231; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_232 = proc_10_io_pipe_phv_out_data_232; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_233 = proc_10_io_pipe_phv_out_data_233; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_234 = proc_10_io_pipe_phv_out_data_234; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_235 = proc_10_io_pipe_phv_out_data_235; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_236 = proc_10_io_pipe_phv_out_data_236; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_237 = proc_10_io_pipe_phv_out_data_237; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_238 = proc_10_io_pipe_phv_out_data_238; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_239 = proc_10_io_pipe_phv_out_data_239; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_240 = proc_10_io_pipe_phv_out_data_240; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_241 = proc_10_io_pipe_phv_out_data_241; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_242 = proc_10_io_pipe_phv_out_data_242; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_243 = proc_10_io_pipe_phv_out_data_243; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_244 = proc_10_io_pipe_phv_out_data_244; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_245 = proc_10_io_pipe_phv_out_data_245; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_246 = proc_10_io_pipe_phv_out_data_246; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_247 = proc_10_io_pipe_phv_out_data_247; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_248 = proc_10_io_pipe_phv_out_data_248; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_249 = proc_10_io_pipe_phv_out_data_249; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_250 = proc_10_io_pipe_phv_out_data_250; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_251 = proc_10_io_pipe_phv_out_data_251; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_252 = proc_10_io_pipe_phv_out_data_252; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_253 = proc_10_io_pipe_phv_out_data_253; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_254 = proc_10_io_pipe_phv_out_data_254; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_255 = proc_10_io_pipe_phv_out_data_255; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_next_processor_id = proc_10_io_pipe_phv_out_next_processor_id; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_next_config_id = proc_10_io_pipe_phv_out_next_config_id; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_is_valid_processor = 4'hb == proc_10_io_pipe_phv_out_next_processor_id; // @[pisa.scala 36:62]
  assign proc_11_io_mod_mat_mod_en = io_mod_proc_mod_11_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_config_id = io_mod_proc_mod_11_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_11_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_11_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_11_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_11_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_11_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_11_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_11_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_11_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_11_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_11_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_11_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_11_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_11_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_w_en = io_mod_proc_mod_11_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_11_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_w_addr = io_mod_proc_mod_11_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_w_data = io_mod_proc_mod_11_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_11_io_mod_exe_mod_en_0 = io_mod_proc_mod_11_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_11_io_mod_exe_mod_en_1 = io_mod_proc_mod_11_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_11_io_mod_exe_mod_addr = io_mod_proc_mod_11_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_11_io_mod_exe_mod_data_0 = io_mod_proc_mod_11_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_11_io_mod_exe_mod_data_1 = io_mod_proc_mod_11_exe_mod_data_1; // @[pisa.scala 29:20]
endmodule
