module MatcherPISA(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [7:0]  io_pipe_phv_in_data_160,
  input  [7:0]  io_pipe_phv_in_data_161,
  input  [7:0]  io_pipe_phv_in_data_162,
  input  [7:0]  io_pipe_phv_in_data_163,
  input  [7:0]  io_pipe_phv_in_data_164,
  input  [7:0]  io_pipe_phv_in_data_165,
  input  [7:0]  io_pipe_phv_in_data_166,
  input  [7:0]  io_pipe_phv_in_data_167,
  input  [7:0]  io_pipe_phv_in_data_168,
  input  [7:0]  io_pipe_phv_in_data_169,
  input  [7:0]  io_pipe_phv_in_data_170,
  input  [7:0]  io_pipe_phv_in_data_171,
  input  [7:0]  io_pipe_phv_in_data_172,
  input  [7:0]  io_pipe_phv_in_data_173,
  input  [7:0]  io_pipe_phv_in_data_174,
  input  [7:0]  io_pipe_phv_in_data_175,
  input  [7:0]  io_pipe_phv_in_data_176,
  input  [7:0]  io_pipe_phv_in_data_177,
  input  [7:0]  io_pipe_phv_in_data_178,
  input  [7:0]  io_pipe_phv_in_data_179,
  input  [7:0]  io_pipe_phv_in_data_180,
  input  [7:0]  io_pipe_phv_in_data_181,
  input  [7:0]  io_pipe_phv_in_data_182,
  input  [7:0]  io_pipe_phv_in_data_183,
  input  [7:0]  io_pipe_phv_in_data_184,
  input  [7:0]  io_pipe_phv_in_data_185,
  input  [7:0]  io_pipe_phv_in_data_186,
  input  [7:0]  io_pipe_phv_in_data_187,
  input  [7:0]  io_pipe_phv_in_data_188,
  input  [7:0]  io_pipe_phv_in_data_189,
  input  [7:0]  io_pipe_phv_in_data_190,
  input  [7:0]  io_pipe_phv_in_data_191,
  input  [7:0]  io_pipe_phv_in_data_192,
  input  [7:0]  io_pipe_phv_in_data_193,
  input  [7:0]  io_pipe_phv_in_data_194,
  input  [7:0]  io_pipe_phv_in_data_195,
  input  [7:0]  io_pipe_phv_in_data_196,
  input  [7:0]  io_pipe_phv_in_data_197,
  input  [7:0]  io_pipe_phv_in_data_198,
  input  [7:0]  io_pipe_phv_in_data_199,
  input  [7:0]  io_pipe_phv_in_data_200,
  input  [7:0]  io_pipe_phv_in_data_201,
  input  [7:0]  io_pipe_phv_in_data_202,
  input  [7:0]  io_pipe_phv_in_data_203,
  input  [7:0]  io_pipe_phv_in_data_204,
  input  [7:0]  io_pipe_phv_in_data_205,
  input  [7:0]  io_pipe_phv_in_data_206,
  input  [7:0]  io_pipe_phv_in_data_207,
  input  [7:0]  io_pipe_phv_in_data_208,
  input  [7:0]  io_pipe_phv_in_data_209,
  input  [7:0]  io_pipe_phv_in_data_210,
  input  [7:0]  io_pipe_phv_in_data_211,
  input  [7:0]  io_pipe_phv_in_data_212,
  input  [7:0]  io_pipe_phv_in_data_213,
  input  [7:0]  io_pipe_phv_in_data_214,
  input  [7:0]  io_pipe_phv_in_data_215,
  input  [7:0]  io_pipe_phv_in_data_216,
  input  [7:0]  io_pipe_phv_in_data_217,
  input  [7:0]  io_pipe_phv_in_data_218,
  input  [7:0]  io_pipe_phv_in_data_219,
  input  [7:0]  io_pipe_phv_in_data_220,
  input  [7:0]  io_pipe_phv_in_data_221,
  input  [7:0]  io_pipe_phv_in_data_222,
  input  [7:0]  io_pipe_phv_in_data_223,
  input  [7:0]  io_pipe_phv_in_data_224,
  input  [7:0]  io_pipe_phv_in_data_225,
  input  [7:0]  io_pipe_phv_in_data_226,
  input  [7:0]  io_pipe_phv_in_data_227,
  input  [7:0]  io_pipe_phv_in_data_228,
  input  [7:0]  io_pipe_phv_in_data_229,
  input  [7:0]  io_pipe_phv_in_data_230,
  input  [7:0]  io_pipe_phv_in_data_231,
  input  [7:0]  io_pipe_phv_in_data_232,
  input  [7:0]  io_pipe_phv_in_data_233,
  input  [7:0]  io_pipe_phv_in_data_234,
  input  [7:0]  io_pipe_phv_in_data_235,
  input  [7:0]  io_pipe_phv_in_data_236,
  input  [7:0]  io_pipe_phv_in_data_237,
  input  [7:0]  io_pipe_phv_in_data_238,
  input  [7:0]  io_pipe_phv_in_data_239,
  input  [7:0]  io_pipe_phv_in_data_240,
  input  [7:0]  io_pipe_phv_in_data_241,
  input  [7:0]  io_pipe_phv_in_data_242,
  input  [7:0]  io_pipe_phv_in_data_243,
  input  [7:0]  io_pipe_phv_in_data_244,
  input  [7:0]  io_pipe_phv_in_data_245,
  input  [7:0]  io_pipe_phv_in_data_246,
  input  [7:0]  io_pipe_phv_in_data_247,
  input  [7:0]  io_pipe_phv_in_data_248,
  input  [7:0]  io_pipe_phv_in_data_249,
  input  [7:0]  io_pipe_phv_in_data_250,
  input  [7:0]  io_pipe_phv_in_data_251,
  input  [7:0]  io_pipe_phv_in_data_252,
  input  [7:0]  io_pipe_phv_in_data_253,
  input  [7:0]  io_pipe_phv_in_data_254,
  input  [7:0]  io_pipe_phv_in_data_255,
  input  [7:0]  io_pipe_phv_in_data_256,
  input  [7:0]  io_pipe_phv_in_data_257,
  input  [7:0]  io_pipe_phv_in_data_258,
  input  [7:0]  io_pipe_phv_in_data_259,
  input  [7:0]  io_pipe_phv_in_data_260,
  input  [7:0]  io_pipe_phv_in_data_261,
  input  [7:0]  io_pipe_phv_in_data_262,
  input  [7:0]  io_pipe_phv_in_data_263,
  input  [7:0]  io_pipe_phv_in_data_264,
  input  [7:0]  io_pipe_phv_in_data_265,
  input  [7:0]  io_pipe_phv_in_data_266,
  input  [7:0]  io_pipe_phv_in_data_267,
  input  [7:0]  io_pipe_phv_in_data_268,
  input  [7:0]  io_pipe_phv_in_data_269,
  input  [7:0]  io_pipe_phv_in_data_270,
  input  [7:0]  io_pipe_phv_in_data_271,
  input  [7:0]  io_pipe_phv_in_data_272,
  input  [7:0]  io_pipe_phv_in_data_273,
  input  [7:0]  io_pipe_phv_in_data_274,
  input  [7:0]  io_pipe_phv_in_data_275,
  input  [7:0]  io_pipe_phv_in_data_276,
  input  [7:0]  io_pipe_phv_in_data_277,
  input  [7:0]  io_pipe_phv_in_data_278,
  input  [7:0]  io_pipe_phv_in_data_279,
  input  [7:0]  io_pipe_phv_in_data_280,
  input  [7:0]  io_pipe_phv_in_data_281,
  input  [7:0]  io_pipe_phv_in_data_282,
  input  [7:0]  io_pipe_phv_in_data_283,
  input  [7:0]  io_pipe_phv_in_data_284,
  input  [7:0]  io_pipe_phv_in_data_285,
  input  [7:0]  io_pipe_phv_in_data_286,
  input  [7:0]  io_pipe_phv_in_data_287,
  input  [7:0]  io_pipe_phv_in_data_288,
  input  [7:0]  io_pipe_phv_in_data_289,
  input  [7:0]  io_pipe_phv_in_data_290,
  input  [7:0]  io_pipe_phv_in_data_291,
  input  [7:0]  io_pipe_phv_in_data_292,
  input  [7:0]  io_pipe_phv_in_data_293,
  input  [7:0]  io_pipe_phv_in_data_294,
  input  [7:0]  io_pipe_phv_in_data_295,
  input  [7:0]  io_pipe_phv_in_data_296,
  input  [7:0]  io_pipe_phv_in_data_297,
  input  [7:0]  io_pipe_phv_in_data_298,
  input  [7:0]  io_pipe_phv_in_data_299,
  input  [7:0]  io_pipe_phv_in_data_300,
  input  [7:0]  io_pipe_phv_in_data_301,
  input  [7:0]  io_pipe_phv_in_data_302,
  input  [7:0]  io_pipe_phv_in_data_303,
  input  [7:0]  io_pipe_phv_in_data_304,
  input  [7:0]  io_pipe_phv_in_data_305,
  input  [7:0]  io_pipe_phv_in_data_306,
  input  [7:0]  io_pipe_phv_in_data_307,
  input  [7:0]  io_pipe_phv_in_data_308,
  input  [7:0]  io_pipe_phv_in_data_309,
  input  [7:0]  io_pipe_phv_in_data_310,
  input  [7:0]  io_pipe_phv_in_data_311,
  input  [7:0]  io_pipe_phv_in_data_312,
  input  [7:0]  io_pipe_phv_in_data_313,
  input  [7:0]  io_pipe_phv_in_data_314,
  input  [7:0]  io_pipe_phv_in_data_315,
  input  [7:0]  io_pipe_phv_in_data_316,
  input  [7:0]  io_pipe_phv_in_data_317,
  input  [7:0]  io_pipe_phv_in_data_318,
  input  [7:0]  io_pipe_phv_in_data_319,
  input  [7:0]  io_pipe_phv_in_data_320,
  input  [7:0]  io_pipe_phv_in_data_321,
  input  [7:0]  io_pipe_phv_in_data_322,
  input  [7:0]  io_pipe_phv_in_data_323,
  input  [7:0]  io_pipe_phv_in_data_324,
  input  [7:0]  io_pipe_phv_in_data_325,
  input  [7:0]  io_pipe_phv_in_data_326,
  input  [7:0]  io_pipe_phv_in_data_327,
  input  [7:0]  io_pipe_phv_in_data_328,
  input  [7:0]  io_pipe_phv_in_data_329,
  input  [7:0]  io_pipe_phv_in_data_330,
  input  [7:0]  io_pipe_phv_in_data_331,
  input  [7:0]  io_pipe_phv_in_data_332,
  input  [7:0]  io_pipe_phv_in_data_333,
  input  [7:0]  io_pipe_phv_in_data_334,
  input  [7:0]  io_pipe_phv_in_data_335,
  input  [7:0]  io_pipe_phv_in_data_336,
  input  [7:0]  io_pipe_phv_in_data_337,
  input  [7:0]  io_pipe_phv_in_data_338,
  input  [7:0]  io_pipe_phv_in_data_339,
  input  [7:0]  io_pipe_phv_in_data_340,
  input  [7:0]  io_pipe_phv_in_data_341,
  input  [7:0]  io_pipe_phv_in_data_342,
  input  [7:0]  io_pipe_phv_in_data_343,
  input  [7:0]  io_pipe_phv_in_data_344,
  input  [7:0]  io_pipe_phv_in_data_345,
  input  [7:0]  io_pipe_phv_in_data_346,
  input  [7:0]  io_pipe_phv_in_data_347,
  input  [7:0]  io_pipe_phv_in_data_348,
  input  [7:0]  io_pipe_phv_in_data_349,
  input  [7:0]  io_pipe_phv_in_data_350,
  input  [7:0]  io_pipe_phv_in_data_351,
  input  [7:0]  io_pipe_phv_in_data_352,
  input  [7:0]  io_pipe_phv_in_data_353,
  input  [7:0]  io_pipe_phv_in_data_354,
  input  [7:0]  io_pipe_phv_in_data_355,
  input  [7:0]  io_pipe_phv_in_data_356,
  input  [7:0]  io_pipe_phv_in_data_357,
  input  [7:0]  io_pipe_phv_in_data_358,
  input  [7:0]  io_pipe_phv_in_data_359,
  input  [7:0]  io_pipe_phv_in_data_360,
  input  [7:0]  io_pipe_phv_in_data_361,
  input  [7:0]  io_pipe_phv_in_data_362,
  input  [7:0]  io_pipe_phv_in_data_363,
  input  [7:0]  io_pipe_phv_in_data_364,
  input  [7:0]  io_pipe_phv_in_data_365,
  input  [7:0]  io_pipe_phv_in_data_366,
  input  [7:0]  io_pipe_phv_in_data_367,
  input  [7:0]  io_pipe_phv_in_data_368,
  input  [7:0]  io_pipe_phv_in_data_369,
  input  [7:0]  io_pipe_phv_in_data_370,
  input  [7:0]  io_pipe_phv_in_data_371,
  input  [7:0]  io_pipe_phv_in_data_372,
  input  [7:0]  io_pipe_phv_in_data_373,
  input  [7:0]  io_pipe_phv_in_data_374,
  input  [7:0]  io_pipe_phv_in_data_375,
  input  [7:0]  io_pipe_phv_in_data_376,
  input  [7:0]  io_pipe_phv_in_data_377,
  input  [7:0]  io_pipe_phv_in_data_378,
  input  [7:0]  io_pipe_phv_in_data_379,
  input  [7:0]  io_pipe_phv_in_data_380,
  input  [7:0]  io_pipe_phv_in_data_381,
  input  [7:0]  io_pipe_phv_in_data_382,
  input  [7:0]  io_pipe_phv_in_data_383,
  input  [7:0]  io_pipe_phv_in_data_384,
  input  [7:0]  io_pipe_phv_in_data_385,
  input  [7:0]  io_pipe_phv_in_data_386,
  input  [7:0]  io_pipe_phv_in_data_387,
  input  [7:0]  io_pipe_phv_in_data_388,
  input  [7:0]  io_pipe_phv_in_data_389,
  input  [7:0]  io_pipe_phv_in_data_390,
  input  [7:0]  io_pipe_phv_in_data_391,
  input  [7:0]  io_pipe_phv_in_data_392,
  input  [7:0]  io_pipe_phv_in_data_393,
  input  [7:0]  io_pipe_phv_in_data_394,
  input  [7:0]  io_pipe_phv_in_data_395,
  input  [7:0]  io_pipe_phv_in_data_396,
  input  [7:0]  io_pipe_phv_in_data_397,
  input  [7:0]  io_pipe_phv_in_data_398,
  input  [7:0]  io_pipe_phv_in_data_399,
  input  [7:0]  io_pipe_phv_in_data_400,
  input  [7:0]  io_pipe_phv_in_data_401,
  input  [7:0]  io_pipe_phv_in_data_402,
  input  [7:0]  io_pipe_phv_in_data_403,
  input  [7:0]  io_pipe_phv_in_data_404,
  input  [7:0]  io_pipe_phv_in_data_405,
  input  [7:0]  io_pipe_phv_in_data_406,
  input  [7:0]  io_pipe_phv_in_data_407,
  input  [7:0]  io_pipe_phv_in_data_408,
  input  [7:0]  io_pipe_phv_in_data_409,
  input  [7:0]  io_pipe_phv_in_data_410,
  input  [7:0]  io_pipe_phv_in_data_411,
  input  [7:0]  io_pipe_phv_in_data_412,
  input  [7:0]  io_pipe_phv_in_data_413,
  input  [7:0]  io_pipe_phv_in_data_414,
  input  [7:0]  io_pipe_phv_in_data_415,
  input  [7:0]  io_pipe_phv_in_data_416,
  input  [7:0]  io_pipe_phv_in_data_417,
  input  [7:0]  io_pipe_phv_in_data_418,
  input  [7:0]  io_pipe_phv_in_data_419,
  input  [7:0]  io_pipe_phv_in_data_420,
  input  [7:0]  io_pipe_phv_in_data_421,
  input  [7:0]  io_pipe_phv_in_data_422,
  input  [7:0]  io_pipe_phv_in_data_423,
  input  [7:0]  io_pipe_phv_in_data_424,
  input  [7:0]  io_pipe_phv_in_data_425,
  input  [7:0]  io_pipe_phv_in_data_426,
  input  [7:0]  io_pipe_phv_in_data_427,
  input  [7:0]  io_pipe_phv_in_data_428,
  input  [7:0]  io_pipe_phv_in_data_429,
  input  [7:0]  io_pipe_phv_in_data_430,
  input  [7:0]  io_pipe_phv_in_data_431,
  input  [7:0]  io_pipe_phv_in_data_432,
  input  [7:0]  io_pipe_phv_in_data_433,
  input  [7:0]  io_pipe_phv_in_data_434,
  input  [7:0]  io_pipe_phv_in_data_435,
  input  [7:0]  io_pipe_phv_in_data_436,
  input  [7:0]  io_pipe_phv_in_data_437,
  input  [7:0]  io_pipe_phv_in_data_438,
  input  [7:0]  io_pipe_phv_in_data_439,
  input  [7:0]  io_pipe_phv_in_data_440,
  input  [7:0]  io_pipe_phv_in_data_441,
  input  [7:0]  io_pipe_phv_in_data_442,
  input  [7:0]  io_pipe_phv_in_data_443,
  input  [7:0]  io_pipe_phv_in_data_444,
  input  [7:0]  io_pipe_phv_in_data_445,
  input  [7:0]  io_pipe_phv_in_data_446,
  input  [7:0]  io_pipe_phv_in_data_447,
  input  [7:0]  io_pipe_phv_in_data_448,
  input  [7:0]  io_pipe_phv_in_data_449,
  input  [7:0]  io_pipe_phv_in_data_450,
  input  [7:0]  io_pipe_phv_in_data_451,
  input  [7:0]  io_pipe_phv_in_data_452,
  input  [7:0]  io_pipe_phv_in_data_453,
  input  [7:0]  io_pipe_phv_in_data_454,
  input  [7:0]  io_pipe_phv_in_data_455,
  input  [7:0]  io_pipe_phv_in_data_456,
  input  [7:0]  io_pipe_phv_in_data_457,
  input  [7:0]  io_pipe_phv_in_data_458,
  input  [7:0]  io_pipe_phv_in_data_459,
  input  [7:0]  io_pipe_phv_in_data_460,
  input  [7:0]  io_pipe_phv_in_data_461,
  input  [7:0]  io_pipe_phv_in_data_462,
  input  [7:0]  io_pipe_phv_in_data_463,
  input  [7:0]  io_pipe_phv_in_data_464,
  input  [7:0]  io_pipe_phv_in_data_465,
  input  [7:0]  io_pipe_phv_in_data_466,
  input  [7:0]  io_pipe_phv_in_data_467,
  input  [7:0]  io_pipe_phv_in_data_468,
  input  [7:0]  io_pipe_phv_in_data_469,
  input  [7:0]  io_pipe_phv_in_data_470,
  input  [7:0]  io_pipe_phv_in_data_471,
  input  [7:0]  io_pipe_phv_in_data_472,
  input  [7:0]  io_pipe_phv_in_data_473,
  input  [7:0]  io_pipe_phv_in_data_474,
  input  [7:0]  io_pipe_phv_in_data_475,
  input  [7:0]  io_pipe_phv_in_data_476,
  input  [7:0]  io_pipe_phv_in_data_477,
  input  [7:0]  io_pipe_phv_in_data_478,
  input  [7:0]  io_pipe_phv_in_data_479,
  input  [7:0]  io_pipe_phv_in_data_480,
  input  [7:0]  io_pipe_phv_in_data_481,
  input  [7:0]  io_pipe_phv_in_data_482,
  input  [7:0]  io_pipe_phv_in_data_483,
  input  [7:0]  io_pipe_phv_in_data_484,
  input  [7:0]  io_pipe_phv_in_data_485,
  input  [7:0]  io_pipe_phv_in_data_486,
  input  [7:0]  io_pipe_phv_in_data_487,
  input  [7:0]  io_pipe_phv_in_data_488,
  input  [7:0]  io_pipe_phv_in_data_489,
  input  [7:0]  io_pipe_phv_in_data_490,
  input  [7:0]  io_pipe_phv_in_data_491,
  input  [7:0]  io_pipe_phv_in_data_492,
  input  [7:0]  io_pipe_phv_in_data_493,
  input  [7:0]  io_pipe_phv_in_data_494,
  input  [7:0]  io_pipe_phv_in_data_495,
  input  [7:0]  io_pipe_phv_in_data_496,
  input  [7:0]  io_pipe_phv_in_data_497,
  input  [7:0]  io_pipe_phv_in_data_498,
  input  [7:0]  io_pipe_phv_in_data_499,
  input  [7:0]  io_pipe_phv_in_data_500,
  input  [7:0]  io_pipe_phv_in_data_501,
  input  [7:0]  io_pipe_phv_in_data_502,
  input  [7:0]  io_pipe_phv_in_data_503,
  input  [7:0]  io_pipe_phv_in_data_504,
  input  [7:0]  io_pipe_phv_in_data_505,
  input  [7:0]  io_pipe_phv_in_data_506,
  input  [7:0]  io_pipe_phv_in_data_507,
  input  [7:0]  io_pipe_phv_in_data_508,
  input  [7:0]  io_pipe_phv_in_data_509,
  input  [7:0]  io_pipe_phv_in_data_510,
  input  [7:0]  io_pipe_phv_in_data_511,
  input  [3:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [7:0]  io_pipe_phv_out_data_160,
  output [7:0]  io_pipe_phv_out_data_161,
  output [7:0]  io_pipe_phv_out_data_162,
  output [7:0]  io_pipe_phv_out_data_163,
  output [7:0]  io_pipe_phv_out_data_164,
  output [7:0]  io_pipe_phv_out_data_165,
  output [7:0]  io_pipe_phv_out_data_166,
  output [7:0]  io_pipe_phv_out_data_167,
  output [7:0]  io_pipe_phv_out_data_168,
  output [7:0]  io_pipe_phv_out_data_169,
  output [7:0]  io_pipe_phv_out_data_170,
  output [7:0]  io_pipe_phv_out_data_171,
  output [7:0]  io_pipe_phv_out_data_172,
  output [7:0]  io_pipe_phv_out_data_173,
  output [7:0]  io_pipe_phv_out_data_174,
  output [7:0]  io_pipe_phv_out_data_175,
  output [7:0]  io_pipe_phv_out_data_176,
  output [7:0]  io_pipe_phv_out_data_177,
  output [7:0]  io_pipe_phv_out_data_178,
  output [7:0]  io_pipe_phv_out_data_179,
  output [7:0]  io_pipe_phv_out_data_180,
  output [7:0]  io_pipe_phv_out_data_181,
  output [7:0]  io_pipe_phv_out_data_182,
  output [7:0]  io_pipe_phv_out_data_183,
  output [7:0]  io_pipe_phv_out_data_184,
  output [7:0]  io_pipe_phv_out_data_185,
  output [7:0]  io_pipe_phv_out_data_186,
  output [7:0]  io_pipe_phv_out_data_187,
  output [7:0]  io_pipe_phv_out_data_188,
  output [7:0]  io_pipe_phv_out_data_189,
  output [7:0]  io_pipe_phv_out_data_190,
  output [7:0]  io_pipe_phv_out_data_191,
  output [7:0]  io_pipe_phv_out_data_192,
  output [7:0]  io_pipe_phv_out_data_193,
  output [7:0]  io_pipe_phv_out_data_194,
  output [7:0]  io_pipe_phv_out_data_195,
  output [7:0]  io_pipe_phv_out_data_196,
  output [7:0]  io_pipe_phv_out_data_197,
  output [7:0]  io_pipe_phv_out_data_198,
  output [7:0]  io_pipe_phv_out_data_199,
  output [7:0]  io_pipe_phv_out_data_200,
  output [7:0]  io_pipe_phv_out_data_201,
  output [7:0]  io_pipe_phv_out_data_202,
  output [7:0]  io_pipe_phv_out_data_203,
  output [7:0]  io_pipe_phv_out_data_204,
  output [7:0]  io_pipe_phv_out_data_205,
  output [7:0]  io_pipe_phv_out_data_206,
  output [7:0]  io_pipe_phv_out_data_207,
  output [7:0]  io_pipe_phv_out_data_208,
  output [7:0]  io_pipe_phv_out_data_209,
  output [7:0]  io_pipe_phv_out_data_210,
  output [7:0]  io_pipe_phv_out_data_211,
  output [7:0]  io_pipe_phv_out_data_212,
  output [7:0]  io_pipe_phv_out_data_213,
  output [7:0]  io_pipe_phv_out_data_214,
  output [7:0]  io_pipe_phv_out_data_215,
  output [7:0]  io_pipe_phv_out_data_216,
  output [7:0]  io_pipe_phv_out_data_217,
  output [7:0]  io_pipe_phv_out_data_218,
  output [7:0]  io_pipe_phv_out_data_219,
  output [7:0]  io_pipe_phv_out_data_220,
  output [7:0]  io_pipe_phv_out_data_221,
  output [7:0]  io_pipe_phv_out_data_222,
  output [7:0]  io_pipe_phv_out_data_223,
  output [7:0]  io_pipe_phv_out_data_224,
  output [7:0]  io_pipe_phv_out_data_225,
  output [7:0]  io_pipe_phv_out_data_226,
  output [7:0]  io_pipe_phv_out_data_227,
  output [7:0]  io_pipe_phv_out_data_228,
  output [7:0]  io_pipe_phv_out_data_229,
  output [7:0]  io_pipe_phv_out_data_230,
  output [7:0]  io_pipe_phv_out_data_231,
  output [7:0]  io_pipe_phv_out_data_232,
  output [7:0]  io_pipe_phv_out_data_233,
  output [7:0]  io_pipe_phv_out_data_234,
  output [7:0]  io_pipe_phv_out_data_235,
  output [7:0]  io_pipe_phv_out_data_236,
  output [7:0]  io_pipe_phv_out_data_237,
  output [7:0]  io_pipe_phv_out_data_238,
  output [7:0]  io_pipe_phv_out_data_239,
  output [7:0]  io_pipe_phv_out_data_240,
  output [7:0]  io_pipe_phv_out_data_241,
  output [7:0]  io_pipe_phv_out_data_242,
  output [7:0]  io_pipe_phv_out_data_243,
  output [7:0]  io_pipe_phv_out_data_244,
  output [7:0]  io_pipe_phv_out_data_245,
  output [7:0]  io_pipe_phv_out_data_246,
  output [7:0]  io_pipe_phv_out_data_247,
  output [7:0]  io_pipe_phv_out_data_248,
  output [7:0]  io_pipe_phv_out_data_249,
  output [7:0]  io_pipe_phv_out_data_250,
  output [7:0]  io_pipe_phv_out_data_251,
  output [7:0]  io_pipe_phv_out_data_252,
  output [7:0]  io_pipe_phv_out_data_253,
  output [7:0]  io_pipe_phv_out_data_254,
  output [7:0]  io_pipe_phv_out_data_255,
  output [7:0]  io_pipe_phv_out_data_256,
  output [7:0]  io_pipe_phv_out_data_257,
  output [7:0]  io_pipe_phv_out_data_258,
  output [7:0]  io_pipe_phv_out_data_259,
  output [7:0]  io_pipe_phv_out_data_260,
  output [7:0]  io_pipe_phv_out_data_261,
  output [7:0]  io_pipe_phv_out_data_262,
  output [7:0]  io_pipe_phv_out_data_263,
  output [7:0]  io_pipe_phv_out_data_264,
  output [7:0]  io_pipe_phv_out_data_265,
  output [7:0]  io_pipe_phv_out_data_266,
  output [7:0]  io_pipe_phv_out_data_267,
  output [7:0]  io_pipe_phv_out_data_268,
  output [7:0]  io_pipe_phv_out_data_269,
  output [7:0]  io_pipe_phv_out_data_270,
  output [7:0]  io_pipe_phv_out_data_271,
  output [7:0]  io_pipe_phv_out_data_272,
  output [7:0]  io_pipe_phv_out_data_273,
  output [7:0]  io_pipe_phv_out_data_274,
  output [7:0]  io_pipe_phv_out_data_275,
  output [7:0]  io_pipe_phv_out_data_276,
  output [7:0]  io_pipe_phv_out_data_277,
  output [7:0]  io_pipe_phv_out_data_278,
  output [7:0]  io_pipe_phv_out_data_279,
  output [7:0]  io_pipe_phv_out_data_280,
  output [7:0]  io_pipe_phv_out_data_281,
  output [7:0]  io_pipe_phv_out_data_282,
  output [7:0]  io_pipe_phv_out_data_283,
  output [7:0]  io_pipe_phv_out_data_284,
  output [7:0]  io_pipe_phv_out_data_285,
  output [7:0]  io_pipe_phv_out_data_286,
  output [7:0]  io_pipe_phv_out_data_287,
  output [7:0]  io_pipe_phv_out_data_288,
  output [7:0]  io_pipe_phv_out_data_289,
  output [7:0]  io_pipe_phv_out_data_290,
  output [7:0]  io_pipe_phv_out_data_291,
  output [7:0]  io_pipe_phv_out_data_292,
  output [7:0]  io_pipe_phv_out_data_293,
  output [7:0]  io_pipe_phv_out_data_294,
  output [7:0]  io_pipe_phv_out_data_295,
  output [7:0]  io_pipe_phv_out_data_296,
  output [7:0]  io_pipe_phv_out_data_297,
  output [7:0]  io_pipe_phv_out_data_298,
  output [7:0]  io_pipe_phv_out_data_299,
  output [7:0]  io_pipe_phv_out_data_300,
  output [7:0]  io_pipe_phv_out_data_301,
  output [7:0]  io_pipe_phv_out_data_302,
  output [7:0]  io_pipe_phv_out_data_303,
  output [7:0]  io_pipe_phv_out_data_304,
  output [7:0]  io_pipe_phv_out_data_305,
  output [7:0]  io_pipe_phv_out_data_306,
  output [7:0]  io_pipe_phv_out_data_307,
  output [7:0]  io_pipe_phv_out_data_308,
  output [7:0]  io_pipe_phv_out_data_309,
  output [7:0]  io_pipe_phv_out_data_310,
  output [7:0]  io_pipe_phv_out_data_311,
  output [7:0]  io_pipe_phv_out_data_312,
  output [7:0]  io_pipe_phv_out_data_313,
  output [7:0]  io_pipe_phv_out_data_314,
  output [7:0]  io_pipe_phv_out_data_315,
  output [7:0]  io_pipe_phv_out_data_316,
  output [7:0]  io_pipe_phv_out_data_317,
  output [7:0]  io_pipe_phv_out_data_318,
  output [7:0]  io_pipe_phv_out_data_319,
  output [7:0]  io_pipe_phv_out_data_320,
  output [7:0]  io_pipe_phv_out_data_321,
  output [7:0]  io_pipe_phv_out_data_322,
  output [7:0]  io_pipe_phv_out_data_323,
  output [7:0]  io_pipe_phv_out_data_324,
  output [7:0]  io_pipe_phv_out_data_325,
  output [7:0]  io_pipe_phv_out_data_326,
  output [7:0]  io_pipe_phv_out_data_327,
  output [7:0]  io_pipe_phv_out_data_328,
  output [7:0]  io_pipe_phv_out_data_329,
  output [7:0]  io_pipe_phv_out_data_330,
  output [7:0]  io_pipe_phv_out_data_331,
  output [7:0]  io_pipe_phv_out_data_332,
  output [7:0]  io_pipe_phv_out_data_333,
  output [7:0]  io_pipe_phv_out_data_334,
  output [7:0]  io_pipe_phv_out_data_335,
  output [7:0]  io_pipe_phv_out_data_336,
  output [7:0]  io_pipe_phv_out_data_337,
  output [7:0]  io_pipe_phv_out_data_338,
  output [7:0]  io_pipe_phv_out_data_339,
  output [7:0]  io_pipe_phv_out_data_340,
  output [7:0]  io_pipe_phv_out_data_341,
  output [7:0]  io_pipe_phv_out_data_342,
  output [7:0]  io_pipe_phv_out_data_343,
  output [7:0]  io_pipe_phv_out_data_344,
  output [7:0]  io_pipe_phv_out_data_345,
  output [7:0]  io_pipe_phv_out_data_346,
  output [7:0]  io_pipe_phv_out_data_347,
  output [7:0]  io_pipe_phv_out_data_348,
  output [7:0]  io_pipe_phv_out_data_349,
  output [7:0]  io_pipe_phv_out_data_350,
  output [7:0]  io_pipe_phv_out_data_351,
  output [7:0]  io_pipe_phv_out_data_352,
  output [7:0]  io_pipe_phv_out_data_353,
  output [7:0]  io_pipe_phv_out_data_354,
  output [7:0]  io_pipe_phv_out_data_355,
  output [7:0]  io_pipe_phv_out_data_356,
  output [7:0]  io_pipe_phv_out_data_357,
  output [7:0]  io_pipe_phv_out_data_358,
  output [7:0]  io_pipe_phv_out_data_359,
  output [7:0]  io_pipe_phv_out_data_360,
  output [7:0]  io_pipe_phv_out_data_361,
  output [7:0]  io_pipe_phv_out_data_362,
  output [7:0]  io_pipe_phv_out_data_363,
  output [7:0]  io_pipe_phv_out_data_364,
  output [7:0]  io_pipe_phv_out_data_365,
  output [7:0]  io_pipe_phv_out_data_366,
  output [7:0]  io_pipe_phv_out_data_367,
  output [7:0]  io_pipe_phv_out_data_368,
  output [7:0]  io_pipe_phv_out_data_369,
  output [7:0]  io_pipe_phv_out_data_370,
  output [7:0]  io_pipe_phv_out_data_371,
  output [7:0]  io_pipe_phv_out_data_372,
  output [7:0]  io_pipe_phv_out_data_373,
  output [7:0]  io_pipe_phv_out_data_374,
  output [7:0]  io_pipe_phv_out_data_375,
  output [7:0]  io_pipe_phv_out_data_376,
  output [7:0]  io_pipe_phv_out_data_377,
  output [7:0]  io_pipe_phv_out_data_378,
  output [7:0]  io_pipe_phv_out_data_379,
  output [7:0]  io_pipe_phv_out_data_380,
  output [7:0]  io_pipe_phv_out_data_381,
  output [7:0]  io_pipe_phv_out_data_382,
  output [7:0]  io_pipe_phv_out_data_383,
  output [7:0]  io_pipe_phv_out_data_384,
  output [7:0]  io_pipe_phv_out_data_385,
  output [7:0]  io_pipe_phv_out_data_386,
  output [7:0]  io_pipe_phv_out_data_387,
  output [7:0]  io_pipe_phv_out_data_388,
  output [7:0]  io_pipe_phv_out_data_389,
  output [7:0]  io_pipe_phv_out_data_390,
  output [7:0]  io_pipe_phv_out_data_391,
  output [7:0]  io_pipe_phv_out_data_392,
  output [7:0]  io_pipe_phv_out_data_393,
  output [7:0]  io_pipe_phv_out_data_394,
  output [7:0]  io_pipe_phv_out_data_395,
  output [7:0]  io_pipe_phv_out_data_396,
  output [7:0]  io_pipe_phv_out_data_397,
  output [7:0]  io_pipe_phv_out_data_398,
  output [7:0]  io_pipe_phv_out_data_399,
  output [7:0]  io_pipe_phv_out_data_400,
  output [7:0]  io_pipe_phv_out_data_401,
  output [7:0]  io_pipe_phv_out_data_402,
  output [7:0]  io_pipe_phv_out_data_403,
  output [7:0]  io_pipe_phv_out_data_404,
  output [7:0]  io_pipe_phv_out_data_405,
  output [7:0]  io_pipe_phv_out_data_406,
  output [7:0]  io_pipe_phv_out_data_407,
  output [7:0]  io_pipe_phv_out_data_408,
  output [7:0]  io_pipe_phv_out_data_409,
  output [7:0]  io_pipe_phv_out_data_410,
  output [7:0]  io_pipe_phv_out_data_411,
  output [7:0]  io_pipe_phv_out_data_412,
  output [7:0]  io_pipe_phv_out_data_413,
  output [7:0]  io_pipe_phv_out_data_414,
  output [7:0]  io_pipe_phv_out_data_415,
  output [7:0]  io_pipe_phv_out_data_416,
  output [7:0]  io_pipe_phv_out_data_417,
  output [7:0]  io_pipe_phv_out_data_418,
  output [7:0]  io_pipe_phv_out_data_419,
  output [7:0]  io_pipe_phv_out_data_420,
  output [7:0]  io_pipe_phv_out_data_421,
  output [7:0]  io_pipe_phv_out_data_422,
  output [7:0]  io_pipe_phv_out_data_423,
  output [7:0]  io_pipe_phv_out_data_424,
  output [7:0]  io_pipe_phv_out_data_425,
  output [7:0]  io_pipe_phv_out_data_426,
  output [7:0]  io_pipe_phv_out_data_427,
  output [7:0]  io_pipe_phv_out_data_428,
  output [7:0]  io_pipe_phv_out_data_429,
  output [7:0]  io_pipe_phv_out_data_430,
  output [7:0]  io_pipe_phv_out_data_431,
  output [7:0]  io_pipe_phv_out_data_432,
  output [7:0]  io_pipe_phv_out_data_433,
  output [7:0]  io_pipe_phv_out_data_434,
  output [7:0]  io_pipe_phv_out_data_435,
  output [7:0]  io_pipe_phv_out_data_436,
  output [7:0]  io_pipe_phv_out_data_437,
  output [7:0]  io_pipe_phv_out_data_438,
  output [7:0]  io_pipe_phv_out_data_439,
  output [7:0]  io_pipe_phv_out_data_440,
  output [7:0]  io_pipe_phv_out_data_441,
  output [7:0]  io_pipe_phv_out_data_442,
  output [7:0]  io_pipe_phv_out_data_443,
  output [7:0]  io_pipe_phv_out_data_444,
  output [7:0]  io_pipe_phv_out_data_445,
  output [7:0]  io_pipe_phv_out_data_446,
  output [7:0]  io_pipe_phv_out_data_447,
  output [7:0]  io_pipe_phv_out_data_448,
  output [7:0]  io_pipe_phv_out_data_449,
  output [7:0]  io_pipe_phv_out_data_450,
  output [7:0]  io_pipe_phv_out_data_451,
  output [7:0]  io_pipe_phv_out_data_452,
  output [7:0]  io_pipe_phv_out_data_453,
  output [7:0]  io_pipe_phv_out_data_454,
  output [7:0]  io_pipe_phv_out_data_455,
  output [7:0]  io_pipe_phv_out_data_456,
  output [7:0]  io_pipe_phv_out_data_457,
  output [7:0]  io_pipe_phv_out_data_458,
  output [7:0]  io_pipe_phv_out_data_459,
  output [7:0]  io_pipe_phv_out_data_460,
  output [7:0]  io_pipe_phv_out_data_461,
  output [7:0]  io_pipe_phv_out_data_462,
  output [7:0]  io_pipe_phv_out_data_463,
  output [7:0]  io_pipe_phv_out_data_464,
  output [7:0]  io_pipe_phv_out_data_465,
  output [7:0]  io_pipe_phv_out_data_466,
  output [7:0]  io_pipe_phv_out_data_467,
  output [7:0]  io_pipe_phv_out_data_468,
  output [7:0]  io_pipe_phv_out_data_469,
  output [7:0]  io_pipe_phv_out_data_470,
  output [7:0]  io_pipe_phv_out_data_471,
  output [7:0]  io_pipe_phv_out_data_472,
  output [7:0]  io_pipe_phv_out_data_473,
  output [7:0]  io_pipe_phv_out_data_474,
  output [7:0]  io_pipe_phv_out_data_475,
  output [7:0]  io_pipe_phv_out_data_476,
  output [7:0]  io_pipe_phv_out_data_477,
  output [7:0]  io_pipe_phv_out_data_478,
  output [7:0]  io_pipe_phv_out_data_479,
  output [7:0]  io_pipe_phv_out_data_480,
  output [7:0]  io_pipe_phv_out_data_481,
  output [7:0]  io_pipe_phv_out_data_482,
  output [7:0]  io_pipe_phv_out_data_483,
  output [7:0]  io_pipe_phv_out_data_484,
  output [7:0]  io_pipe_phv_out_data_485,
  output [7:0]  io_pipe_phv_out_data_486,
  output [7:0]  io_pipe_phv_out_data_487,
  output [7:0]  io_pipe_phv_out_data_488,
  output [7:0]  io_pipe_phv_out_data_489,
  output [7:0]  io_pipe_phv_out_data_490,
  output [7:0]  io_pipe_phv_out_data_491,
  output [7:0]  io_pipe_phv_out_data_492,
  output [7:0]  io_pipe_phv_out_data_493,
  output [7:0]  io_pipe_phv_out_data_494,
  output [7:0]  io_pipe_phv_out_data_495,
  output [7:0]  io_pipe_phv_out_data_496,
  output [7:0]  io_pipe_phv_out_data_497,
  output [7:0]  io_pipe_phv_out_data_498,
  output [7:0]  io_pipe_phv_out_data_499,
  output [7:0]  io_pipe_phv_out_data_500,
  output [7:0]  io_pipe_phv_out_data_501,
  output [7:0]  io_pipe_phv_out_data_502,
  output [7:0]  io_pipe_phv_out_data_503,
  output [7:0]  io_pipe_phv_out_data_504,
  output [7:0]  io_pipe_phv_out_data_505,
  output [7:0]  io_pipe_phv_out_data_506,
  output [7:0]  io_pipe_phv_out_data_507,
  output [7:0]  io_pipe_phv_out_data_508,
  output [7:0]  io_pipe_phv_out_data_509,
  output [7:0]  io_pipe_phv_out_data_510,
  output [7:0]  io_pipe_phv_out_data_511,
  output [3:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input         io_mod_en,
  input         io_mod_config_id,
  input         io_mod_key_mod_en,
  input  [2:0]  io_mod_key_mod_group_index,
  input  [1:0]  io_mod_key_mod_group_config,
  input         io_mod_key_mod_group_mask_0,
  input         io_mod_key_mod_group_mask_1,
  input         io_mod_key_mod_group_mask_2,
  input         io_mod_key_mod_group_mask_3,
  input  [7:0]  io_mod_key_mod_group_id_0,
  input  [7:0]  io_mod_key_mod_group_id_1,
  input  [7:0]  io_mod_key_mod_group_id_2,
  input  [7:0]  io_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_table_mod_table_depth,
  input  [4:0]  io_mod_table_mod_table_width,
  input         io_mod_w_en,
  input  [3:0]  io_mod_w_sram_id,
  input  [7:0]  io_mod_w_addr,
  input  [63:0] io_mod_w_data,
  output        io_hit,
  output [63:0] io_match_value
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
`endif // RANDOMIZE_REG_INIT
  wire  pipe1_clock; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_4; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_5; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_6; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_7; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_8; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_9; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_10; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_11; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_12; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_13; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_14; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_15; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_16; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_17; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_18; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_19; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_20; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_21; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_22; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_23; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_24; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_25; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_26; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_27; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_28; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_29; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_30; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_31; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_32; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_33; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_34; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_35; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_36; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_37; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_38; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_39; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_40; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_41; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_42; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_43; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_44; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_45; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_46; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_47; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_48; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_49; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_50; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_51; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_52; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_53; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_54; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_55; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_56; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_57; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_58; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_59; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_60; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_61; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_62; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_63; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_64; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_65; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_66; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_67; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_68; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_69; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_70; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_71; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_72; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_73; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_74; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_75; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_76; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_77; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_78; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_79; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_80; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_81; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_82; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_83; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_84; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_85; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_86; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_87; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_88; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_89; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_90; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_91; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_92; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_93; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_94; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_95; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_96; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_97; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_98; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_99; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_100; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_101; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_102; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_103; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_104; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_105; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_106; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_107; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_108; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_109; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_110; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_111; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_112; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_113; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_114; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_115; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_116; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_117; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_118; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_119; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_120; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_121; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_122; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_123; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_124; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_125; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_126; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_127; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_128; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_129; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_130; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_131; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_132; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_133; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_134; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_135; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_136; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_137; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_138; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_139; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_140; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_141; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_142; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_143; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_144; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_145; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_146; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_147; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_148; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_149; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_150; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_151; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_152; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_153; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_154; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_155; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_156; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_157; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_158; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_159; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_160; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_161; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_162; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_163; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_164; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_165; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_166; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_167; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_168; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_169; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_170; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_171; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_172; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_173; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_174; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_175; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_176; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_177; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_178; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_179; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_180; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_181; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_182; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_183; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_184; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_185; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_186; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_187; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_188; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_189; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_190; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_191; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_192; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_193; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_194; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_195; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_196; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_197; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_198; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_199; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_200; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_201; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_202; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_203; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_204; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_205; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_206; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_207; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_208; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_209; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_210; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_211; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_212; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_213; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_214; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_215; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_216; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_217; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_218; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_219; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_220; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_221; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_222; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_223; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_224; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_225; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_226; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_227; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_228; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_229; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_230; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_231; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_232; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_233; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_234; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_235; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_236; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_237; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_238; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_239; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_240; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_241; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_242; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_243; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_244; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_245; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_246; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_247; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_248; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_249; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_250; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_251; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_252; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_253; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_254; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_255; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_256; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_257; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_258; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_259; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_260; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_261; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_262; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_263; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_264; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_265; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_266; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_267; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_268; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_269; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_270; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_271; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_272; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_273; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_274; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_275; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_276; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_277; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_278; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_279; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_280; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_281; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_282; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_283; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_284; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_285; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_286; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_287; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_288; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_289; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_290; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_291; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_292; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_293; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_294; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_295; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_296; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_297; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_298; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_299; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_300; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_301; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_302; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_303; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_304; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_305; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_306; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_307; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_308; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_309; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_310; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_311; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_312; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_313; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_314; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_315; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_316; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_317; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_318; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_319; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_320; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_321; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_322; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_323; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_324; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_325; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_326; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_327; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_328; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_329; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_330; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_331; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_332; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_333; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_334; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_335; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_336; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_337; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_338; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_339; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_340; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_341; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_342; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_343; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_344; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_345; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_346; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_347; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_348; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_349; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_350; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_351; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_352; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_353; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_354; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_355; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_356; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_357; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_358; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_359; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_360; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_361; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_362; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_363; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_364; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_365; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_366; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_367; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_368; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_369; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_370; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_371; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_372; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_373; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_374; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_375; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_376; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_377; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_378; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_379; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_380; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_381; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_382; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_383; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_384; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_385; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_386; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_387; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_388; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_389; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_390; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_391; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_392; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_393; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_394; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_395; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_396; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_397; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_398; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_399; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_400; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_401; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_402; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_403; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_404; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_405; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_406; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_407; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_408; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_409; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_410; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_411; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_412; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_413; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_414; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_415; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_416; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_417; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_418; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_419; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_420; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_421; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_422; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_423; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_424; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_425; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_426; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_427; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_428; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_429; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_430; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_431; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_432; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_433; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_434; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_435; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_436; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_437; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_438; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_439; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_440; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_441; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_442; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_443; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_444; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_445; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_446; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_447; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_448; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_449; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_450; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_451; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_452; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_453; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_454; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_455; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_456; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_457; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_458; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_459; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_460; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_461; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_462; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_463; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_464; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_465; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_466; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_467; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_468; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_469; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_470; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_471; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_472; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_473; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_474; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_475; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_476; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_477; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_478; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_479; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_480; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_481; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_482; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_483; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_484; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_485; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_486; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_487; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_488; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_489; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_490; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_491; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_492; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_493; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_494; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_495; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_496; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_497; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_498; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_499; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_500; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_501; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_502; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_503; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_504; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_505; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_506; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_507; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_508; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_509; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_510; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_511; // @[matcher_pisa.scala 333:23]
  wire [3:0] pipe1_io_pipe_phv_in_next_processor_id; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_pipe_phv_in_next_config_id; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_pipe_phv_in_is_valid_processor; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_4; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_5; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_6; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_7; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_8; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_9; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_10; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_11; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_12; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_13; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_14; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_15; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_16; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_17; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_18; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_19; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_20; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_21; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_22; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_23; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_24; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_25; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_26; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_27; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_28; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_29; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_30; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_31; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_32; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_33; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_34; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_35; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_36; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_37; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_38; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_39; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_40; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_41; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_42; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_43; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_44; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_45; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_46; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_47; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_48; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_49; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_50; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_51; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_52; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_53; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_54; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_55; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_56; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_57; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_58; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_59; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_60; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_61; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_62; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_63; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_64; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_65; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_66; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_67; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_68; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_69; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_70; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_71; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_72; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_73; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_74; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_75; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_76; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_77; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_78; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_79; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_80; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_81; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_82; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_83; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_84; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_85; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_86; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_87; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_88; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_89; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_90; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_91; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_92; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_93; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_94; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_95; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_96; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_97; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_98; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_99; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_100; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_101; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_102; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_103; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_104; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_105; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_106; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_107; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_108; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_109; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_110; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_111; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_112; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_113; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_114; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_115; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_116; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_117; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_118; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_119; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_120; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_121; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_122; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_123; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_124; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_125; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_126; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_127; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_128; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_129; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_130; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_131; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_132; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_133; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_134; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_135; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_136; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_137; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_138; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_139; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_140; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_141; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_142; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_143; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_144; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_145; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_146; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_147; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_148; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_149; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_150; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_151; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_152; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_153; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_154; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_155; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_156; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_157; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_158; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_159; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_160; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_161; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_162; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_163; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_164; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_165; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_166; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_167; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_168; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_169; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_170; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_171; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_172; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_173; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_174; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_175; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_176; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_177; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_178; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_179; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_180; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_181; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_182; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_183; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_184; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_185; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_186; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_187; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_188; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_189; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_190; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_191; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_192; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_193; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_194; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_195; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_196; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_197; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_198; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_199; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_200; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_201; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_202; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_203; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_204; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_205; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_206; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_207; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_208; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_209; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_210; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_211; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_212; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_213; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_214; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_215; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_216; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_217; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_218; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_219; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_220; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_221; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_222; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_223; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_224; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_225; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_226; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_227; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_228; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_229; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_230; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_231; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_232; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_233; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_234; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_235; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_236; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_237; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_238; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_239; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_240; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_241; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_242; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_243; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_244; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_245; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_246; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_247; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_248; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_249; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_250; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_251; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_252; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_253; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_254; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_255; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_256; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_257; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_258; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_259; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_260; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_261; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_262; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_263; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_264; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_265; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_266; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_267; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_268; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_269; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_270; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_271; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_272; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_273; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_274; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_275; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_276; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_277; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_278; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_279; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_280; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_281; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_282; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_283; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_284; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_285; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_286; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_287; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_288; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_289; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_290; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_291; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_292; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_293; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_294; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_295; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_296; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_297; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_298; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_299; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_300; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_301; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_302; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_303; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_304; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_305; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_306; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_307; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_308; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_309; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_310; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_311; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_312; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_313; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_314; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_315; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_316; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_317; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_318; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_319; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_320; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_321; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_322; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_323; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_324; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_325; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_326; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_327; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_328; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_329; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_330; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_331; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_332; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_333; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_334; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_335; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_336; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_337; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_338; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_339; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_340; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_341; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_342; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_343; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_344; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_345; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_346; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_347; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_348; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_349; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_350; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_351; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_352; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_353; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_354; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_355; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_356; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_357; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_358; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_359; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_360; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_361; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_362; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_363; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_364; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_365; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_366; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_367; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_368; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_369; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_370; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_371; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_372; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_373; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_374; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_375; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_376; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_377; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_378; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_379; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_380; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_381; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_382; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_383; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_384; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_385; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_386; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_387; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_388; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_389; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_390; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_391; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_392; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_393; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_394; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_395; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_396; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_397; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_398; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_399; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_400; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_401; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_402; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_403; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_404; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_405; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_406; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_407; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_408; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_409; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_410; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_411; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_412; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_413; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_414; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_415; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_416; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_417; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_418; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_419; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_420; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_421; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_422; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_423; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_424; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_425; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_426; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_427; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_428; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_429; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_430; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_431; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_432; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_433; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_434; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_435; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_436; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_437; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_438; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_439; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_440; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_441; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_442; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_443; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_444; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_445; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_446; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_447; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_448; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_449; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_450; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_451; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_452; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_453; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_454; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_455; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_456; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_457; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_458; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_459; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_460; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_461; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_462; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_463; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_464; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_465; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_466; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_467; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_468; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_469; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_470; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_471; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_472; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_473; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_474; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_475; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_476; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_477; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_478; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_479; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_480; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_481; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_482; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_483; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_484; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_485; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_486; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_487; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_488; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_489; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_490; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_491; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_492; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_493; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_494; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_495; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_496; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_497; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_498; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_499; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_500; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_501; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_502; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_503; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_504; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_505; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_506; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_507; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_508; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_509; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_510; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_511; // @[matcher_pisa.scala 333:23]
  wire [3:0] pipe1_io_pipe_phv_out_next_processor_id; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_pipe_phv_out_next_config_id; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_pipe_phv_out_is_valid_processor; // @[matcher_pisa.scala 333:23]
  wire [1:0] pipe1_io_key_config_0_field_config_0; // @[matcher_pisa.scala 333:23]
  wire [1:0] pipe1_io_key_config_0_field_config_1; // @[matcher_pisa.scala 333:23]
  wire [1:0] pipe1_io_key_config_0_field_config_2; // @[matcher_pisa.scala 333:23]
  wire [1:0] pipe1_io_key_config_0_field_config_3; // @[matcher_pisa.scala 333:23]
  wire [1:0] pipe1_io_key_config_0_field_config_4; // @[matcher_pisa.scala 333:23]
  wire [1:0] pipe1_io_key_config_0_field_config_5; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_0_0; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_0_1; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_0_2; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_0_3; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_1_0; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_1_1; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_1_2; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_1_3; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_2_0; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_2_1; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_2_2; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_2_3; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_3_0; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_3_1; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_3_2; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_3_3; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_4_0; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_4_1; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_4_2; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_4_3; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_5_0; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_5_1; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_5_2; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_0_field_mask_5_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_0_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_0_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_0_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_0_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_1_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_1_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_1_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_1_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_2_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_2_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_2_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_2_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_3_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_3_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_3_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_3_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_4_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_4_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_4_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_4_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_5_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_5_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_5_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_0_field_id_5_3; // @[matcher_pisa.scala 333:23]
  wire [1:0] pipe1_io_key_config_1_field_config_0; // @[matcher_pisa.scala 333:23]
  wire [1:0] pipe1_io_key_config_1_field_config_1; // @[matcher_pisa.scala 333:23]
  wire [1:0] pipe1_io_key_config_1_field_config_2; // @[matcher_pisa.scala 333:23]
  wire [1:0] pipe1_io_key_config_1_field_config_3; // @[matcher_pisa.scala 333:23]
  wire [1:0] pipe1_io_key_config_1_field_config_4; // @[matcher_pisa.scala 333:23]
  wire [1:0] pipe1_io_key_config_1_field_config_5; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_0_0; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_0_1; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_0_2; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_0_3; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_1_0; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_1_1; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_1_2; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_1_3; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_2_0; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_2_1; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_2_2; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_2_3; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_3_0; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_3_1; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_3_2; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_3_3; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_4_0; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_4_1; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_4_2; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_4_3; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_5_0; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_5_1; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_5_2; // @[matcher_pisa.scala 333:23]
  wire  pipe1_io_key_config_1_field_mask_5_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_0_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_0_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_0_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_0_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_1_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_1_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_1_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_1_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_2_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_2_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_2_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_2_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_3_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_3_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_3_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_3_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_4_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_4_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_4_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_4_3; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_5_0; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_5_1; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_5_2; // @[matcher_pisa.scala 333:23]
  wire [7:0] pipe1_io_key_config_1_field_id_5_3; // @[matcher_pisa.scala 333:23]
  wire [191:0] pipe1_io_match_key; // @[matcher_pisa.scala 333:23]
  wire  pipe2_clock; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_0; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_1; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_2; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_3; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_4; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_5; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_6; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_7; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_8; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_9; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_10; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_11; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_12; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_13; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_14; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_15; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_16; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_17; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_18; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_19; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_20; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_21; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_22; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_23; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_24; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_25; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_26; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_27; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_28; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_29; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_30; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_31; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_32; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_33; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_34; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_35; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_36; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_37; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_38; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_39; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_40; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_41; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_42; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_43; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_44; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_45; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_46; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_47; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_48; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_49; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_50; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_51; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_52; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_53; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_54; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_55; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_56; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_57; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_58; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_59; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_60; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_61; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_62; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_63; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_64; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_65; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_66; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_67; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_68; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_69; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_70; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_71; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_72; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_73; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_74; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_75; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_76; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_77; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_78; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_79; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_80; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_81; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_82; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_83; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_84; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_85; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_86; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_87; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_88; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_89; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_90; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_91; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_92; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_93; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_94; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_95; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_96; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_97; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_98; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_99; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_100; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_101; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_102; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_103; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_104; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_105; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_106; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_107; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_108; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_109; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_110; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_111; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_112; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_113; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_114; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_115; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_116; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_117; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_118; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_119; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_120; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_121; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_122; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_123; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_124; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_125; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_126; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_127; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_128; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_129; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_130; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_131; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_132; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_133; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_134; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_135; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_136; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_137; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_138; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_139; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_140; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_141; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_142; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_143; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_144; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_145; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_146; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_147; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_148; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_149; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_150; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_151; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_152; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_153; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_154; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_155; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_156; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_157; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_158; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_159; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_160; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_161; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_162; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_163; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_164; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_165; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_166; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_167; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_168; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_169; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_170; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_171; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_172; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_173; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_174; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_175; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_176; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_177; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_178; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_179; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_180; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_181; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_182; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_183; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_184; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_185; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_186; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_187; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_188; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_189; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_190; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_191; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_192; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_193; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_194; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_195; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_196; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_197; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_198; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_199; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_200; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_201; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_202; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_203; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_204; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_205; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_206; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_207; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_208; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_209; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_210; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_211; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_212; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_213; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_214; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_215; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_216; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_217; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_218; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_219; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_220; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_221; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_222; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_223; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_224; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_225; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_226; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_227; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_228; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_229; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_230; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_231; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_232; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_233; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_234; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_235; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_236; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_237; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_238; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_239; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_240; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_241; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_242; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_243; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_244; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_245; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_246; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_247; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_248; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_249; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_250; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_251; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_252; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_253; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_254; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_255; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_256; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_257; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_258; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_259; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_260; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_261; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_262; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_263; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_264; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_265; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_266; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_267; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_268; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_269; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_270; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_271; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_272; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_273; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_274; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_275; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_276; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_277; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_278; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_279; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_280; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_281; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_282; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_283; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_284; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_285; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_286; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_287; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_288; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_289; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_290; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_291; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_292; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_293; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_294; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_295; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_296; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_297; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_298; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_299; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_300; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_301; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_302; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_303; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_304; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_305; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_306; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_307; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_308; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_309; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_310; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_311; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_312; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_313; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_314; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_315; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_316; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_317; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_318; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_319; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_320; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_321; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_322; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_323; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_324; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_325; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_326; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_327; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_328; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_329; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_330; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_331; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_332; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_333; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_334; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_335; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_336; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_337; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_338; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_339; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_340; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_341; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_342; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_343; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_344; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_345; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_346; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_347; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_348; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_349; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_350; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_351; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_352; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_353; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_354; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_355; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_356; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_357; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_358; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_359; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_360; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_361; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_362; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_363; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_364; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_365; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_366; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_367; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_368; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_369; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_370; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_371; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_372; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_373; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_374; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_375; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_376; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_377; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_378; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_379; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_380; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_381; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_382; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_383; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_384; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_385; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_386; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_387; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_388; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_389; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_390; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_391; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_392; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_393; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_394; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_395; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_396; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_397; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_398; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_399; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_400; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_401; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_402; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_403; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_404; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_405; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_406; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_407; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_408; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_409; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_410; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_411; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_412; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_413; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_414; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_415; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_416; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_417; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_418; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_419; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_420; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_421; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_422; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_423; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_424; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_425; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_426; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_427; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_428; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_429; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_430; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_431; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_432; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_433; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_434; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_435; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_436; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_437; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_438; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_439; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_440; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_441; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_442; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_443; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_444; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_445; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_446; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_447; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_448; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_449; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_450; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_451; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_452; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_453; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_454; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_455; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_456; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_457; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_458; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_459; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_460; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_461; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_462; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_463; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_464; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_465; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_466; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_467; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_468; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_469; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_470; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_471; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_472; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_473; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_474; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_475; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_476; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_477; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_478; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_479; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_480; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_481; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_482; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_483; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_484; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_485; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_486; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_487; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_488; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_489; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_490; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_491; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_492; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_493; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_494; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_495; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_496; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_497; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_498; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_499; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_500; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_501; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_502; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_503; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_504; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_505; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_506; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_507; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_508; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_509; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_510; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_511; // @[matcher_pisa.scala 334:23]
  wire [3:0] pipe2_io_pipe_phv_in_next_processor_id; // @[matcher_pisa.scala 334:23]
  wire  pipe2_io_pipe_phv_in_next_config_id; // @[matcher_pisa.scala 334:23]
  wire  pipe2_io_pipe_phv_in_is_valid_processor; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_0; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_1; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_2; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_3; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_4; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_5; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_6; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_7; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_8; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_9; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_10; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_11; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_12; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_13; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_14; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_15; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_16; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_17; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_18; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_19; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_20; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_21; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_22; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_23; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_24; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_25; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_26; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_27; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_28; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_29; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_30; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_31; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_32; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_33; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_34; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_35; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_36; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_37; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_38; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_39; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_40; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_41; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_42; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_43; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_44; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_45; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_46; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_47; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_48; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_49; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_50; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_51; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_52; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_53; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_54; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_55; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_56; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_57; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_58; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_59; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_60; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_61; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_62; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_63; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_64; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_65; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_66; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_67; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_68; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_69; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_70; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_71; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_72; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_73; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_74; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_75; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_76; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_77; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_78; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_79; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_80; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_81; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_82; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_83; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_84; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_85; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_86; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_87; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_88; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_89; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_90; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_91; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_92; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_93; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_94; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_95; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_96; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_97; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_98; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_99; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_100; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_101; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_102; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_103; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_104; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_105; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_106; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_107; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_108; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_109; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_110; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_111; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_112; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_113; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_114; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_115; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_116; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_117; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_118; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_119; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_120; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_121; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_122; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_123; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_124; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_125; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_126; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_127; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_128; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_129; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_130; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_131; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_132; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_133; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_134; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_135; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_136; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_137; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_138; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_139; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_140; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_141; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_142; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_143; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_144; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_145; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_146; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_147; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_148; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_149; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_150; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_151; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_152; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_153; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_154; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_155; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_156; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_157; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_158; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_159; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_160; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_161; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_162; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_163; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_164; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_165; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_166; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_167; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_168; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_169; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_170; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_171; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_172; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_173; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_174; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_175; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_176; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_177; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_178; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_179; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_180; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_181; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_182; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_183; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_184; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_185; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_186; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_187; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_188; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_189; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_190; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_191; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_192; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_193; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_194; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_195; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_196; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_197; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_198; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_199; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_200; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_201; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_202; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_203; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_204; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_205; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_206; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_207; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_208; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_209; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_210; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_211; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_212; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_213; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_214; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_215; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_216; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_217; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_218; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_219; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_220; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_221; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_222; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_223; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_224; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_225; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_226; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_227; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_228; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_229; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_230; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_231; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_232; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_233; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_234; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_235; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_236; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_237; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_238; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_239; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_240; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_241; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_242; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_243; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_244; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_245; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_246; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_247; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_248; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_249; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_250; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_251; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_252; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_253; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_254; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_255; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_256; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_257; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_258; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_259; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_260; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_261; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_262; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_263; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_264; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_265; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_266; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_267; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_268; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_269; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_270; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_271; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_272; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_273; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_274; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_275; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_276; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_277; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_278; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_279; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_280; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_281; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_282; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_283; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_284; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_285; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_286; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_287; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_288; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_289; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_290; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_291; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_292; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_293; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_294; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_295; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_296; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_297; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_298; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_299; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_300; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_301; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_302; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_303; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_304; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_305; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_306; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_307; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_308; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_309; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_310; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_311; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_312; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_313; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_314; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_315; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_316; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_317; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_318; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_319; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_320; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_321; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_322; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_323; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_324; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_325; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_326; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_327; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_328; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_329; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_330; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_331; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_332; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_333; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_334; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_335; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_336; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_337; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_338; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_339; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_340; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_341; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_342; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_343; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_344; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_345; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_346; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_347; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_348; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_349; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_350; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_351; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_352; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_353; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_354; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_355; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_356; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_357; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_358; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_359; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_360; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_361; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_362; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_363; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_364; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_365; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_366; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_367; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_368; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_369; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_370; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_371; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_372; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_373; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_374; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_375; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_376; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_377; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_378; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_379; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_380; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_381; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_382; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_383; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_384; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_385; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_386; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_387; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_388; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_389; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_390; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_391; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_392; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_393; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_394; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_395; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_396; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_397; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_398; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_399; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_400; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_401; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_402; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_403; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_404; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_405; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_406; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_407; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_408; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_409; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_410; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_411; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_412; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_413; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_414; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_415; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_416; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_417; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_418; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_419; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_420; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_421; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_422; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_423; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_424; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_425; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_426; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_427; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_428; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_429; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_430; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_431; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_432; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_433; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_434; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_435; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_436; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_437; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_438; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_439; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_440; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_441; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_442; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_443; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_444; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_445; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_446; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_447; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_448; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_449; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_450; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_451; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_452; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_453; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_454; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_455; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_456; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_457; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_458; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_459; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_460; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_461; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_462; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_463; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_464; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_465; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_466; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_467; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_468; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_469; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_470; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_471; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_472; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_473; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_474; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_475; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_476; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_477; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_478; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_479; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_480; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_481; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_482; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_483; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_484; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_485; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_486; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_487; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_488; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_489; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_490; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_491; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_492; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_493; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_494; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_495; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_496; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_497; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_498; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_499; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_500; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_501; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_502; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_503; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_504; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_505; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_506; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_507; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_508; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_509; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_510; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_511; // @[matcher_pisa.scala 334:23]
  wire [3:0] pipe2_io_pipe_phv_out_next_processor_id; // @[matcher_pisa.scala 334:23]
  wire  pipe2_io_pipe_phv_out_next_config_id; // @[matcher_pisa.scala 334:23]
  wire  pipe2_io_pipe_phv_out_is_valid_processor; // @[matcher_pisa.scala 334:23]
  wire  pipe2_io_mod_hash_depth_mod; // @[matcher_pisa.scala 334:23]
  wire  pipe2_io_mod_config_id; // @[matcher_pisa.scala 334:23]
  wire [3:0] pipe2_io_mod_hash_depth; // @[matcher_pisa.scala 334:23]
  wire [191:0] pipe2_io_key_in; // @[matcher_pisa.scala 334:23]
  wire [191:0] pipe2_io_key_out; // @[matcher_pisa.scala 334:23]
  wire [7:0] pipe2_io_hash_val; // @[matcher_pisa.scala 334:23]
  wire [3:0] pipe2_io_hash_val_cs; // @[matcher_pisa.scala 334:23]
  wire  pipe3_clock; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_0; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_1; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_2; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_3; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_4; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_5; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_6; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_7; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_8; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_9; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_10; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_11; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_12; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_13; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_14; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_15; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_16; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_17; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_18; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_19; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_20; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_21; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_22; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_23; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_24; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_25; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_26; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_27; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_28; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_29; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_30; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_31; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_32; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_33; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_34; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_35; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_36; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_37; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_38; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_39; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_40; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_41; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_42; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_43; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_44; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_45; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_46; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_47; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_48; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_49; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_50; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_51; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_52; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_53; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_54; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_55; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_56; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_57; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_58; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_59; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_60; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_61; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_62; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_63; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_64; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_65; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_66; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_67; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_68; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_69; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_70; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_71; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_72; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_73; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_74; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_75; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_76; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_77; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_78; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_79; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_80; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_81; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_82; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_83; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_84; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_85; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_86; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_87; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_88; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_89; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_90; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_91; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_92; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_93; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_94; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_95; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_96; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_97; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_98; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_99; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_100; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_101; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_102; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_103; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_104; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_105; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_106; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_107; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_108; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_109; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_110; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_111; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_112; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_113; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_114; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_115; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_116; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_117; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_118; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_119; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_120; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_121; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_122; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_123; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_124; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_125; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_126; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_127; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_128; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_129; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_130; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_131; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_132; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_133; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_134; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_135; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_136; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_137; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_138; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_139; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_140; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_141; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_142; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_143; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_144; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_145; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_146; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_147; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_148; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_149; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_150; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_151; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_152; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_153; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_154; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_155; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_156; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_157; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_158; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_159; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_160; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_161; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_162; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_163; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_164; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_165; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_166; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_167; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_168; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_169; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_170; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_171; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_172; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_173; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_174; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_175; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_176; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_177; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_178; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_179; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_180; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_181; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_182; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_183; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_184; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_185; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_186; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_187; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_188; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_189; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_190; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_191; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_192; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_193; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_194; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_195; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_196; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_197; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_198; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_199; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_200; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_201; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_202; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_203; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_204; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_205; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_206; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_207; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_208; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_209; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_210; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_211; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_212; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_213; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_214; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_215; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_216; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_217; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_218; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_219; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_220; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_221; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_222; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_223; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_224; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_225; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_226; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_227; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_228; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_229; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_230; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_231; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_232; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_233; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_234; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_235; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_236; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_237; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_238; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_239; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_240; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_241; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_242; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_243; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_244; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_245; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_246; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_247; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_248; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_249; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_250; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_251; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_252; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_253; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_254; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_255; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_256; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_257; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_258; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_259; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_260; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_261; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_262; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_263; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_264; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_265; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_266; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_267; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_268; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_269; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_270; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_271; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_272; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_273; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_274; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_275; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_276; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_277; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_278; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_279; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_280; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_281; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_282; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_283; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_284; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_285; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_286; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_287; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_288; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_289; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_290; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_291; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_292; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_293; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_294; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_295; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_296; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_297; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_298; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_299; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_300; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_301; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_302; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_303; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_304; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_305; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_306; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_307; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_308; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_309; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_310; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_311; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_312; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_313; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_314; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_315; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_316; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_317; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_318; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_319; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_320; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_321; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_322; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_323; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_324; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_325; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_326; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_327; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_328; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_329; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_330; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_331; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_332; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_333; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_334; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_335; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_336; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_337; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_338; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_339; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_340; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_341; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_342; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_343; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_344; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_345; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_346; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_347; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_348; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_349; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_350; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_351; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_352; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_353; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_354; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_355; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_356; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_357; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_358; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_359; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_360; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_361; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_362; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_363; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_364; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_365; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_366; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_367; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_368; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_369; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_370; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_371; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_372; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_373; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_374; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_375; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_376; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_377; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_378; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_379; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_380; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_381; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_382; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_383; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_384; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_385; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_386; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_387; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_388; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_389; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_390; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_391; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_392; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_393; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_394; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_395; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_396; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_397; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_398; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_399; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_400; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_401; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_402; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_403; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_404; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_405; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_406; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_407; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_408; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_409; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_410; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_411; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_412; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_413; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_414; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_415; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_416; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_417; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_418; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_419; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_420; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_421; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_422; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_423; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_424; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_425; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_426; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_427; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_428; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_429; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_430; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_431; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_432; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_433; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_434; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_435; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_436; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_437; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_438; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_439; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_440; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_441; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_442; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_443; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_444; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_445; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_446; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_447; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_448; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_449; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_450; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_451; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_452; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_453; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_454; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_455; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_456; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_457; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_458; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_459; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_460; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_461; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_462; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_463; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_464; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_465; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_466; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_467; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_468; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_469; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_470; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_471; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_472; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_473; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_474; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_475; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_476; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_477; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_478; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_479; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_480; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_481; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_482; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_483; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_484; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_485; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_486; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_487; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_488; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_489; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_490; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_491; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_492; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_493; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_494; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_495; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_496; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_497; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_498; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_499; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_500; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_501; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_502; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_503; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_504; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_505; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_506; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_507; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_508; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_509; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_510; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_511; // @[matcher_pisa.scala 335:23]
  wire [3:0] pipe3_io_pipe_phv_in_next_processor_id; // @[matcher_pisa.scala 335:23]
  wire  pipe3_io_pipe_phv_in_next_config_id; // @[matcher_pisa.scala 335:23]
  wire  pipe3_io_pipe_phv_in_is_valid_processor; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_0; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_1; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_2; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_3; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_4; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_5; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_6; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_7; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_8; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_9; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_10; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_11; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_12; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_13; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_14; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_15; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_16; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_17; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_18; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_19; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_20; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_21; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_22; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_23; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_24; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_25; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_26; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_27; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_28; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_29; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_30; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_31; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_32; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_33; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_34; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_35; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_36; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_37; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_38; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_39; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_40; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_41; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_42; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_43; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_44; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_45; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_46; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_47; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_48; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_49; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_50; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_51; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_52; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_53; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_54; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_55; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_56; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_57; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_58; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_59; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_60; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_61; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_62; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_63; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_64; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_65; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_66; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_67; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_68; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_69; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_70; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_71; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_72; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_73; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_74; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_75; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_76; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_77; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_78; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_79; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_80; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_81; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_82; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_83; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_84; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_85; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_86; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_87; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_88; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_89; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_90; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_91; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_92; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_93; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_94; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_95; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_96; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_97; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_98; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_99; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_100; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_101; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_102; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_103; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_104; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_105; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_106; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_107; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_108; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_109; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_110; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_111; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_112; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_113; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_114; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_115; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_116; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_117; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_118; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_119; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_120; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_121; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_122; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_123; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_124; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_125; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_126; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_127; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_128; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_129; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_130; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_131; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_132; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_133; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_134; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_135; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_136; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_137; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_138; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_139; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_140; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_141; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_142; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_143; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_144; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_145; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_146; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_147; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_148; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_149; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_150; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_151; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_152; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_153; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_154; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_155; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_156; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_157; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_158; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_159; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_160; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_161; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_162; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_163; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_164; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_165; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_166; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_167; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_168; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_169; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_170; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_171; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_172; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_173; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_174; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_175; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_176; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_177; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_178; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_179; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_180; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_181; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_182; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_183; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_184; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_185; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_186; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_187; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_188; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_189; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_190; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_191; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_192; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_193; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_194; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_195; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_196; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_197; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_198; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_199; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_200; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_201; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_202; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_203; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_204; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_205; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_206; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_207; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_208; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_209; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_210; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_211; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_212; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_213; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_214; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_215; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_216; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_217; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_218; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_219; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_220; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_221; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_222; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_223; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_224; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_225; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_226; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_227; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_228; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_229; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_230; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_231; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_232; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_233; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_234; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_235; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_236; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_237; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_238; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_239; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_240; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_241; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_242; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_243; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_244; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_245; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_246; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_247; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_248; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_249; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_250; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_251; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_252; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_253; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_254; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_255; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_256; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_257; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_258; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_259; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_260; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_261; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_262; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_263; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_264; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_265; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_266; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_267; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_268; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_269; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_270; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_271; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_272; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_273; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_274; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_275; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_276; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_277; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_278; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_279; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_280; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_281; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_282; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_283; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_284; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_285; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_286; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_287; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_288; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_289; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_290; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_291; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_292; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_293; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_294; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_295; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_296; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_297; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_298; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_299; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_300; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_301; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_302; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_303; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_304; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_305; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_306; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_307; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_308; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_309; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_310; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_311; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_312; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_313; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_314; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_315; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_316; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_317; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_318; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_319; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_320; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_321; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_322; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_323; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_324; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_325; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_326; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_327; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_328; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_329; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_330; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_331; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_332; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_333; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_334; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_335; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_336; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_337; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_338; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_339; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_340; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_341; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_342; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_343; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_344; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_345; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_346; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_347; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_348; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_349; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_350; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_351; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_352; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_353; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_354; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_355; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_356; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_357; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_358; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_359; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_360; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_361; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_362; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_363; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_364; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_365; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_366; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_367; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_368; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_369; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_370; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_371; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_372; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_373; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_374; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_375; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_376; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_377; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_378; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_379; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_380; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_381; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_382; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_383; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_384; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_385; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_386; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_387; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_388; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_389; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_390; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_391; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_392; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_393; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_394; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_395; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_396; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_397; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_398; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_399; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_400; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_401; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_402; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_403; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_404; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_405; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_406; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_407; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_408; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_409; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_410; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_411; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_412; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_413; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_414; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_415; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_416; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_417; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_418; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_419; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_420; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_421; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_422; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_423; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_424; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_425; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_426; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_427; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_428; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_429; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_430; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_431; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_432; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_433; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_434; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_435; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_436; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_437; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_438; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_439; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_440; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_441; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_442; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_443; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_444; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_445; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_446; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_447; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_448; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_449; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_450; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_451; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_452; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_453; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_454; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_455; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_456; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_457; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_458; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_459; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_460; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_461; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_462; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_463; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_464; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_465; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_466; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_467; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_468; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_469; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_470; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_471; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_472; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_473; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_474; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_475; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_476; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_477; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_478; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_479; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_480; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_481; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_482; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_483; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_484; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_485; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_486; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_487; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_488; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_489; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_490; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_491; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_492; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_493; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_494; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_495; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_496; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_497; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_498; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_499; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_500; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_501; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_502; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_503; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_504; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_505; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_506; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_507; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_508; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_509; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_510; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_511; // @[matcher_pisa.scala 335:23]
  wire [3:0] pipe3_io_pipe_phv_out_next_processor_id; // @[matcher_pisa.scala 335:23]
  wire  pipe3_io_pipe_phv_out_next_config_id; // @[matcher_pisa.scala 335:23]
  wire  pipe3_io_pipe_phv_out_is_valid_processor; // @[matcher_pisa.scala 335:23]
  wire [4:0] pipe3_io_table_config_0_table_depth; // @[matcher_pisa.scala 335:23]
  wire [4:0] pipe3_io_table_config_0_table_width; // @[matcher_pisa.scala 335:23]
  wire [4:0] pipe3_io_table_config_1_table_depth; // @[matcher_pisa.scala 335:23]
  wire [4:0] pipe3_io_table_config_1_table_width; // @[matcher_pisa.scala 335:23]
  wire [191:0] pipe3_io_key_in; // @[matcher_pisa.scala 335:23]
  wire [191:0] pipe3_io_key_out; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_addr_in; // @[matcher_pisa.scala 335:23]
  wire [3:0] pipe3_io_cs_in; // @[matcher_pisa.scala 335:23]
  wire [255:0] pipe3_io_data_out; // @[matcher_pisa.scala 335:23]
  wire  pipe3_io_w_en; // @[matcher_pisa.scala 335:23]
  wire [3:0] pipe3_io_w_sram_id; // @[matcher_pisa.scala 335:23]
  wire [7:0] pipe3_io_w_addr; // @[matcher_pisa.scala 335:23]
  wire [63:0] pipe3_io_w_data; // @[matcher_pisa.scala 335:23]
  wire  pipe4_clock; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_0; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_1; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_2; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_3; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_4; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_5; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_6; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_7; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_8; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_9; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_10; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_11; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_12; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_13; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_14; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_15; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_16; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_17; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_18; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_19; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_20; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_21; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_22; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_23; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_24; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_25; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_26; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_27; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_28; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_29; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_30; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_31; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_32; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_33; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_34; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_35; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_36; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_37; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_38; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_39; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_40; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_41; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_42; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_43; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_44; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_45; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_46; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_47; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_48; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_49; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_50; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_51; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_52; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_53; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_54; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_55; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_56; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_57; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_58; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_59; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_60; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_61; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_62; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_63; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_64; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_65; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_66; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_67; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_68; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_69; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_70; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_71; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_72; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_73; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_74; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_75; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_76; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_77; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_78; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_79; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_80; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_81; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_82; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_83; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_84; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_85; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_86; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_87; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_88; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_89; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_90; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_91; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_92; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_93; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_94; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_95; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_96; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_97; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_98; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_99; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_100; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_101; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_102; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_103; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_104; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_105; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_106; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_107; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_108; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_109; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_110; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_111; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_112; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_113; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_114; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_115; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_116; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_117; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_118; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_119; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_120; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_121; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_122; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_123; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_124; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_125; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_126; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_127; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_128; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_129; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_130; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_131; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_132; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_133; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_134; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_135; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_136; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_137; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_138; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_139; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_140; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_141; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_142; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_143; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_144; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_145; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_146; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_147; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_148; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_149; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_150; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_151; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_152; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_153; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_154; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_155; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_156; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_157; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_158; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_159; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_160; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_161; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_162; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_163; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_164; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_165; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_166; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_167; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_168; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_169; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_170; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_171; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_172; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_173; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_174; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_175; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_176; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_177; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_178; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_179; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_180; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_181; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_182; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_183; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_184; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_185; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_186; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_187; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_188; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_189; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_190; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_191; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_192; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_193; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_194; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_195; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_196; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_197; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_198; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_199; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_200; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_201; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_202; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_203; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_204; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_205; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_206; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_207; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_208; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_209; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_210; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_211; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_212; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_213; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_214; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_215; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_216; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_217; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_218; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_219; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_220; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_221; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_222; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_223; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_224; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_225; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_226; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_227; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_228; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_229; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_230; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_231; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_232; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_233; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_234; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_235; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_236; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_237; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_238; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_239; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_240; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_241; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_242; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_243; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_244; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_245; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_246; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_247; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_248; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_249; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_250; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_251; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_252; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_253; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_254; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_255; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_256; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_257; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_258; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_259; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_260; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_261; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_262; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_263; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_264; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_265; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_266; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_267; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_268; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_269; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_270; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_271; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_272; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_273; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_274; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_275; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_276; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_277; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_278; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_279; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_280; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_281; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_282; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_283; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_284; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_285; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_286; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_287; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_288; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_289; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_290; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_291; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_292; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_293; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_294; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_295; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_296; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_297; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_298; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_299; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_300; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_301; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_302; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_303; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_304; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_305; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_306; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_307; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_308; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_309; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_310; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_311; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_312; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_313; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_314; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_315; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_316; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_317; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_318; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_319; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_320; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_321; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_322; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_323; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_324; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_325; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_326; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_327; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_328; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_329; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_330; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_331; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_332; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_333; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_334; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_335; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_336; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_337; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_338; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_339; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_340; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_341; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_342; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_343; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_344; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_345; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_346; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_347; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_348; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_349; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_350; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_351; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_352; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_353; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_354; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_355; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_356; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_357; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_358; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_359; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_360; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_361; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_362; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_363; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_364; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_365; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_366; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_367; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_368; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_369; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_370; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_371; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_372; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_373; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_374; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_375; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_376; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_377; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_378; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_379; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_380; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_381; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_382; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_383; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_384; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_385; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_386; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_387; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_388; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_389; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_390; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_391; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_392; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_393; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_394; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_395; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_396; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_397; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_398; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_399; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_400; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_401; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_402; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_403; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_404; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_405; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_406; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_407; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_408; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_409; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_410; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_411; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_412; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_413; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_414; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_415; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_416; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_417; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_418; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_419; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_420; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_421; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_422; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_423; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_424; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_425; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_426; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_427; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_428; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_429; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_430; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_431; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_432; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_433; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_434; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_435; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_436; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_437; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_438; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_439; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_440; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_441; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_442; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_443; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_444; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_445; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_446; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_447; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_448; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_449; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_450; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_451; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_452; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_453; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_454; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_455; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_456; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_457; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_458; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_459; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_460; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_461; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_462; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_463; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_464; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_465; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_466; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_467; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_468; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_469; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_470; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_471; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_472; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_473; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_474; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_475; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_476; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_477; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_478; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_479; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_480; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_481; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_482; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_483; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_484; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_485; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_486; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_487; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_488; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_489; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_490; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_491; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_492; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_493; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_494; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_495; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_496; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_497; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_498; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_499; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_500; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_501; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_502; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_503; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_504; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_505; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_506; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_507; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_508; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_509; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_510; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_511; // @[matcher_pisa.scala 336:23]
  wire [3:0] pipe4_io_pipe_phv_in_next_processor_id; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_pipe_phv_in_next_config_id; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_pipe_phv_in_is_valid_processor; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_0; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_1; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_2; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_3; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_4; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_5; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_6; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_7; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_8; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_9; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_10; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_11; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_12; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_13; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_14; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_15; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_16; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_17; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_18; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_19; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_20; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_21; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_22; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_23; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_24; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_25; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_26; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_27; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_28; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_29; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_30; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_31; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_32; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_33; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_34; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_35; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_36; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_37; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_38; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_39; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_40; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_41; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_42; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_43; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_44; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_45; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_46; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_47; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_48; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_49; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_50; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_51; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_52; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_53; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_54; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_55; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_56; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_57; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_58; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_59; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_60; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_61; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_62; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_63; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_64; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_65; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_66; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_67; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_68; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_69; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_70; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_71; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_72; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_73; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_74; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_75; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_76; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_77; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_78; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_79; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_80; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_81; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_82; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_83; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_84; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_85; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_86; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_87; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_88; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_89; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_90; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_91; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_92; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_93; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_94; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_95; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_96; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_97; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_98; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_99; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_100; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_101; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_102; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_103; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_104; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_105; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_106; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_107; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_108; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_109; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_110; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_111; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_112; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_113; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_114; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_115; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_116; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_117; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_118; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_119; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_120; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_121; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_122; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_123; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_124; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_125; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_126; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_127; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_128; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_129; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_130; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_131; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_132; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_133; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_134; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_135; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_136; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_137; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_138; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_139; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_140; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_141; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_142; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_143; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_144; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_145; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_146; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_147; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_148; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_149; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_150; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_151; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_152; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_153; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_154; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_155; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_156; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_157; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_158; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_159; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_160; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_161; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_162; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_163; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_164; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_165; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_166; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_167; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_168; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_169; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_170; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_171; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_172; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_173; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_174; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_175; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_176; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_177; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_178; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_179; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_180; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_181; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_182; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_183; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_184; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_185; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_186; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_187; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_188; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_189; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_190; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_191; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_192; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_193; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_194; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_195; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_196; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_197; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_198; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_199; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_200; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_201; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_202; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_203; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_204; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_205; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_206; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_207; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_208; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_209; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_210; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_211; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_212; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_213; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_214; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_215; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_216; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_217; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_218; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_219; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_220; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_221; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_222; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_223; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_224; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_225; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_226; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_227; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_228; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_229; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_230; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_231; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_232; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_233; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_234; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_235; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_236; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_237; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_238; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_239; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_240; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_241; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_242; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_243; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_244; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_245; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_246; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_247; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_248; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_249; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_250; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_251; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_252; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_253; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_254; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_255; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_256; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_257; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_258; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_259; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_260; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_261; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_262; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_263; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_264; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_265; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_266; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_267; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_268; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_269; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_270; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_271; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_272; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_273; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_274; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_275; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_276; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_277; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_278; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_279; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_280; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_281; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_282; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_283; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_284; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_285; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_286; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_287; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_288; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_289; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_290; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_291; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_292; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_293; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_294; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_295; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_296; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_297; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_298; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_299; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_300; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_301; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_302; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_303; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_304; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_305; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_306; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_307; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_308; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_309; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_310; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_311; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_312; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_313; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_314; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_315; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_316; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_317; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_318; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_319; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_320; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_321; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_322; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_323; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_324; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_325; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_326; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_327; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_328; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_329; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_330; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_331; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_332; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_333; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_334; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_335; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_336; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_337; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_338; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_339; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_340; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_341; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_342; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_343; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_344; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_345; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_346; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_347; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_348; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_349; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_350; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_351; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_352; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_353; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_354; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_355; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_356; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_357; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_358; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_359; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_360; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_361; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_362; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_363; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_364; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_365; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_366; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_367; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_368; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_369; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_370; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_371; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_372; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_373; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_374; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_375; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_376; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_377; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_378; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_379; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_380; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_381; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_382; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_383; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_384; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_385; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_386; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_387; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_388; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_389; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_390; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_391; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_392; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_393; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_394; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_395; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_396; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_397; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_398; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_399; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_400; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_401; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_402; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_403; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_404; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_405; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_406; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_407; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_408; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_409; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_410; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_411; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_412; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_413; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_414; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_415; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_416; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_417; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_418; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_419; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_420; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_421; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_422; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_423; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_424; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_425; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_426; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_427; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_428; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_429; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_430; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_431; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_432; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_433; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_434; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_435; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_436; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_437; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_438; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_439; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_440; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_441; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_442; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_443; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_444; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_445; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_446; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_447; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_448; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_449; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_450; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_451; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_452; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_453; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_454; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_455; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_456; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_457; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_458; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_459; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_460; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_461; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_462; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_463; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_464; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_465; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_466; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_467; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_468; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_469; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_470; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_471; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_472; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_473; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_474; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_475; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_476; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_477; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_478; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_479; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_480; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_481; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_482; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_483; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_484; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_485; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_486; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_487; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_488; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_489; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_490; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_491; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_492; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_493; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_494; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_495; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_496; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_497; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_498; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_499; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_500; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_501; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_502; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_503; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_504; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_505; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_506; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_507; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_508; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_509; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_510; // @[matcher_pisa.scala 336:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_511; // @[matcher_pisa.scala 336:23]
  wire [3:0] pipe4_io_pipe_phv_out_next_processor_id; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_pipe_phv_out_next_config_id; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_pipe_phv_out_is_valid_processor; // @[matcher_pisa.scala 336:23]
  wire [1:0] pipe4_io_key_config_0_field_config_0; // @[matcher_pisa.scala 336:23]
  wire [1:0] pipe4_io_key_config_0_field_config_1; // @[matcher_pisa.scala 336:23]
  wire [1:0] pipe4_io_key_config_0_field_config_2; // @[matcher_pisa.scala 336:23]
  wire [1:0] pipe4_io_key_config_0_field_config_3; // @[matcher_pisa.scala 336:23]
  wire [1:0] pipe4_io_key_config_0_field_config_4; // @[matcher_pisa.scala 336:23]
  wire [1:0] pipe4_io_key_config_0_field_config_5; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_0_0; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_0_1; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_0_2; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_0_3; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_1_0; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_1_1; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_1_2; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_1_3; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_2_0; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_2_1; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_2_2; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_2_3; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_3_0; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_3_1; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_3_2; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_3_3; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_4_0; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_4_1; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_4_2; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_4_3; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_5_0; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_5_1; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_5_2; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_0_field_mask_5_3; // @[matcher_pisa.scala 336:23]
  wire [1:0] pipe4_io_key_config_1_field_config_0; // @[matcher_pisa.scala 336:23]
  wire [1:0] pipe4_io_key_config_1_field_config_1; // @[matcher_pisa.scala 336:23]
  wire [1:0] pipe4_io_key_config_1_field_config_2; // @[matcher_pisa.scala 336:23]
  wire [1:0] pipe4_io_key_config_1_field_config_3; // @[matcher_pisa.scala 336:23]
  wire [1:0] pipe4_io_key_config_1_field_config_4; // @[matcher_pisa.scala 336:23]
  wire [1:0] pipe4_io_key_config_1_field_config_5; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_0_0; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_0_1; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_0_2; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_0_3; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_1_0; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_1_1; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_1_2; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_1_3; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_2_0; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_2_1; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_2_2; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_2_3; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_3_0; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_3_1; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_3_2; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_3_3; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_4_0; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_4_1; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_4_2; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_4_3; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_5_0; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_5_1; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_5_2; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_key_config_1_field_mask_5_3; // @[matcher_pisa.scala 336:23]
  wire [191:0] pipe4_io_key_in; // @[matcher_pisa.scala 336:23]
  wire [255:0] pipe4_io_data_in; // @[matcher_pisa.scala 336:23]
  wire  pipe4_io_hit; // @[matcher_pisa.scala 336:23]
  wire [63:0] pipe4_io_match_value; // @[matcher_pisa.scala 336:23]
  reg [1:0] key_config_0_field_config_0; // @[matcher_pisa.scala 70:25]
  reg [1:0] key_config_0_field_config_1; // @[matcher_pisa.scala 70:25]
  reg [1:0] key_config_0_field_config_2; // @[matcher_pisa.scala 70:25]
  reg [1:0] key_config_0_field_config_3; // @[matcher_pisa.scala 70:25]
  reg [1:0] key_config_0_field_config_4; // @[matcher_pisa.scala 70:25]
  reg [1:0] key_config_0_field_config_5; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_0_0; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_0_1; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_0_2; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_0_3; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_1_0; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_1_1; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_1_2; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_1_3; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_2_0; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_2_1; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_2_2; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_2_3; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_3_0; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_3_1; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_3_2; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_3_3; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_4_0; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_4_1; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_4_2; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_4_3; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_5_0; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_5_1; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_5_2; // @[matcher_pisa.scala 70:25]
  reg  key_config_0_field_mask_5_3; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_0_0; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_0_1; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_0_2; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_0_3; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_1_0; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_1_1; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_1_2; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_1_3; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_2_0; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_2_1; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_2_2; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_2_3; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_3_0; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_3_1; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_3_2; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_3_3; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_4_0; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_4_1; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_4_2; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_4_3; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_5_0; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_5_1; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_5_2; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_0_field_id_5_3; // @[matcher_pisa.scala 70:25]
  reg [1:0] key_config_1_field_config_0; // @[matcher_pisa.scala 70:25]
  reg [1:0] key_config_1_field_config_1; // @[matcher_pisa.scala 70:25]
  reg [1:0] key_config_1_field_config_2; // @[matcher_pisa.scala 70:25]
  reg [1:0] key_config_1_field_config_3; // @[matcher_pisa.scala 70:25]
  reg [1:0] key_config_1_field_config_4; // @[matcher_pisa.scala 70:25]
  reg [1:0] key_config_1_field_config_5; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_0_0; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_0_1; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_0_2; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_0_3; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_1_0; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_1_1; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_1_2; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_1_3; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_2_0; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_2_1; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_2_2; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_2_3; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_3_0; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_3_1; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_3_2; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_3_3; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_4_0; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_4_1; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_4_2; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_4_3; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_5_0; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_5_1; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_5_2; // @[matcher_pisa.scala 70:25]
  reg  key_config_1_field_mask_5_3; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_0_0; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_0_1; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_0_2; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_0_3; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_1_0; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_1_1; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_1_2; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_1_3; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_2_0; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_2_1; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_2_2; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_2_3; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_3_0; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_3_1; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_3_2; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_3_3; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_4_0; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_4_1; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_4_2; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_4_3; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_5_0; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_5_1; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_5_2; // @[matcher_pisa.scala 70:25]
  reg [7:0] key_config_1_field_id_5_3; // @[matcher_pisa.scala 70:25]
  reg [4:0] table_config_0_table_depth; // @[matcher_pisa.scala 71:27]
  reg [4:0] table_config_0_table_width; // @[matcher_pisa.scala 71:27]
  reg [4:0] table_config_1_table_depth; // @[matcher_pisa.scala 71:27]
  reg [4:0] table_config_1_table_width; // @[matcher_pisa.scala 71:27]
  wire  _GEN_338 = ~io_mod_config_id; // @[matcher_pisa.scala 74:83 matcher_pisa.scala 74:83 matcher_pisa.scala 70:25]
  wire  _GEN_339 = 3'h0 == io_mod_key_mod_group_index; // @[matcher_pisa.scala 74:83 matcher_pisa.scala 74:83 matcher_pisa.scala 70:25]
  wire  _GEN_341 = 3'h1 == io_mod_key_mod_group_index; // @[matcher_pisa.scala 74:83 matcher_pisa.scala 74:83 matcher_pisa.scala 70:25]
  wire  _GEN_343 = 3'h2 == io_mod_key_mod_group_index; // @[matcher_pisa.scala 74:83 matcher_pisa.scala 74:83 matcher_pisa.scala 70:25]
  wire  _GEN_345 = 3'h3 == io_mod_key_mod_group_index; // @[matcher_pisa.scala 74:83 matcher_pisa.scala 74:83 matcher_pisa.scala 70:25]
  wire  _GEN_347 = 3'h4 == io_mod_key_mod_group_index; // @[matcher_pisa.scala 74:83 matcher_pisa.scala 74:83 matcher_pisa.scala 70:25]
  wire  _GEN_349 = 3'h5 == io_mod_key_mod_group_index; // @[matcher_pisa.scala 74:83 matcher_pisa.scala 74:83 matcher_pisa.scala 70:25]
  MatchGetKeyPISA pipe1 ( // @[matcher_pisa.scala 333:23]
    .clock(pipe1_clock),
    .io_pipe_phv_in_data_0(pipe1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe1_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe1_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe1_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe1_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe1_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe1_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe1_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe1_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe1_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe1_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe1_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe1_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe1_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe1_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe1_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe1_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe1_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe1_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe1_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe1_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe1_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe1_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe1_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe1_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe1_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe1_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe1_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe1_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe1_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe1_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe1_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe1_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe1_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe1_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe1_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe1_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe1_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe1_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe1_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe1_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe1_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe1_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe1_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe1_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe1_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe1_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe1_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe1_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe1_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe1_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe1_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe1_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe1_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe1_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe1_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe1_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe1_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe1_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe1_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe1_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe1_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe1_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe1_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe1_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe1_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe1_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe1_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe1_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe1_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe1_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe1_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe1_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe1_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe1_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe1_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe1_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe1_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe1_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe1_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe1_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe1_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe1_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe1_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe1_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe1_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe1_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe1_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe1_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe1_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe1_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe1_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe1_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe1_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe1_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe1_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe1_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe1_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe1_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe1_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe1_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe1_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe1_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe1_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe1_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe1_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe1_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe1_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe1_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe1_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe1_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe1_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe1_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe1_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe1_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe1_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe1_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe1_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe1_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe1_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe1_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe1_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe1_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe1_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe1_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe1_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe1_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe1_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe1_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe1_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe1_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe1_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe1_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe1_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe1_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe1_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe1_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe1_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe1_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe1_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe1_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe1_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe1_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe1_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe1_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe1_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe1_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe1_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe1_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe1_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe1_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe1_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe1_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe1_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe1_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe1_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe1_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe1_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe1_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe1_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe1_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(pipe1_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(pipe1_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(pipe1_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(pipe1_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(pipe1_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(pipe1_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(pipe1_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(pipe1_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(pipe1_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(pipe1_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(pipe1_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(pipe1_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(pipe1_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(pipe1_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(pipe1_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(pipe1_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(pipe1_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(pipe1_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(pipe1_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(pipe1_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(pipe1_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(pipe1_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(pipe1_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(pipe1_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(pipe1_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(pipe1_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(pipe1_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(pipe1_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(pipe1_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(pipe1_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(pipe1_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(pipe1_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(pipe1_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(pipe1_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(pipe1_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(pipe1_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(pipe1_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(pipe1_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(pipe1_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(pipe1_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(pipe1_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(pipe1_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(pipe1_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(pipe1_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(pipe1_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(pipe1_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(pipe1_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(pipe1_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(pipe1_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(pipe1_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(pipe1_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(pipe1_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(pipe1_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(pipe1_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(pipe1_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(pipe1_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(pipe1_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(pipe1_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(pipe1_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(pipe1_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(pipe1_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(pipe1_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(pipe1_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(pipe1_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(pipe1_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(pipe1_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(pipe1_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(pipe1_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(pipe1_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(pipe1_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(pipe1_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(pipe1_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(pipe1_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(pipe1_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(pipe1_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(pipe1_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(pipe1_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(pipe1_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(pipe1_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(pipe1_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(pipe1_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(pipe1_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(pipe1_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(pipe1_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(pipe1_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(pipe1_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(pipe1_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(pipe1_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(pipe1_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(pipe1_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(pipe1_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(pipe1_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(pipe1_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(pipe1_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(pipe1_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(pipe1_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(pipe1_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(pipe1_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(pipe1_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(pipe1_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(pipe1_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(pipe1_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(pipe1_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(pipe1_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(pipe1_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(pipe1_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(pipe1_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(pipe1_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(pipe1_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(pipe1_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(pipe1_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(pipe1_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(pipe1_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(pipe1_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(pipe1_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(pipe1_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(pipe1_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(pipe1_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(pipe1_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(pipe1_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(pipe1_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(pipe1_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(pipe1_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(pipe1_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(pipe1_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(pipe1_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(pipe1_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(pipe1_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(pipe1_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(pipe1_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(pipe1_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(pipe1_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(pipe1_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(pipe1_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(pipe1_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(pipe1_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(pipe1_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(pipe1_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(pipe1_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(pipe1_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(pipe1_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(pipe1_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(pipe1_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(pipe1_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(pipe1_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(pipe1_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(pipe1_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(pipe1_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(pipe1_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(pipe1_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(pipe1_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(pipe1_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(pipe1_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(pipe1_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(pipe1_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(pipe1_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(pipe1_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(pipe1_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(pipe1_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(pipe1_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(pipe1_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(pipe1_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(pipe1_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(pipe1_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(pipe1_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(pipe1_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(pipe1_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(pipe1_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(pipe1_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(pipe1_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(pipe1_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(pipe1_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(pipe1_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(pipe1_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(pipe1_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(pipe1_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(pipe1_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(pipe1_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(pipe1_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(pipe1_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(pipe1_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(pipe1_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(pipe1_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(pipe1_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(pipe1_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(pipe1_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(pipe1_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(pipe1_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(pipe1_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(pipe1_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(pipe1_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(pipe1_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(pipe1_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(pipe1_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(pipe1_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(pipe1_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(pipe1_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(pipe1_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(pipe1_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(pipe1_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(pipe1_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(pipe1_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(pipe1_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(pipe1_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(pipe1_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(pipe1_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(pipe1_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(pipe1_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(pipe1_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(pipe1_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(pipe1_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(pipe1_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(pipe1_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(pipe1_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(pipe1_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(pipe1_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(pipe1_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(pipe1_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(pipe1_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(pipe1_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(pipe1_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(pipe1_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(pipe1_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(pipe1_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(pipe1_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(pipe1_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(pipe1_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(pipe1_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(pipe1_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(pipe1_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(pipe1_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(pipe1_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(pipe1_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(pipe1_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(pipe1_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(pipe1_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(pipe1_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(pipe1_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(pipe1_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(pipe1_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(pipe1_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(pipe1_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(pipe1_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(pipe1_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(pipe1_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(pipe1_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(pipe1_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(pipe1_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(pipe1_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(pipe1_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(pipe1_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(pipe1_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(pipe1_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(pipe1_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(pipe1_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(pipe1_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_next_processor_id(pipe1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe1_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe1_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe1_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe1_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe1_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe1_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe1_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe1_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe1_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe1_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe1_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe1_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe1_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe1_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe1_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe1_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe1_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe1_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe1_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe1_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe1_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe1_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe1_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe1_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe1_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe1_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe1_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe1_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe1_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe1_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe1_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe1_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe1_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe1_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe1_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe1_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe1_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe1_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe1_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe1_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe1_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe1_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe1_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe1_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe1_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe1_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe1_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe1_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe1_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe1_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe1_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe1_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe1_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe1_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe1_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe1_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe1_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe1_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe1_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe1_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe1_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe1_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe1_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe1_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe1_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe1_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe1_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe1_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe1_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe1_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe1_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe1_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe1_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe1_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe1_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe1_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe1_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe1_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe1_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe1_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe1_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe1_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe1_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe1_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe1_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe1_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe1_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe1_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe1_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe1_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe1_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe1_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe1_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe1_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe1_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe1_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe1_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe1_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe1_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe1_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe1_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe1_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe1_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe1_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe1_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe1_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe1_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe1_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe1_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe1_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe1_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe1_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe1_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe1_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe1_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe1_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe1_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe1_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe1_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe1_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe1_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe1_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe1_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe1_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe1_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe1_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe1_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe1_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe1_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe1_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe1_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe1_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe1_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe1_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe1_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe1_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe1_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe1_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe1_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe1_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe1_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe1_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe1_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe1_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe1_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe1_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe1_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe1_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe1_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe1_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe1_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe1_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe1_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe1_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe1_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe1_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe1_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe1_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe1_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe1_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe1_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(pipe1_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(pipe1_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(pipe1_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(pipe1_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(pipe1_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(pipe1_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(pipe1_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(pipe1_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(pipe1_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(pipe1_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(pipe1_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(pipe1_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(pipe1_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(pipe1_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(pipe1_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(pipe1_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(pipe1_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(pipe1_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(pipe1_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(pipe1_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(pipe1_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(pipe1_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(pipe1_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(pipe1_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(pipe1_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(pipe1_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(pipe1_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(pipe1_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(pipe1_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(pipe1_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(pipe1_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(pipe1_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(pipe1_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(pipe1_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(pipe1_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(pipe1_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(pipe1_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(pipe1_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(pipe1_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(pipe1_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(pipe1_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(pipe1_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(pipe1_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(pipe1_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(pipe1_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(pipe1_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(pipe1_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(pipe1_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(pipe1_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(pipe1_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(pipe1_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(pipe1_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(pipe1_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(pipe1_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(pipe1_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(pipe1_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(pipe1_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(pipe1_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(pipe1_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(pipe1_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(pipe1_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(pipe1_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(pipe1_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(pipe1_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(pipe1_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(pipe1_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(pipe1_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(pipe1_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(pipe1_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(pipe1_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(pipe1_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(pipe1_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(pipe1_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(pipe1_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(pipe1_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(pipe1_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(pipe1_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(pipe1_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(pipe1_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(pipe1_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(pipe1_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(pipe1_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(pipe1_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(pipe1_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(pipe1_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(pipe1_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(pipe1_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(pipe1_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(pipe1_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(pipe1_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(pipe1_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(pipe1_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(pipe1_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(pipe1_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(pipe1_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(pipe1_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(pipe1_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(pipe1_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(pipe1_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(pipe1_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(pipe1_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(pipe1_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(pipe1_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(pipe1_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(pipe1_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(pipe1_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(pipe1_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(pipe1_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(pipe1_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(pipe1_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(pipe1_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(pipe1_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(pipe1_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(pipe1_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(pipe1_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(pipe1_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(pipe1_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(pipe1_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(pipe1_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(pipe1_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(pipe1_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(pipe1_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(pipe1_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(pipe1_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(pipe1_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(pipe1_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(pipe1_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(pipe1_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(pipe1_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(pipe1_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(pipe1_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(pipe1_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(pipe1_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(pipe1_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(pipe1_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(pipe1_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(pipe1_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(pipe1_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(pipe1_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(pipe1_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(pipe1_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(pipe1_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(pipe1_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(pipe1_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(pipe1_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(pipe1_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(pipe1_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(pipe1_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(pipe1_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(pipe1_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(pipe1_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(pipe1_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(pipe1_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(pipe1_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(pipe1_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(pipe1_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(pipe1_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(pipe1_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(pipe1_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(pipe1_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(pipe1_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(pipe1_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(pipe1_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(pipe1_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(pipe1_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(pipe1_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(pipe1_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(pipe1_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(pipe1_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(pipe1_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(pipe1_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(pipe1_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(pipe1_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(pipe1_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(pipe1_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(pipe1_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(pipe1_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(pipe1_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(pipe1_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(pipe1_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(pipe1_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(pipe1_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(pipe1_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(pipe1_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(pipe1_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(pipe1_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(pipe1_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(pipe1_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(pipe1_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(pipe1_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(pipe1_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(pipe1_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(pipe1_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(pipe1_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(pipe1_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(pipe1_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(pipe1_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(pipe1_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(pipe1_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(pipe1_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(pipe1_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(pipe1_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(pipe1_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(pipe1_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(pipe1_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(pipe1_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(pipe1_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(pipe1_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(pipe1_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(pipe1_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(pipe1_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(pipe1_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(pipe1_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(pipe1_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(pipe1_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(pipe1_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(pipe1_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(pipe1_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(pipe1_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(pipe1_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(pipe1_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(pipe1_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(pipe1_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(pipe1_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(pipe1_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(pipe1_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(pipe1_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(pipe1_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(pipe1_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(pipe1_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(pipe1_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(pipe1_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(pipe1_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(pipe1_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(pipe1_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(pipe1_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(pipe1_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(pipe1_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(pipe1_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(pipe1_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(pipe1_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(pipe1_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(pipe1_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(pipe1_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(pipe1_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(pipe1_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(pipe1_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(pipe1_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(pipe1_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(pipe1_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(pipe1_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(pipe1_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(pipe1_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(pipe1_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(pipe1_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(pipe1_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_next_processor_id(pipe1_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe1_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe1_io_pipe_phv_out_is_valid_processor),
    .io_key_config_0_field_config_0(pipe1_io_key_config_0_field_config_0),
    .io_key_config_0_field_config_1(pipe1_io_key_config_0_field_config_1),
    .io_key_config_0_field_config_2(pipe1_io_key_config_0_field_config_2),
    .io_key_config_0_field_config_3(pipe1_io_key_config_0_field_config_3),
    .io_key_config_0_field_config_4(pipe1_io_key_config_0_field_config_4),
    .io_key_config_0_field_config_5(pipe1_io_key_config_0_field_config_5),
    .io_key_config_0_field_mask_0_0(pipe1_io_key_config_0_field_mask_0_0),
    .io_key_config_0_field_mask_0_1(pipe1_io_key_config_0_field_mask_0_1),
    .io_key_config_0_field_mask_0_2(pipe1_io_key_config_0_field_mask_0_2),
    .io_key_config_0_field_mask_0_3(pipe1_io_key_config_0_field_mask_0_3),
    .io_key_config_0_field_mask_1_0(pipe1_io_key_config_0_field_mask_1_0),
    .io_key_config_0_field_mask_1_1(pipe1_io_key_config_0_field_mask_1_1),
    .io_key_config_0_field_mask_1_2(pipe1_io_key_config_0_field_mask_1_2),
    .io_key_config_0_field_mask_1_3(pipe1_io_key_config_0_field_mask_1_3),
    .io_key_config_0_field_mask_2_0(pipe1_io_key_config_0_field_mask_2_0),
    .io_key_config_0_field_mask_2_1(pipe1_io_key_config_0_field_mask_2_1),
    .io_key_config_0_field_mask_2_2(pipe1_io_key_config_0_field_mask_2_2),
    .io_key_config_0_field_mask_2_3(pipe1_io_key_config_0_field_mask_2_3),
    .io_key_config_0_field_mask_3_0(pipe1_io_key_config_0_field_mask_3_0),
    .io_key_config_0_field_mask_3_1(pipe1_io_key_config_0_field_mask_3_1),
    .io_key_config_0_field_mask_3_2(pipe1_io_key_config_0_field_mask_3_2),
    .io_key_config_0_field_mask_3_3(pipe1_io_key_config_0_field_mask_3_3),
    .io_key_config_0_field_mask_4_0(pipe1_io_key_config_0_field_mask_4_0),
    .io_key_config_0_field_mask_4_1(pipe1_io_key_config_0_field_mask_4_1),
    .io_key_config_0_field_mask_4_2(pipe1_io_key_config_0_field_mask_4_2),
    .io_key_config_0_field_mask_4_3(pipe1_io_key_config_0_field_mask_4_3),
    .io_key_config_0_field_mask_5_0(pipe1_io_key_config_0_field_mask_5_0),
    .io_key_config_0_field_mask_5_1(pipe1_io_key_config_0_field_mask_5_1),
    .io_key_config_0_field_mask_5_2(pipe1_io_key_config_0_field_mask_5_2),
    .io_key_config_0_field_mask_5_3(pipe1_io_key_config_0_field_mask_5_3),
    .io_key_config_0_field_id_0_0(pipe1_io_key_config_0_field_id_0_0),
    .io_key_config_0_field_id_0_1(pipe1_io_key_config_0_field_id_0_1),
    .io_key_config_0_field_id_0_2(pipe1_io_key_config_0_field_id_0_2),
    .io_key_config_0_field_id_0_3(pipe1_io_key_config_0_field_id_0_3),
    .io_key_config_0_field_id_1_0(pipe1_io_key_config_0_field_id_1_0),
    .io_key_config_0_field_id_1_1(pipe1_io_key_config_0_field_id_1_1),
    .io_key_config_0_field_id_1_2(pipe1_io_key_config_0_field_id_1_2),
    .io_key_config_0_field_id_1_3(pipe1_io_key_config_0_field_id_1_3),
    .io_key_config_0_field_id_2_0(pipe1_io_key_config_0_field_id_2_0),
    .io_key_config_0_field_id_2_1(pipe1_io_key_config_0_field_id_2_1),
    .io_key_config_0_field_id_2_2(pipe1_io_key_config_0_field_id_2_2),
    .io_key_config_0_field_id_2_3(pipe1_io_key_config_0_field_id_2_3),
    .io_key_config_0_field_id_3_0(pipe1_io_key_config_0_field_id_3_0),
    .io_key_config_0_field_id_3_1(pipe1_io_key_config_0_field_id_3_1),
    .io_key_config_0_field_id_3_2(pipe1_io_key_config_0_field_id_3_2),
    .io_key_config_0_field_id_3_3(pipe1_io_key_config_0_field_id_3_3),
    .io_key_config_0_field_id_4_0(pipe1_io_key_config_0_field_id_4_0),
    .io_key_config_0_field_id_4_1(pipe1_io_key_config_0_field_id_4_1),
    .io_key_config_0_field_id_4_2(pipe1_io_key_config_0_field_id_4_2),
    .io_key_config_0_field_id_4_3(pipe1_io_key_config_0_field_id_4_3),
    .io_key_config_0_field_id_5_0(pipe1_io_key_config_0_field_id_5_0),
    .io_key_config_0_field_id_5_1(pipe1_io_key_config_0_field_id_5_1),
    .io_key_config_0_field_id_5_2(pipe1_io_key_config_0_field_id_5_2),
    .io_key_config_0_field_id_5_3(pipe1_io_key_config_0_field_id_5_3),
    .io_key_config_1_field_config_0(pipe1_io_key_config_1_field_config_0),
    .io_key_config_1_field_config_1(pipe1_io_key_config_1_field_config_1),
    .io_key_config_1_field_config_2(pipe1_io_key_config_1_field_config_2),
    .io_key_config_1_field_config_3(pipe1_io_key_config_1_field_config_3),
    .io_key_config_1_field_config_4(pipe1_io_key_config_1_field_config_4),
    .io_key_config_1_field_config_5(pipe1_io_key_config_1_field_config_5),
    .io_key_config_1_field_mask_0_0(pipe1_io_key_config_1_field_mask_0_0),
    .io_key_config_1_field_mask_0_1(pipe1_io_key_config_1_field_mask_0_1),
    .io_key_config_1_field_mask_0_2(pipe1_io_key_config_1_field_mask_0_2),
    .io_key_config_1_field_mask_0_3(pipe1_io_key_config_1_field_mask_0_3),
    .io_key_config_1_field_mask_1_0(pipe1_io_key_config_1_field_mask_1_0),
    .io_key_config_1_field_mask_1_1(pipe1_io_key_config_1_field_mask_1_1),
    .io_key_config_1_field_mask_1_2(pipe1_io_key_config_1_field_mask_1_2),
    .io_key_config_1_field_mask_1_3(pipe1_io_key_config_1_field_mask_1_3),
    .io_key_config_1_field_mask_2_0(pipe1_io_key_config_1_field_mask_2_0),
    .io_key_config_1_field_mask_2_1(pipe1_io_key_config_1_field_mask_2_1),
    .io_key_config_1_field_mask_2_2(pipe1_io_key_config_1_field_mask_2_2),
    .io_key_config_1_field_mask_2_3(pipe1_io_key_config_1_field_mask_2_3),
    .io_key_config_1_field_mask_3_0(pipe1_io_key_config_1_field_mask_3_0),
    .io_key_config_1_field_mask_3_1(pipe1_io_key_config_1_field_mask_3_1),
    .io_key_config_1_field_mask_3_2(pipe1_io_key_config_1_field_mask_3_2),
    .io_key_config_1_field_mask_3_3(pipe1_io_key_config_1_field_mask_3_3),
    .io_key_config_1_field_mask_4_0(pipe1_io_key_config_1_field_mask_4_0),
    .io_key_config_1_field_mask_4_1(pipe1_io_key_config_1_field_mask_4_1),
    .io_key_config_1_field_mask_4_2(pipe1_io_key_config_1_field_mask_4_2),
    .io_key_config_1_field_mask_4_3(pipe1_io_key_config_1_field_mask_4_3),
    .io_key_config_1_field_mask_5_0(pipe1_io_key_config_1_field_mask_5_0),
    .io_key_config_1_field_mask_5_1(pipe1_io_key_config_1_field_mask_5_1),
    .io_key_config_1_field_mask_5_2(pipe1_io_key_config_1_field_mask_5_2),
    .io_key_config_1_field_mask_5_3(pipe1_io_key_config_1_field_mask_5_3),
    .io_key_config_1_field_id_0_0(pipe1_io_key_config_1_field_id_0_0),
    .io_key_config_1_field_id_0_1(pipe1_io_key_config_1_field_id_0_1),
    .io_key_config_1_field_id_0_2(pipe1_io_key_config_1_field_id_0_2),
    .io_key_config_1_field_id_0_3(pipe1_io_key_config_1_field_id_0_3),
    .io_key_config_1_field_id_1_0(pipe1_io_key_config_1_field_id_1_0),
    .io_key_config_1_field_id_1_1(pipe1_io_key_config_1_field_id_1_1),
    .io_key_config_1_field_id_1_2(pipe1_io_key_config_1_field_id_1_2),
    .io_key_config_1_field_id_1_3(pipe1_io_key_config_1_field_id_1_3),
    .io_key_config_1_field_id_2_0(pipe1_io_key_config_1_field_id_2_0),
    .io_key_config_1_field_id_2_1(pipe1_io_key_config_1_field_id_2_1),
    .io_key_config_1_field_id_2_2(pipe1_io_key_config_1_field_id_2_2),
    .io_key_config_1_field_id_2_3(pipe1_io_key_config_1_field_id_2_3),
    .io_key_config_1_field_id_3_0(pipe1_io_key_config_1_field_id_3_0),
    .io_key_config_1_field_id_3_1(pipe1_io_key_config_1_field_id_3_1),
    .io_key_config_1_field_id_3_2(pipe1_io_key_config_1_field_id_3_2),
    .io_key_config_1_field_id_3_3(pipe1_io_key_config_1_field_id_3_3),
    .io_key_config_1_field_id_4_0(pipe1_io_key_config_1_field_id_4_0),
    .io_key_config_1_field_id_4_1(pipe1_io_key_config_1_field_id_4_1),
    .io_key_config_1_field_id_4_2(pipe1_io_key_config_1_field_id_4_2),
    .io_key_config_1_field_id_4_3(pipe1_io_key_config_1_field_id_4_3),
    .io_key_config_1_field_id_5_0(pipe1_io_key_config_1_field_id_5_0),
    .io_key_config_1_field_id_5_1(pipe1_io_key_config_1_field_id_5_1),
    .io_key_config_1_field_id_5_2(pipe1_io_key_config_1_field_id_5_2),
    .io_key_config_1_field_id_5_3(pipe1_io_key_config_1_field_id_5_3),
    .io_match_key(pipe1_io_match_key)
  );
  Hash pipe2 ( // @[matcher_pisa.scala 334:23]
    .clock(pipe2_clock),
    .io_pipe_phv_in_data_0(pipe2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe2_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe2_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe2_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe2_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe2_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe2_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe2_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe2_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe2_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe2_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe2_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe2_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe2_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe2_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe2_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe2_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe2_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe2_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe2_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe2_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe2_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe2_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe2_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe2_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe2_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe2_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe2_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe2_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe2_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe2_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe2_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe2_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe2_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe2_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe2_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe2_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe2_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe2_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe2_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe2_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe2_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe2_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe2_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe2_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe2_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe2_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe2_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe2_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe2_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe2_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe2_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe2_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe2_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe2_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe2_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe2_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe2_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe2_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe2_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe2_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe2_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe2_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe2_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe2_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe2_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe2_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe2_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe2_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe2_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe2_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe2_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe2_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe2_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe2_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe2_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe2_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe2_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe2_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe2_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe2_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe2_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe2_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe2_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe2_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe2_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe2_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe2_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe2_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe2_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe2_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe2_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe2_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe2_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe2_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe2_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe2_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe2_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe2_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe2_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe2_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe2_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe2_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe2_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe2_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe2_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe2_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe2_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe2_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe2_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe2_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe2_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe2_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe2_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe2_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe2_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe2_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe2_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe2_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe2_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe2_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe2_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe2_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe2_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe2_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe2_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe2_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe2_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe2_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe2_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe2_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe2_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe2_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe2_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe2_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe2_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe2_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe2_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe2_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe2_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe2_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe2_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe2_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe2_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe2_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe2_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe2_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe2_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe2_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe2_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe2_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe2_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe2_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe2_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe2_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe2_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe2_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe2_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe2_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe2_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe2_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(pipe2_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(pipe2_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(pipe2_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(pipe2_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(pipe2_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(pipe2_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(pipe2_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(pipe2_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(pipe2_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(pipe2_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(pipe2_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(pipe2_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(pipe2_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(pipe2_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(pipe2_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(pipe2_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(pipe2_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(pipe2_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(pipe2_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(pipe2_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(pipe2_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(pipe2_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(pipe2_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(pipe2_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(pipe2_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(pipe2_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(pipe2_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(pipe2_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(pipe2_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(pipe2_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(pipe2_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(pipe2_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(pipe2_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(pipe2_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(pipe2_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(pipe2_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(pipe2_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(pipe2_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(pipe2_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(pipe2_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(pipe2_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(pipe2_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(pipe2_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(pipe2_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(pipe2_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(pipe2_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(pipe2_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(pipe2_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(pipe2_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(pipe2_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(pipe2_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(pipe2_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(pipe2_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(pipe2_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(pipe2_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(pipe2_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(pipe2_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(pipe2_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(pipe2_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(pipe2_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(pipe2_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(pipe2_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(pipe2_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(pipe2_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(pipe2_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(pipe2_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(pipe2_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(pipe2_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(pipe2_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(pipe2_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(pipe2_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(pipe2_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(pipe2_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(pipe2_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(pipe2_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(pipe2_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(pipe2_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(pipe2_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(pipe2_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(pipe2_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(pipe2_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(pipe2_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(pipe2_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(pipe2_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(pipe2_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(pipe2_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(pipe2_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(pipe2_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(pipe2_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(pipe2_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(pipe2_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(pipe2_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(pipe2_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(pipe2_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(pipe2_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(pipe2_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(pipe2_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(pipe2_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(pipe2_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(pipe2_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(pipe2_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(pipe2_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(pipe2_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(pipe2_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(pipe2_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(pipe2_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(pipe2_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(pipe2_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(pipe2_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(pipe2_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(pipe2_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(pipe2_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(pipe2_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(pipe2_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(pipe2_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(pipe2_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(pipe2_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(pipe2_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(pipe2_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(pipe2_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(pipe2_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(pipe2_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(pipe2_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(pipe2_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(pipe2_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(pipe2_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(pipe2_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(pipe2_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(pipe2_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(pipe2_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(pipe2_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(pipe2_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(pipe2_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(pipe2_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(pipe2_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(pipe2_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(pipe2_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(pipe2_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(pipe2_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(pipe2_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(pipe2_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(pipe2_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(pipe2_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(pipe2_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(pipe2_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(pipe2_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(pipe2_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(pipe2_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(pipe2_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(pipe2_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(pipe2_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(pipe2_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(pipe2_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(pipe2_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(pipe2_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(pipe2_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(pipe2_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(pipe2_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(pipe2_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(pipe2_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(pipe2_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(pipe2_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(pipe2_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(pipe2_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(pipe2_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(pipe2_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(pipe2_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(pipe2_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(pipe2_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(pipe2_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(pipe2_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(pipe2_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(pipe2_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(pipe2_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(pipe2_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(pipe2_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(pipe2_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(pipe2_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(pipe2_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(pipe2_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(pipe2_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(pipe2_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(pipe2_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(pipe2_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(pipe2_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(pipe2_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(pipe2_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(pipe2_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(pipe2_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(pipe2_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(pipe2_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(pipe2_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(pipe2_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(pipe2_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(pipe2_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(pipe2_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(pipe2_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(pipe2_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(pipe2_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(pipe2_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(pipe2_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(pipe2_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(pipe2_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(pipe2_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(pipe2_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(pipe2_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(pipe2_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(pipe2_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(pipe2_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(pipe2_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(pipe2_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(pipe2_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(pipe2_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(pipe2_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(pipe2_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(pipe2_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(pipe2_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(pipe2_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(pipe2_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(pipe2_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(pipe2_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(pipe2_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(pipe2_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(pipe2_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(pipe2_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(pipe2_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(pipe2_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(pipe2_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(pipe2_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(pipe2_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(pipe2_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(pipe2_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(pipe2_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(pipe2_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(pipe2_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(pipe2_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(pipe2_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(pipe2_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(pipe2_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(pipe2_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(pipe2_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(pipe2_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(pipe2_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(pipe2_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(pipe2_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(pipe2_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(pipe2_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(pipe2_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(pipe2_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(pipe2_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(pipe2_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(pipe2_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(pipe2_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(pipe2_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(pipe2_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(pipe2_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_next_processor_id(pipe2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe2_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe2_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe2_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe2_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe2_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe2_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe2_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe2_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe2_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe2_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe2_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe2_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe2_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe2_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe2_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe2_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe2_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe2_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe2_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe2_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe2_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe2_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe2_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe2_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe2_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe2_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe2_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe2_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe2_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe2_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe2_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe2_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe2_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe2_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe2_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe2_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe2_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe2_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe2_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe2_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe2_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe2_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe2_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe2_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe2_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe2_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe2_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe2_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe2_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe2_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe2_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe2_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe2_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe2_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe2_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe2_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe2_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe2_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe2_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe2_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe2_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe2_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe2_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe2_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe2_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe2_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe2_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe2_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe2_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe2_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe2_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe2_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe2_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe2_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe2_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe2_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe2_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe2_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe2_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe2_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe2_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe2_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe2_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe2_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe2_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe2_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe2_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe2_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe2_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe2_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe2_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe2_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe2_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe2_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe2_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe2_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe2_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe2_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe2_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe2_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe2_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe2_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe2_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe2_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe2_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe2_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe2_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe2_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe2_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe2_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe2_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe2_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe2_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe2_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe2_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe2_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe2_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe2_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe2_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe2_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe2_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe2_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe2_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe2_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe2_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe2_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe2_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe2_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe2_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe2_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe2_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe2_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe2_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe2_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe2_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe2_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe2_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe2_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe2_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe2_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe2_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe2_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe2_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe2_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe2_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe2_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe2_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe2_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe2_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe2_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe2_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe2_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe2_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe2_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe2_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe2_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe2_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe2_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe2_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe2_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe2_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(pipe2_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(pipe2_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(pipe2_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(pipe2_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(pipe2_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(pipe2_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(pipe2_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(pipe2_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(pipe2_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(pipe2_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(pipe2_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(pipe2_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(pipe2_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(pipe2_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(pipe2_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(pipe2_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(pipe2_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(pipe2_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(pipe2_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(pipe2_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(pipe2_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(pipe2_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(pipe2_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(pipe2_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(pipe2_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(pipe2_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(pipe2_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(pipe2_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(pipe2_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(pipe2_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(pipe2_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(pipe2_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(pipe2_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(pipe2_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(pipe2_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(pipe2_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(pipe2_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(pipe2_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(pipe2_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(pipe2_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(pipe2_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(pipe2_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(pipe2_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(pipe2_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(pipe2_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(pipe2_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(pipe2_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(pipe2_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(pipe2_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(pipe2_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(pipe2_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(pipe2_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(pipe2_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(pipe2_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(pipe2_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(pipe2_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(pipe2_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(pipe2_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(pipe2_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(pipe2_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(pipe2_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(pipe2_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(pipe2_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(pipe2_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(pipe2_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(pipe2_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(pipe2_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(pipe2_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(pipe2_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(pipe2_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(pipe2_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(pipe2_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(pipe2_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(pipe2_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(pipe2_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(pipe2_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(pipe2_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(pipe2_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(pipe2_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(pipe2_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(pipe2_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(pipe2_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(pipe2_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(pipe2_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(pipe2_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(pipe2_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(pipe2_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(pipe2_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(pipe2_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(pipe2_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(pipe2_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(pipe2_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(pipe2_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(pipe2_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(pipe2_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(pipe2_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(pipe2_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(pipe2_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(pipe2_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(pipe2_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(pipe2_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(pipe2_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(pipe2_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(pipe2_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(pipe2_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(pipe2_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(pipe2_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(pipe2_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(pipe2_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(pipe2_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(pipe2_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(pipe2_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(pipe2_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(pipe2_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(pipe2_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(pipe2_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(pipe2_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(pipe2_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(pipe2_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(pipe2_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(pipe2_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(pipe2_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(pipe2_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(pipe2_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(pipe2_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(pipe2_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(pipe2_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(pipe2_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(pipe2_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(pipe2_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(pipe2_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(pipe2_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(pipe2_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(pipe2_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(pipe2_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(pipe2_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(pipe2_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(pipe2_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(pipe2_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(pipe2_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(pipe2_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(pipe2_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(pipe2_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(pipe2_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(pipe2_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(pipe2_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(pipe2_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(pipe2_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(pipe2_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(pipe2_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(pipe2_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(pipe2_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(pipe2_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(pipe2_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(pipe2_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(pipe2_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(pipe2_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(pipe2_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(pipe2_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(pipe2_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(pipe2_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(pipe2_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(pipe2_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(pipe2_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(pipe2_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(pipe2_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(pipe2_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(pipe2_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(pipe2_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(pipe2_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(pipe2_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(pipe2_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(pipe2_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(pipe2_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(pipe2_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(pipe2_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(pipe2_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(pipe2_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(pipe2_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(pipe2_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(pipe2_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(pipe2_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(pipe2_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(pipe2_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(pipe2_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(pipe2_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(pipe2_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(pipe2_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(pipe2_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(pipe2_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(pipe2_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(pipe2_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(pipe2_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(pipe2_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(pipe2_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(pipe2_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(pipe2_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(pipe2_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(pipe2_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(pipe2_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(pipe2_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(pipe2_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(pipe2_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(pipe2_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(pipe2_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(pipe2_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(pipe2_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(pipe2_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(pipe2_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(pipe2_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(pipe2_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(pipe2_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(pipe2_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(pipe2_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(pipe2_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(pipe2_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(pipe2_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(pipe2_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(pipe2_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(pipe2_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(pipe2_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(pipe2_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(pipe2_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(pipe2_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(pipe2_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(pipe2_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(pipe2_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(pipe2_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(pipe2_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(pipe2_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(pipe2_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(pipe2_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(pipe2_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(pipe2_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(pipe2_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(pipe2_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(pipe2_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(pipe2_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(pipe2_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(pipe2_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(pipe2_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(pipe2_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(pipe2_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(pipe2_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(pipe2_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(pipe2_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(pipe2_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(pipe2_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(pipe2_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(pipe2_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(pipe2_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(pipe2_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(pipe2_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(pipe2_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(pipe2_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(pipe2_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_next_processor_id(pipe2_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe2_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe2_io_pipe_phv_out_is_valid_processor),
    .io_mod_hash_depth_mod(pipe2_io_mod_hash_depth_mod),
    .io_mod_config_id(pipe2_io_mod_config_id),
    .io_mod_hash_depth(pipe2_io_mod_hash_depth),
    .io_key_in(pipe2_io_key_in),
    .io_key_out(pipe2_io_key_out),
    .io_hash_val(pipe2_io_hash_val),
    .io_hash_val_cs(pipe2_io_hash_val_cs)
  );
  MatchReadDataPISA pipe3 ( // @[matcher_pisa.scala 335:23]
    .clock(pipe3_clock),
    .io_pipe_phv_in_data_0(pipe3_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe3_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe3_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe3_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe3_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe3_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe3_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe3_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe3_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe3_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe3_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe3_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe3_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe3_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe3_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe3_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe3_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe3_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe3_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe3_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe3_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe3_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe3_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe3_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe3_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe3_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe3_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe3_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe3_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe3_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe3_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe3_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe3_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe3_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe3_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe3_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe3_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe3_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe3_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe3_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe3_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe3_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe3_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe3_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe3_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe3_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe3_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe3_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe3_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe3_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe3_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe3_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe3_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe3_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe3_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe3_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe3_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe3_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe3_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe3_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe3_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe3_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe3_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe3_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe3_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe3_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe3_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe3_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe3_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe3_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe3_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe3_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe3_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe3_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe3_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe3_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe3_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe3_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe3_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe3_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe3_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe3_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe3_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe3_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe3_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe3_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe3_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe3_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe3_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe3_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe3_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe3_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe3_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe3_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe3_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe3_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe3_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe3_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe3_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe3_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe3_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe3_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe3_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe3_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe3_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe3_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe3_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe3_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe3_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe3_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe3_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe3_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe3_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe3_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe3_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe3_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe3_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe3_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe3_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe3_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe3_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe3_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe3_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe3_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe3_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe3_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe3_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe3_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe3_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe3_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe3_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe3_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe3_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe3_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe3_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe3_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe3_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe3_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe3_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe3_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe3_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe3_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe3_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe3_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe3_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe3_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe3_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe3_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe3_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe3_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe3_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe3_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe3_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe3_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe3_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe3_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe3_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe3_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe3_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe3_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe3_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe3_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe3_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe3_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe3_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe3_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe3_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe3_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe3_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe3_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe3_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe3_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe3_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe3_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe3_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe3_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe3_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe3_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe3_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe3_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe3_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe3_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe3_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe3_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe3_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe3_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe3_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe3_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe3_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe3_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe3_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe3_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe3_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe3_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe3_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe3_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe3_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe3_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe3_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe3_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe3_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe3_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe3_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe3_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe3_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe3_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe3_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe3_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe3_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe3_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe3_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe3_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe3_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe3_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe3_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe3_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe3_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe3_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe3_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe3_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe3_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe3_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe3_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe3_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe3_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe3_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe3_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe3_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe3_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe3_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe3_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe3_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe3_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe3_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe3_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe3_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe3_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe3_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe3_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe3_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe3_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe3_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe3_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe3_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe3_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe3_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe3_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe3_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe3_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe3_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe3_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe3_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe3_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe3_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe3_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe3_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(pipe3_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(pipe3_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(pipe3_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(pipe3_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(pipe3_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(pipe3_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(pipe3_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(pipe3_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(pipe3_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(pipe3_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(pipe3_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(pipe3_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(pipe3_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(pipe3_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(pipe3_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(pipe3_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(pipe3_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(pipe3_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(pipe3_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(pipe3_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(pipe3_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(pipe3_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(pipe3_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(pipe3_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(pipe3_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(pipe3_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(pipe3_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(pipe3_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(pipe3_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(pipe3_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(pipe3_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(pipe3_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(pipe3_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(pipe3_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(pipe3_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(pipe3_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(pipe3_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(pipe3_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(pipe3_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(pipe3_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(pipe3_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(pipe3_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(pipe3_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(pipe3_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(pipe3_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(pipe3_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(pipe3_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(pipe3_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(pipe3_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(pipe3_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(pipe3_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(pipe3_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(pipe3_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(pipe3_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(pipe3_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(pipe3_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(pipe3_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(pipe3_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(pipe3_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(pipe3_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(pipe3_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(pipe3_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(pipe3_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(pipe3_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(pipe3_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(pipe3_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(pipe3_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(pipe3_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(pipe3_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(pipe3_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(pipe3_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(pipe3_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(pipe3_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(pipe3_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(pipe3_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(pipe3_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(pipe3_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(pipe3_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(pipe3_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(pipe3_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(pipe3_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(pipe3_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(pipe3_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(pipe3_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(pipe3_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(pipe3_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(pipe3_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(pipe3_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(pipe3_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(pipe3_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(pipe3_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(pipe3_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(pipe3_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(pipe3_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(pipe3_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(pipe3_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(pipe3_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(pipe3_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(pipe3_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(pipe3_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(pipe3_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(pipe3_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(pipe3_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(pipe3_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(pipe3_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(pipe3_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(pipe3_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(pipe3_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(pipe3_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(pipe3_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(pipe3_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(pipe3_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(pipe3_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(pipe3_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(pipe3_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(pipe3_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(pipe3_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(pipe3_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(pipe3_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(pipe3_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(pipe3_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(pipe3_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(pipe3_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(pipe3_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(pipe3_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(pipe3_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(pipe3_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(pipe3_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(pipe3_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(pipe3_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(pipe3_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(pipe3_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(pipe3_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(pipe3_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(pipe3_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(pipe3_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(pipe3_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(pipe3_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(pipe3_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(pipe3_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(pipe3_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(pipe3_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(pipe3_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(pipe3_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(pipe3_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(pipe3_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(pipe3_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(pipe3_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(pipe3_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(pipe3_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(pipe3_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(pipe3_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(pipe3_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(pipe3_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(pipe3_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(pipe3_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(pipe3_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(pipe3_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(pipe3_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(pipe3_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(pipe3_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(pipe3_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(pipe3_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(pipe3_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(pipe3_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(pipe3_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(pipe3_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(pipe3_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(pipe3_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(pipe3_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(pipe3_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(pipe3_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(pipe3_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(pipe3_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(pipe3_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(pipe3_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(pipe3_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(pipe3_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(pipe3_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(pipe3_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(pipe3_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(pipe3_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(pipe3_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(pipe3_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(pipe3_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(pipe3_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(pipe3_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(pipe3_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(pipe3_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(pipe3_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(pipe3_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(pipe3_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(pipe3_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(pipe3_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(pipe3_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(pipe3_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(pipe3_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(pipe3_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(pipe3_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(pipe3_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(pipe3_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(pipe3_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(pipe3_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(pipe3_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(pipe3_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(pipe3_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(pipe3_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(pipe3_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(pipe3_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(pipe3_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(pipe3_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(pipe3_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(pipe3_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(pipe3_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(pipe3_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(pipe3_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(pipe3_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(pipe3_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(pipe3_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(pipe3_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(pipe3_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(pipe3_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(pipe3_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(pipe3_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(pipe3_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(pipe3_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(pipe3_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(pipe3_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(pipe3_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(pipe3_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(pipe3_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(pipe3_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(pipe3_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(pipe3_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(pipe3_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(pipe3_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(pipe3_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(pipe3_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(pipe3_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(pipe3_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(pipe3_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(pipe3_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(pipe3_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(pipe3_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(pipe3_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(pipe3_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(pipe3_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(pipe3_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(pipe3_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(pipe3_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(pipe3_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(pipe3_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(pipe3_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(pipe3_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(pipe3_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(pipe3_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_next_processor_id(pipe3_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe3_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe3_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe3_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe3_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe3_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe3_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe3_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe3_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe3_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe3_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe3_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe3_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe3_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe3_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe3_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe3_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe3_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe3_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe3_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe3_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe3_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe3_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe3_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe3_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe3_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe3_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe3_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe3_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe3_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe3_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe3_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe3_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe3_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe3_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe3_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe3_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe3_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe3_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe3_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe3_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe3_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe3_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe3_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe3_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe3_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe3_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe3_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe3_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe3_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe3_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe3_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe3_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe3_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe3_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe3_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe3_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe3_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe3_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe3_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe3_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe3_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe3_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe3_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe3_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe3_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe3_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe3_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe3_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe3_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe3_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe3_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe3_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe3_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe3_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe3_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe3_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe3_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe3_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe3_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe3_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe3_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe3_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe3_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe3_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe3_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe3_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe3_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe3_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe3_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe3_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe3_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe3_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe3_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe3_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe3_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe3_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe3_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe3_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe3_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe3_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe3_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe3_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe3_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe3_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe3_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe3_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe3_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe3_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe3_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe3_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe3_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe3_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe3_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe3_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe3_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe3_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe3_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe3_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe3_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe3_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe3_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe3_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe3_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe3_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe3_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe3_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe3_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe3_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe3_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe3_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe3_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe3_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe3_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe3_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe3_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe3_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe3_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe3_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe3_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe3_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe3_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe3_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe3_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe3_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe3_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe3_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe3_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe3_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe3_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe3_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe3_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe3_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe3_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe3_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe3_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe3_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe3_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe3_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe3_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe3_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe3_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe3_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe3_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe3_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe3_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe3_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe3_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe3_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe3_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe3_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe3_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe3_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe3_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe3_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe3_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe3_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe3_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe3_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe3_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe3_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe3_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe3_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe3_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe3_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe3_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe3_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe3_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe3_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe3_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe3_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe3_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe3_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe3_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe3_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe3_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe3_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe3_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe3_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe3_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe3_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe3_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe3_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe3_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe3_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe3_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe3_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe3_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe3_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe3_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe3_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe3_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe3_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe3_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe3_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe3_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe3_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe3_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe3_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe3_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe3_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe3_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe3_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe3_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe3_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe3_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe3_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe3_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe3_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe3_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe3_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe3_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe3_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe3_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe3_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe3_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe3_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe3_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe3_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe3_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe3_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe3_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe3_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe3_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe3_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe3_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe3_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe3_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe3_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe3_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe3_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe3_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe3_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe3_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe3_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe3_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe3_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe3_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe3_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(pipe3_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(pipe3_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(pipe3_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(pipe3_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(pipe3_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(pipe3_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(pipe3_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(pipe3_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(pipe3_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(pipe3_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(pipe3_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(pipe3_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(pipe3_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(pipe3_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(pipe3_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(pipe3_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(pipe3_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(pipe3_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(pipe3_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(pipe3_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(pipe3_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(pipe3_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(pipe3_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(pipe3_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(pipe3_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(pipe3_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(pipe3_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(pipe3_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(pipe3_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(pipe3_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(pipe3_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(pipe3_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(pipe3_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(pipe3_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(pipe3_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(pipe3_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(pipe3_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(pipe3_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(pipe3_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(pipe3_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(pipe3_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(pipe3_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(pipe3_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(pipe3_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(pipe3_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(pipe3_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(pipe3_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(pipe3_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(pipe3_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(pipe3_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(pipe3_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(pipe3_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(pipe3_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(pipe3_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(pipe3_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(pipe3_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(pipe3_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(pipe3_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(pipe3_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(pipe3_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(pipe3_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(pipe3_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(pipe3_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(pipe3_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(pipe3_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(pipe3_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(pipe3_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(pipe3_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(pipe3_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(pipe3_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(pipe3_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(pipe3_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(pipe3_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(pipe3_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(pipe3_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(pipe3_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(pipe3_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(pipe3_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(pipe3_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(pipe3_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(pipe3_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(pipe3_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(pipe3_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(pipe3_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(pipe3_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(pipe3_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(pipe3_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(pipe3_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(pipe3_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(pipe3_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(pipe3_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(pipe3_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(pipe3_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(pipe3_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(pipe3_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(pipe3_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(pipe3_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(pipe3_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(pipe3_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(pipe3_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(pipe3_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(pipe3_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(pipe3_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(pipe3_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(pipe3_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(pipe3_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(pipe3_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(pipe3_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(pipe3_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(pipe3_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(pipe3_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(pipe3_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(pipe3_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(pipe3_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(pipe3_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(pipe3_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(pipe3_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(pipe3_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(pipe3_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(pipe3_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(pipe3_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(pipe3_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(pipe3_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(pipe3_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(pipe3_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(pipe3_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(pipe3_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(pipe3_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(pipe3_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(pipe3_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(pipe3_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(pipe3_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(pipe3_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(pipe3_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(pipe3_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(pipe3_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(pipe3_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(pipe3_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(pipe3_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(pipe3_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(pipe3_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(pipe3_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(pipe3_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(pipe3_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(pipe3_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(pipe3_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(pipe3_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(pipe3_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(pipe3_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(pipe3_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(pipe3_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(pipe3_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(pipe3_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(pipe3_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(pipe3_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(pipe3_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(pipe3_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(pipe3_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(pipe3_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(pipe3_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(pipe3_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(pipe3_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(pipe3_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(pipe3_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(pipe3_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(pipe3_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(pipe3_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(pipe3_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(pipe3_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(pipe3_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(pipe3_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(pipe3_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(pipe3_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(pipe3_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(pipe3_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(pipe3_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(pipe3_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(pipe3_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(pipe3_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(pipe3_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(pipe3_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(pipe3_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(pipe3_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(pipe3_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(pipe3_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(pipe3_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(pipe3_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(pipe3_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(pipe3_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(pipe3_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(pipe3_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(pipe3_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(pipe3_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(pipe3_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(pipe3_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(pipe3_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(pipe3_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(pipe3_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(pipe3_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(pipe3_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(pipe3_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(pipe3_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(pipe3_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(pipe3_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(pipe3_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(pipe3_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(pipe3_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(pipe3_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(pipe3_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(pipe3_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(pipe3_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(pipe3_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(pipe3_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(pipe3_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(pipe3_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(pipe3_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(pipe3_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(pipe3_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(pipe3_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(pipe3_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(pipe3_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(pipe3_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(pipe3_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(pipe3_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(pipe3_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(pipe3_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(pipe3_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(pipe3_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(pipe3_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(pipe3_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(pipe3_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(pipe3_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(pipe3_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(pipe3_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(pipe3_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(pipe3_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(pipe3_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(pipe3_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(pipe3_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(pipe3_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(pipe3_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(pipe3_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(pipe3_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(pipe3_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(pipe3_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(pipe3_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(pipe3_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(pipe3_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(pipe3_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(pipe3_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(pipe3_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(pipe3_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(pipe3_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(pipe3_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(pipe3_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(pipe3_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_next_processor_id(pipe3_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe3_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe3_io_pipe_phv_out_is_valid_processor),
    .io_table_config_0_table_depth(pipe3_io_table_config_0_table_depth),
    .io_table_config_0_table_width(pipe3_io_table_config_0_table_width),
    .io_table_config_1_table_depth(pipe3_io_table_config_1_table_depth),
    .io_table_config_1_table_width(pipe3_io_table_config_1_table_width),
    .io_key_in(pipe3_io_key_in),
    .io_key_out(pipe3_io_key_out),
    .io_addr_in(pipe3_io_addr_in),
    .io_cs_in(pipe3_io_cs_in),
    .io_data_out(pipe3_io_data_out),
    .io_w_en(pipe3_io_w_en),
    .io_w_sram_id(pipe3_io_w_sram_id),
    .io_w_addr(pipe3_io_w_addr),
    .io_w_data(pipe3_io_w_data)
  );
  MatchResultPISA pipe4 ( // @[matcher_pisa.scala 336:23]
    .clock(pipe4_clock),
    .io_pipe_phv_in_data_0(pipe4_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe4_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe4_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe4_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe4_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe4_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe4_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe4_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe4_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe4_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe4_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe4_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe4_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe4_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe4_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe4_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe4_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe4_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe4_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe4_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe4_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe4_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe4_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe4_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe4_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe4_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe4_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe4_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe4_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe4_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe4_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe4_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe4_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe4_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe4_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe4_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe4_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe4_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe4_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe4_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe4_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe4_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe4_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe4_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe4_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe4_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe4_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe4_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe4_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe4_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe4_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe4_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe4_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe4_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe4_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe4_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe4_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe4_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe4_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe4_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe4_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe4_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe4_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe4_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe4_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe4_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe4_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe4_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe4_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe4_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe4_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe4_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe4_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe4_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe4_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe4_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe4_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe4_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe4_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe4_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe4_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe4_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe4_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe4_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe4_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe4_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe4_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe4_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe4_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe4_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe4_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe4_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe4_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe4_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe4_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe4_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe4_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe4_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe4_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe4_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe4_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe4_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe4_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe4_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe4_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe4_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe4_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe4_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe4_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe4_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe4_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe4_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe4_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe4_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe4_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe4_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe4_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe4_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe4_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe4_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe4_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe4_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe4_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe4_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe4_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe4_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe4_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe4_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe4_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe4_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe4_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe4_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe4_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe4_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe4_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe4_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe4_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe4_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe4_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe4_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe4_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe4_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe4_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe4_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe4_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe4_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe4_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe4_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe4_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe4_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe4_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe4_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe4_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe4_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe4_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe4_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe4_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe4_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe4_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe4_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe4_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe4_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe4_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe4_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe4_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe4_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe4_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe4_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe4_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe4_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe4_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe4_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe4_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe4_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe4_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe4_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe4_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe4_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe4_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe4_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe4_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe4_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe4_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe4_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe4_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe4_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe4_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe4_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe4_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe4_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe4_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe4_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe4_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe4_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe4_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe4_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe4_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe4_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe4_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe4_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe4_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe4_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe4_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe4_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe4_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe4_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe4_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe4_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe4_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe4_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe4_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe4_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe4_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe4_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe4_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe4_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe4_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe4_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe4_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe4_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe4_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe4_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe4_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe4_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe4_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe4_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe4_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe4_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe4_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe4_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe4_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe4_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe4_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe4_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe4_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe4_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe4_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe4_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe4_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe4_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe4_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe4_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe4_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe4_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe4_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe4_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe4_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe4_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe4_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe4_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe4_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe4_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe4_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe4_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe4_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe4_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(pipe4_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(pipe4_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(pipe4_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(pipe4_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(pipe4_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(pipe4_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(pipe4_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(pipe4_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(pipe4_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(pipe4_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(pipe4_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(pipe4_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(pipe4_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(pipe4_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(pipe4_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(pipe4_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(pipe4_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(pipe4_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(pipe4_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(pipe4_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(pipe4_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(pipe4_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(pipe4_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(pipe4_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(pipe4_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(pipe4_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(pipe4_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(pipe4_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(pipe4_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(pipe4_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(pipe4_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(pipe4_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(pipe4_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(pipe4_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(pipe4_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(pipe4_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(pipe4_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(pipe4_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(pipe4_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(pipe4_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(pipe4_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(pipe4_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(pipe4_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(pipe4_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(pipe4_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(pipe4_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(pipe4_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(pipe4_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(pipe4_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(pipe4_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(pipe4_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(pipe4_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(pipe4_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(pipe4_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(pipe4_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(pipe4_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(pipe4_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(pipe4_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(pipe4_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(pipe4_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(pipe4_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(pipe4_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(pipe4_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(pipe4_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(pipe4_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(pipe4_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(pipe4_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(pipe4_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(pipe4_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(pipe4_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(pipe4_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(pipe4_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(pipe4_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(pipe4_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(pipe4_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(pipe4_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(pipe4_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(pipe4_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(pipe4_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(pipe4_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(pipe4_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(pipe4_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(pipe4_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(pipe4_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(pipe4_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(pipe4_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(pipe4_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(pipe4_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(pipe4_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(pipe4_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(pipe4_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(pipe4_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(pipe4_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(pipe4_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(pipe4_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(pipe4_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(pipe4_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(pipe4_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(pipe4_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(pipe4_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(pipe4_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(pipe4_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(pipe4_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(pipe4_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(pipe4_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(pipe4_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(pipe4_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(pipe4_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(pipe4_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(pipe4_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(pipe4_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(pipe4_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(pipe4_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(pipe4_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(pipe4_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(pipe4_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(pipe4_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(pipe4_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(pipe4_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(pipe4_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(pipe4_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(pipe4_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(pipe4_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(pipe4_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(pipe4_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(pipe4_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(pipe4_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(pipe4_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(pipe4_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(pipe4_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(pipe4_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(pipe4_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(pipe4_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(pipe4_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(pipe4_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(pipe4_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(pipe4_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(pipe4_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(pipe4_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(pipe4_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(pipe4_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(pipe4_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(pipe4_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(pipe4_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(pipe4_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(pipe4_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(pipe4_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(pipe4_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(pipe4_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(pipe4_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(pipe4_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(pipe4_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(pipe4_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(pipe4_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(pipe4_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(pipe4_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(pipe4_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(pipe4_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(pipe4_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(pipe4_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(pipe4_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(pipe4_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(pipe4_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(pipe4_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(pipe4_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(pipe4_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(pipe4_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(pipe4_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(pipe4_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(pipe4_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(pipe4_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(pipe4_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(pipe4_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(pipe4_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(pipe4_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(pipe4_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(pipe4_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(pipe4_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(pipe4_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(pipe4_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(pipe4_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(pipe4_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(pipe4_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(pipe4_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(pipe4_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(pipe4_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(pipe4_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(pipe4_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(pipe4_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(pipe4_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(pipe4_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(pipe4_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(pipe4_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(pipe4_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(pipe4_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(pipe4_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(pipe4_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(pipe4_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(pipe4_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(pipe4_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(pipe4_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(pipe4_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(pipe4_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(pipe4_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(pipe4_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(pipe4_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(pipe4_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(pipe4_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(pipe4_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(pipe4_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(pipe4_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(pipe4_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(pipe4_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(pipe4_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(pipe4_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(pipe4_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(pipe4_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(pipe4_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(pipe4_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(pipe4_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(pipe4_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(pipe4_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(pipe4_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(pipe4_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(pipe4_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(pipe4_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(pipe4_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(pipe4_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(pipe4_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(pipe4_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(pipe4_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(pipe4_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(pipe4_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(pipe4_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(pipe4_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(pipe4_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(pipe4_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(pipe4_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(pipe4_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(pipe4_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(pipe4_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(pipe4_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(pipe4_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(pipe4_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(pipe4_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(pipe4_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(pipe4_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(pipe4_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(pipe4_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(pipe4_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(pipe4_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(pipe4_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(pipe4_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(pipe4_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(pipe4_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(pipe4_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_next_processor_id(pipe4_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe4_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe4_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe4_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe4_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe4_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe4_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe4_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe4_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe4_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe4_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe4_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe4_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe4_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe4_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe4_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe4_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe4_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe4_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe4_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe4_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe4_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe4_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe4_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe4_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe4_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe4_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe4_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe4_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe4_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe4_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe4_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe4_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe4_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe4_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe4_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe4_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe4_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe4_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe4_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe4_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe4_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe4_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe4_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe4_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe4_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe4_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe4_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe4_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe4_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe4_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe4_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe4_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe4_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe4_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe4_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe4_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe4_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe4_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe4_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe4_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe4_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe4_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe4_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe4_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe4_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe4_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe4_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe4_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe4_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe4_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe4_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe4_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe4_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe4_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe4_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe4_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe4_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe4_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe4_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe4_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe4_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe4_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe4_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe4_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe4_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe4_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe4_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe4_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe4_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe4_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe4_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe4_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe4_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe4_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe4_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe4_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe4_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe4_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe4_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe4_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe4_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe4_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe4_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe4_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe4_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe4_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe4_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe4_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe4_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe4_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe4_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe4_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe4_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe4_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe4_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe4_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe4_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe4_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe4_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe4_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe4_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe4_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe4_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe4_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe4_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe4_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe4_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe4_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe4_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe4_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe4_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe4_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe4_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe4_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe4_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe4_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe4_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe4_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe4_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe4_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe4_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe4_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe4_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe4_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe4_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe4_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe4_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe4_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe4_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe4_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe4_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe4_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe4_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe4_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe4_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe4_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe4_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe4_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe4_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe4_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe4_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe4_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe4_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe4_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe4_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe4_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe4_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe4_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe4_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe4_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe4_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe4_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe4_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe4_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe4_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe4_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe4_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe4_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe4_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe4_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe4_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe4_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe4_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe4_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe4_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe4_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe4_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe4_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe4_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe4_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe4_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe4_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe4_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe4_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe4_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe4_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe4_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe4_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe4_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe4_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe4_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe4_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe4_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe4_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe4_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe4_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe4_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe4_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe4_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe4_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe4_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe4_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe4_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe4_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe4_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe4_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe4_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe4_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe4_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe4_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe4_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe4_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe4_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe4_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe4_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe4_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe4_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe4_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe4_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe4_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe4_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe4_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe4_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe4_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe4_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe4_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe4_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe4_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe4_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe4_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe4_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe4_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe4_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe4_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe4_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe4_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe4_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe4_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe4_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe4_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe4_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe4_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe4_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe4_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe4_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe4_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe4_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe4_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(pipe4_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(pipe4_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(pipe4_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(pipe4_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(pipe4_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(pipe4_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(pipe4_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(pipe4_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(pipe4_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(pipe4_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(pipe4_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(pipe4_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(pipe4_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(pipe4_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(pipe4_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(pipe4_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(pipe4_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(pipe4_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(pipe4_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(pipe4_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(pipe4_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(pipe4_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(pipe4_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(pipe4_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(pipe4_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(pipe4_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(pipe4_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(pipe4_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(pipe4_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(pipe4_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(pipe4_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(pipe4_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(pipe4_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(pipe4_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(pipe4_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(pipe4_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(pipe4_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(pipe4_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(pipe4_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(pipe4_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(pipe4_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(pipe4_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(pipe4_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(pipe4_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(pipe4_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(pipe4_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(pipe4_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(pipe4_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(pipe4_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(pipe4_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(pipe4_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(pipe4_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(pipe4_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(pipe4_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(pipe4_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(pipe4_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(pipe4_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(pipe4_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(pipe4_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(pipe4_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(pipe4_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(pipe4_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(pipe4_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(pipe4_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(pipe4_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(pipe4_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(pipe4_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(pipe4_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(pipe4_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(pipe4_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(pipe4_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(pipe4_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(pipe4_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(pipe4_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(pipe4_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(pipe4_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(pipe4_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(pipe4_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(pipe4_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(pipe4_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(pipe4_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(pipe4_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(pipe4_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(pipe4_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(pipe4_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(pipe4_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(pipe4_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(pipe4_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(pipe4_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(pipe4_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(pipe4_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(pipe4_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(pipe4_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(pipe4_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(pipe4_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(pipe4_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(pipe4_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(pipe4_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(pipe4_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(pipe4_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(pipe4_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(pipe4_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(pipe4_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(pipe4_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(pipe4_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(pipe4_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(pipe4_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(pipe4_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(pipe4_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(pipe4_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(pipe4_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(pipe4_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(pipe4_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(pipe4_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(pipe4_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(pipe4_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(pipe4_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(pipe4_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(pipe4_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(pipe4_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(pipe4_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(pipe4_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(pipe4_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(pipe4_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(pipe4_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(pipe4_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(pipe4_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(pipe4_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(pipe4_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(pipe4_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(pipe4_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(pipe4_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(pipe4_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(pipe4_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(pipe4_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(pipe4_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(pipe4_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(pipe4_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(pipe4_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(pipe4_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(pipe4_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(pipe4_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(pipe4_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(pipe4_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(pipe4_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(pipe4_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(pipe4_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(pipe4_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(pipe4_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(pipe4_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(pipe4_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(pipe4_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(pipe4_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(pipe4_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(pipe4_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(pipe4_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(pipe4_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(pipe4_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(pipe4_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(pipe4_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(pipe4_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(pipe4_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(pipe4_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(pipe4_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(pipe4_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(pipe4_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(pipe4_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(pipe4_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(pipe4_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(pipe4_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(pipe4_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(pipe4_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(pipe4_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(pipe4_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(pipe4_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(pipe4_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(pipe4_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(pipe4_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(pipe4_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(pipe4_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(pipe4_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(pipe4_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(pipe4_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(pipe4_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(pipe4_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(pipe4_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(pipe4_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(pipe4_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(pipe4_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(pipe4_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(pipe4_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(pipe4_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(pipe4_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(pipe4_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(pipe4_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(pipe4_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(pipe4_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(pipe4_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(pipe4_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(pipe4_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(pipe4_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(pipe4_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(pipe4_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(pipe4_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(pipe4_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(pipe4_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(pipe4_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(pipe4_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(pipe4_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(pipe4_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(pipe4_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(pipe4_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(pipe4_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(pipe4_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(pipe4_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(pipe4_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(pipe4_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(pipe4_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(pipe4_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(pipe4_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(pipe4_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(pipe4_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(pipe4_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(pipe4_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(pipe4_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(pipe4_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(pipe4_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(pipe4_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(pipe4_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(pipe4_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(pipe4_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(pipe4_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(pipe4_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(pipe4_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(pipe4_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(pipe4_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(pipe4_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(pipe4_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(pipe4_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(pipe4_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(pipe4_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(pipe4_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(pipe4_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(pipe4_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(pipe4_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(pipe4_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(pipe4_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(pipe4_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(pipe4_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(pipe4_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(pipe4_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(pipe4_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(pipe4_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(pipe4_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(pipe4_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(pipe4_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_next_processor_id(pipe4_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe4_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe4_io_pipe_phv_out_is_valid_processor),
    .io_key_config_0_field_config_0(pipe4_io_key_config_0_field_config_0),
    .io_key_config_0_field_config_1(pipe4_io_key_config_0_field_config_1),
    .io_key_config_0_field_config_2(pipe4_io_key_config_0_field_config_2),
    .io_key_config_0_field_config_3(pipe4_io_key_config_0_field_config_3),
    .io_key_config_0_field_config_4(pipe4_io_key_config_0_field_config_4),
    .io_key_config_0_field_config_5(pipe4_io_key_config_0_field_config_5),
    .io_key_config_0_field_mask_0_0(pipe4_io_key_config_0_field_mask_0_0),
    .io_key_config_0_field_mask_0_1(pipe4_io_key_config_0_field_mask_0_1),
    .io_key_config_0_field_mask_0_2(pipe4_io_key_config_0_field_mask_0_2),
    .io_key_config_0_field_mask_0_3(pipe4_io_key_config_0_field_mask_0_3),
    .io_key_config_0_field_mask_1_0(pipe4_io_key_config_0_field_mask_1_0),
    .io_key_config_0_field_mask_1_1(pipe4_io_key_config_0_field_mask_1_1),
    .io_key_config_0_field_mask_1_2(pipe4_io_key_config_0_field_mask_1_2),
    .io_key_config_0_field_mask_1_3(pipe4_io_key_config_0_field_mask_1_3),
    .io_key_config_0_field_mask_2_0(pipe4_io_key_config_0_field_mask_2_0),
    .io_key_config_0_field_mask_2_1(pipe4_io_key_config_0_field_mask_2_1),
    .io_key_config_0_field_mask_2_2(pipe4_io_key_config_0_field_mask_2_2),
    .io_key_config_0_field_mask_2_3(pipe4_io_key_config_0_field_mask_2_3),
    .io_key_config_0_field_mask_3_0(pipe4_io_key_config_0_field_mask_3_0),
    .io_key_config_0_field_mask_3_1(pipe4_io_key_config_0_field_mask_3_1),
    .io_key_config_0_field_mask_3_2(pipe4_io_key_config_0_field_mask_3_2),
    .io_key_config_0_field_mask_3_3(pipe4_io_key_config_0_field_mask_3_3),
    .io_key_config_0_field_mask_4_0(pipe4_io_key_config_0_field_mask_4_0),
    .io_key_config_0_field_mask_4_1(pipe4_io_key_config_0_field_mask_4_1),
    .io_key_config_0_field_mask_4_2(pipe4_io_key_config_0_field_mask_4_2),
    .io_key_config_0_field_mask_4_3(pipe4_io_key_config_0_field_mask_4_3),
    .io_key_config_0_field_mask_5_0(pipe4_io_key_config_0_field_mask_5_0),
    .io_key_config_0_field_mask_5_1(pipe4_io_key_config_0_field_mask_5_1),
    .io_key_config_0_field_mask_5_2(pipe4_io_key_config_0_field_mask_5_2),
    .io_key_config_0_field_mask_5_3(pipe4_io_key_config_0_field_mask_5_3),
    .io_key_config_1_field_config_0(pipe4_io_key_config_1_field_config_0),
    .io_key_config_1_field_config_1(pipe4_io_key_config_1_field_config_1),
    .io_key_config_1_field_config_2(pipe4_io_key_config_1_field_config_2),
    .io_key_config_1_field_config_3(pipe4_io_key_config_1_field_config_3),
    .io_key_config_1_field_config_4(pipe4_io_key_config_1_field_config_4),
    .io_key_config_1_field_config_5(pipe4_io_key_config_1_field_config_5),
    .io_key_config_1_field_mask_0_0(pipe4_io_key_config_1_field_mask_0_0),
    .io_key_config_1_field_mask_0_1(pipe4_io_key_config_1_field_mask_0_1),
    .io_key_config_1_field_mask_0_2(pipe4_io_key_config_1_field_mask_0_2),
    .io_key_config_1_field_mask_0_3(pipe4_io_key_config_1_field_mask_0_3),
    .io_key_config_1_field_mask_1_0(pipe4_io_key_config_1_field_mask_1_0),
    .io_key_config_1_field_mask_1_1(pipe4_io_key_config_1_field_mask_1_1),
    .io_key_config_1_field_mask_1_2(pipe4_io_key_config_1_field_mask_1_2),
    .io_key_config_1_field_mask_1_3(pipe4_io_key_config_1_field_mask_1_3),
    .io_key_config_1_field_mask_2_0(pipe4_io_key_config_1_field_mask_2_0),
    .io_key_config_1_field_mask_2_1(pipe4_io_key_config_1_field_mask_2_1),
    .io_key_config_1_field_mask_2_2(pipe4_io_key_config_1_field_mask_2_2),
    .io_key_config_1_field_mask_2_3(pipe4_io_key_config_1_field_mask_2_3),
    .io_key_config_1_field_mask_3_0(pipe4_io_key_config_1_field_mask_3_0),
    .io_key_config_1_field_mask_3_1(pipe4_io_key_config_1_field_mask_3_1),
    .io_key_config_1_field_mask_3_2(pipe4_io_key_config_1_field_mask_3_2),
    .io_key_config_1_field_mask_3_3(pipe4_io_key_config_1_field_mask_3_3),
    .io_key_config_1_field_mask_4_0(pipe4_io_key_config_1_field_mask_4_0),
    .io_key_config_1_field_mask_4_1(pipe4_io_key_config_1_field_mask_4_1),
    .io_key_config_1_field_mask_4_2(pipe4_io_key_config_1_field_mask_4_2),
    .io_key_config_1_field_mask_4_3(pipe4_io_key_config_1_field_mask_4_3),
    .io_key_config_1_field_mask_5_0(pipe4_io_key_config_1_field_mask_5_0),
    .io_key_config_1_field_mask_5_1(pipe4_io_key_config_1_field_mask_5_1),
    .io_key_config_1_field_mask_5_2(pipe4_io_key_config_1_field_mask_5_2),
    .io_key_config_1_field_mask_5_3(pipe4_io_key_config_1_field_mask_5_3),
    .io_key_in(pipe4_io_key_in),
    .io_data_in(pipe4_io_data_in),
    .io_hit(pipe4_io_hit),
    .io_match_value(pipe4_io_match_value)
  );
  assign io_pipe_phv_out_data_0 = pipe4_io_pipe_phv_out_data_0; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_1 = pipe4_io_pipe_phv_out_data_1; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_2 = pipe4_io_pipe_phv_out_data_2; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_3 = pipe4_io_pipe_phv_out_data_3; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_4 = pipe4_io_pipe_phv_out_data_4; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_5 = pipe4_io_pipe_phv_out_data_5; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_6 = pipe4_io_pipe_phv_out_data_6; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_7 = pipe4_io_pipe_phv_out_data_7; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_8 = pipe4_io_pipe_phv_out_data_8; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_9 = pipe4_io_pipe_phv_out_data_9; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_10 = pipe4_io_pipe_phv_out_data_10; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_11 = pipe4_io_pipe_phv_out_data_11; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_12 = pipe4_io_pipe_phv_out_data_12; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_13 = pipe4_io_pipe_phv_out_data_13; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_14 = pipe4_io_pipe_phv_out_data_14; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_15 = pipe4_io_pipe_phv_out_data_15; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_16 = pipe4_io_pipe_phv_out_data_16; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_17 = pipe4_io_pipe_phv_out_data_17; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_18 = pipe4_io_pipe_phv_out_data_18; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_19 = pipe4_io_pipe_phv_out_data_19; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_20 = pipe4_io_pipe_phv_out_data_20; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_21 = pipe4_io_pipe_phv_out_data_21; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_22 = pipe4_io_pipe_phv_out_data_22; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_23 = pipe4_io_pipe_phv_out_data_23; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_24 = pipe4_io_pipe_phv_out_data_24; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_25 = pipe4_io_pipe_phv_out_data_25; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_26 = pipe4_io_pipe_phv_out_data_26; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_27 = pipe4_io_pipe_phv_out_data_27; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_28 = pipe4_io_pipe_phv_out_data_28; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_29 = pipe4_io_pipe_phv_out_data_29; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_30 = pipe4_io_pipe_phv_out_data_30; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_31 = pipe4_io_pipe_phv_out_data_31; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_32 = pipe4_io_pipe_phv_out_data_32; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_33 = pipe4_io_pipe_phv_out_data_33; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_34 = pipe4_io_pipe_phv_out_data_34; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_35 = pipe4_io_pipe_phv_out_data_35; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_36 = pipe4_io_pipe_phv_out_data_36; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_37 = pipe4_io_pipe_phv_out_data_37; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_38 = pipe4_io_pipe_phv_out_data_38; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_39 = pipe4_io_pipe_phv_out_data_39; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_40 = pipe4_io_pipe_phv_out_data_40; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_41 = pipe4_io_pipe_phv_out_data_41; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_42 = pipe4_io_pipe_phv_out_data_42; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_43 = pipe4_io_pipe_phv_out_data_43; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_44 = pipe4_io_pipe_phv_out_data_44; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_45 = pipe4_io_pipe_phv_out_data_45; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_46 = pipe4_io_pipe_phv_out_data_46; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_47 = pipe4_io_pipe_phv_out_data_47; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_48 = pipe4_io_pipe_phv_out_data_48; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_49 = pipe4_io_pipe_phv_out_data_49; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_50 = pipe4_io_pipe_phv_out_data_50; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_51 = pipe4_io_pipe_phv_out_data_51; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_52 = pipe4_io_pipe_phv_out_data_52; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_53 = pipe4_io_pipe_phv_out_data_53; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_54 = pipe4_io_pipe_phv_out_data_54; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_55 = pipe4_io_pipe_phv_out_data_55; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_56 = pipe4_io_pipe_phv_out_data_56; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_57 = pipe4_io_pipe_phv_out_data_57; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_58 = pipe4_io_pipe_phv_out_data_58; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_59 = pipe4_io_pipe_phv_out_data_59; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_60 = pipe4_io_pipe_phv_out_data_60; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_61 = pipe4_io_pipe_phv_out_data_61; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_62 = pipe4_io_pipe_phv_out_data_62; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_63 = pipe4_io_pipe_phv_out_data_63; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_64 = pipe4_io_pipe_phv_out_data_64; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_65 = pipe4_io_pipe_phv_out_data_65; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_66 = pipe4_io_pipe_phv_out_data_66; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_67 = pipe4_io_pipe_phv_out_data_67; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_68 = pipe4_io_pipe_phv_out_data_68; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_69 = pipe4_io_pipe_phv_out_data_69; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_70 = pipe4_io_pipe_phv_out_data_70; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_71 = pipe4_io_pipe_phv_out_data_71; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_72 = pipe4_io_pipe_phv_out_data_72; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_73 = pipe4_io_pipe_phv_out_data_73; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_74 = pipe4_io_pipe_phv_out_data_74; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_75 = pipe4_io_pipe_phv_out_data_75; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_76 = pipe4_io_pipe_phv_out_data_76; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_77 = pipe4_io_pipe_phv_out_data_77; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_78 = pipe4_io_pipe_phv_out_data_78; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_79 = pipe4_io_pipe_phv_out_data_79; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_80 = pipe4_io_pipe_phv_out_data_80; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_81 = pipe4_io_pipe_phv_out_data_81; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_82 = pipe4_io_pipe_phv_out_data_82; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_83 = pipe4_io_pipe_phv_out_data_83; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_84 = pipe4_io_pipe_phv_out_data_84; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_85 = pipe4_io_pipe_phv_out_data_85; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_86 = pipe4_io_pipe_phv_out_data_86; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_87 = pipe4_io_pipe_phv_out_data_87; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_88 = pipe4_io_pipe_phv_out_data_88; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_89 = pipe4_io_pipe_phv_out_data_89; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_90 = pipe4_io_pipe_phv_out_data_90; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_91 = pipe4_io_pipe_phv_out_data_91; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_92 = pipe4_io_pipe_phv_out_data_92; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_93 = pipe4_io_pipe_phv_out_data_93; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_94 = pipe4_io_pipe_phv_out_data_94; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_95 = pipe4_io_pipe_phv_out_data_95; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_96 = pipe4_io_pipe_phv_out_data_96; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_97 = pipe4_io_pipe_phv_out_data_97; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_98 = pipe4_io_pipe_phv_out_data_98; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_99 = pipe4_io_pipe_phv_out_data_99; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_100 = pipe4_io_pipe_phv_out_data_100; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_101 = pipe4_io_pipe_phv_out_data_101; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_102 = pipe4_io_pipe_phv_out_data_102; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_103 = pipe4_io_pipe_phv_out_data_103; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_104 = pipe4_io_pipe_phv_out_data_104; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_105 = pipe4_io_pipe_phv_out_data_105; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_106 = pipe4_io_pipe_phv_out_data_106; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_107 = pipe4_io_pipe_phv_out_data_107; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_108 = pipe4_io_pipe_phv_out_data_108; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_109 = pipe4_io_pipe_phv_out_data_109; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_110 = pipe4_io_pipe_phv_out_data_110; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_111 = pipe4_io_pipe_phv_out_data_111; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_112 = pipe4_io_pipe_phv_out_data_112; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_113 = pipe4_io_pipe_phv_out_data_113; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_114 = pipe4_io_pipe_phv_out_data_114; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_115 = pipe4_io_pipe_phv_out_data_115; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_116 = pipe4_io_pipe_phv_out_data_116; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_117 = pipe4_io_pipe_phv_out_data_117; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_118 = pipe4_io_pipe_phv_out_data_118; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_119 = pipe4_io_pipe_phv_out_data_119; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_120 = pipe4_io_pipe_phv_out_data_120; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_121 = pipe4_io_pipe_phv_out_data_121; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_122 = pipe4_io_pipe_phv_out_data_122; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_123 = pipe4_io_pipe_phv_out_data_123; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_124 = pipe4_io_pipe_phv_out_data_124; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_125 = pipe4_io_pipe_phv_out_data_125; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_126 = pipe4_io_pipe_phv_out_data_126; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_127 = pipe4_io_pipe_phv_out_data_127; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_128 = pipe4_io_pipe_phv_out_data_128; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_129 = pipe4_io_pipe_phv_out_data_129; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_130 = pipe4_io_pipe_phv_out_data_130; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_131 = pipe4_io_pipe_phv_out_data_131; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_132 = pipe4_io_pipe_phv_out_data_132; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_133 = pipe4_io_pipe_phv_out_data_133; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_134 = pipe4_io_pipe_phv_out_data_134; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_135 = pipe4_io_pipe_phv_out_data_135; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_136 = pipe4_io_pipe_phv_out_data_136; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_137 = pipe4_io_pipe_phv_out_data_137; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_138 = pipe4_io_pipe_phv_out_data_138; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_139 = pipe4_io_pipe_phv_out_data_139; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_140 = pipe4_io_pipe_phv_out_data_140; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_141 = pipe4_io_pipe_phv_out_data_141; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_142 = pipe4_io_pipe_phv_out_data_142; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_143 = pipe4_io_pipe_phv_out_data_143; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_144 = pipe4_io_pipe_phv_out_data_144; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_145 = pipe4_io_pipe_phv_out_data_145; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_146 = pipe4_io_pipe_phv_out_data_146; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_147 = pipe4_io_pipe_phv_out_data_147; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_148 = pipe4_io_pipe_phv_out_data_148; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_149 = pipe4_io_pipe_phv_out_data_149; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_150 = pipe4_io_pipe_phv_out_data_150; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_151 = pipe4_io_pipe_phv_out_data_151; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_152 = pipe4_io_pipe_phv_out_data_152; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_153 = pipe4_io_pipe_phv_out_data_153; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_154 = pipe4_io_pipe_phv_out_data_154; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_155 = pipe4_io_pipe_phv_out_data_155; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_156 = pipe4_io_pipe_phv_out_data_156; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_157 = pipe4_io_pipe_phv_out_data_157; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_158 = pipe4_io_pipe_phv_out_data_158; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_159 = pipe4_io_pipe_phv_out_data_159; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_160 = pipe4_io_pipe_phv_out_data_160; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_161 = pipe4_io_pipe_phv_out_data_161; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_162 = pipe4_io_pipe_phv_out_data_162; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_163 = pipe4_io_pipe_phv_out_data_163; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_164 = pipe4_io_pipe_phv_out_data_164; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_165 = pipe4_io_pipe_phv_out_data_165; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_166 = pipe4_io_pipe_phv_out_data_166; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_167 = pipe4_io_pipe_phv_out_data_167; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_168 = pipe4_io_pipe_phv_out_data_168; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_169 = pipe4_io_pipe_phv_out_data_169; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_170 = pipe4_io_pipe_phv_out_data_170; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_171 = pipe4_io_pipe_phv_out_data_171; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_172 = pipe4_io_pipe_phv_out_data_172; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_173 = pipe4_io_pipe_phv_out_data_173; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_174 = pipe4_io_pipe_phv_out_data_174; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_175 = pipe4_io_pipe_phv_out_data_175; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_176 = pipe4_io_pipe_phv_out_data_176; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_177 = pipe4_io_pipe_phv_out_data_177; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_178 = pipe4_io_pipe_phv_out_data_178; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_179 = pipe4_io_pipe_phv_out_data_179; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_180 = pipe4_io_pipe_phv_out_data_180; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_181 = pipe4_io_pipe_phv_out_data_181; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_182 = pipe4_io_pipe_phv_out_data_182; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_183 = pipe4_io_pipe_phv_out_data_183; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_184 = pipe4_io_pipe_phv_out_data_184; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_185 = pipe4_io_pipe_phv_out_data_185; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_186 = pipe4_io_pipe_phv_out_data_186; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_187 = pipe4_io_pipe_phv_out_data_187; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_188 = pipe4_io_pipe_phv_out_data_188; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_189 = pipe4_io_pipe_phv_out_data_189; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_190 = pipe4_io_pipe_phv_out_data_190; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_191 = pipe4_io_pipe_phv_out_data_191; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_192 = pipe4_io_pipe_phv_out_data_192; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_193 = pipe4_io_pipe_phv_out_data_193; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_194 = pipe4_io_pipe_phv_out_data_194; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_195 = pipe4_io_pipe_phv_out_data_195; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_196 = pipe4_io_pipe_phv_out_data_196; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_197 = pipe4_io_pipe_phv_out_data_197; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_198 = pipe4_io_pipe_phv_out_data_198; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_199 = pipe4_io_pipe_phv_out_data_199; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_200 = pipe4_io_pipe_phv_out_data_200; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_201 = pipe4_io_pipe_phv_out_data_201; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_202 = pipe4_io_pipe_phv_out_data_202; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_203 = pipe4_io_pipe_phv_out_data_203; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_204 = pipe4_io_pipe_phv_out_data_204; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_205 = pipe4_io_pipe_phv_out_data_205; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_206 = pipe4_io_pipe_phv_out_data_206; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_207 = pipe4_io_pipe_phv_out_data_207; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_208 = pipe4_io_pipe_phv_out_data_208; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_209 = pipe4_io_pipe_phv_out_data_209; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_210 = pipe4_io_pipe_phv_out_data_210; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_211 = pipe4_io_pipe_phv_out_data_211; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_212 = pipe4_io_pipe_phv_out_data_212; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_213 = pipe4_io_pipe_phv_out_data_213; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_214 = pipe4_io_pipe_phv_out_data_214; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_215 = pipe4_io_pipe_phv_out_data_215; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_216 = pipe4_io_pipe_phv_out_data_216; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_217 = pipe4_io_pipe_phv_out_data_217; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_218 = pipe4_io_pipe_phv_out_data_218; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_219 = pipe4_io_pipe_phv_out_data_219; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_220 = pipe4_io_pipe_phv_out_data_220; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_221 = pipe4_io_pipe_phv_out_data_221; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_222 = pipe4_io_pipe_phv_out_data_222; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_223 = pipe4_io_pipe_phv_out_data_223; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_224 = pipe4_io_pipe_phv_out_data_224; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_225 = pipe4_io_pipe_phv_out_data_225; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_226 = pipe4_io_pipe_phv_out_data_226; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_227 = pipe4_io_pipe_phv_out_data_227; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_228 = pipe4_io_pipe_phv_out_data_228; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_229 = pipe4_io_pipe_phv_out_data_229; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_230 = pipe4_io_pipe_phv_out_data_230; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_231 = pipe4_io_pipe_phv_out_data_231; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_232 = pipe4_io_pipe_phv_out_data_232; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_233 = pipe4_io_pipe_phv_out_data_233; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_234 = pipe4_io_pipe_phv_out_data_234; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_235 = pipe4_io_pipe_phv_out_data_235; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_236 = pipe4_io_pipe_phv_out_data_236; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_237 = pipe4_io_pipe_phv_out_data_237; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_238 = pipe4_io_pipe_phv_out_data_238; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_239 = pipe4_io_pipe_phv_out_data_239; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_240 = pipe4_io_pipe_phv_out_data_240; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_241 = pipe4_io_pipe_phv_out_data_241; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_242 = pipe4_io_pipe_phv_out_data_242; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_243 = pipe4_io_pipe_phv_out_data_243; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_244 = pipe4_io_pipe_phv_out_data_244; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_245 = pipe4_io_pipe_phv_out_data_245; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_246 = pipe4_io_pipe_phv_out_data_246; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_247 = pipe4_io_pipe_phv_out_data_247; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_248 = pipe4_io_pipe_phv_out_data_248; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_249 = pipe4_io_pipe_phv_out_data_249; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_250 = pipe4_io_pipe_phv_out_data_250; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_251 = pipe4_io_pipe_phv_out_data_251; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_252 = pipe4_io_pipe_phv_out_data_252; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_253 = pipe4_io_pipe_phv_out_data_253; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_254 = pipe4_io_pipe_phv_out_data_254; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_255 = pipe4_io_pipe_phv_out_data_255; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_256 = pipe4_io_pipe_phv_out_data_256; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_257 = pipe4_io_pipe_phv_out_data_257; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_258 = pipe4_io_pipe_phv_out_data_258; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_259 = pipe4_io_pipe_phv_out_data_259; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_260 = pipe4_io_pipe_phv_out_data_260; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_261 = pipe4_io_pipe_phv_out_data_261; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_262 = pipe4_io_pipe_phv_out_data_262; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_263 = pipe4_io_pipe_phv_out_data_263; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_264 = pipe4_io_pipe_phv_out_data_264; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_265 = pipe4_io_pipe_phv_out_data_265; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_266 = pipe4_io_pipe_phv_out_data_266; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_267 = pipe4_io_pipe_phv_out_data_267; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_268 = pipe4_io_pipe_phv_out_data_268; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_269 = pipe4_io_pipe_phv_out_data_269; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_270 = pipe4_io_pipe_phv_out_data_270; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_271 = pipe4_io_pipe_phv_out_data_271; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_272 = pipe4_io_pipe_phv_out_data_272; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_273 = pipe4_io_pipe_phv_out_data_273; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_274 = pipe4_io_pipe_phv_out_data_274; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_275 = pipe4_io_pipe_phv_out_data_275; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_276 = pipe4_io_pipe_phv_out_data_276; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_277 = pipe4_io_pipe_phv_out_data_277; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_278 = pipe4_io_pipe_phv_out_data_278; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_279 = pipe4_io_pipe_phv_out_data_279; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_280 = pipe4_io_pipe_phv_out_data_280; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_281 = pipe4_io_pipe_phv_out_data_281; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_282 = pipe4_io_pipe_phv_out_data_282; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_283 = pipe4_io_pipe_phv_out_data_283; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_284 = pipe4_io_pipe_phv_out_data_284; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_285 = pipe4_io_pipe_phv_out_data_285; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_286 = pipe4_io_pipe_phv_out_data_286; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_287 = pipe4_io_pipe_phv_out_data_287; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_288 = pipe4_io_pipe_phv_out_data_288; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_289 = pipe4_io_pipe_phv_out_data_289; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_290 = pipe4_io_pipe_phv_out_data_290; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_291 = pipe4_io_pipe_phv_out_data_291; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_292 = pipe4_io_pipe_phv_out_data_292; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_293 = pipe4_io_pipe_phv_out_data_293; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_294 = pipe4_io_pipe_phv_out_data_294; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_295 = pipe4_io_pipe_phv_out_data_295; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_296 = pipe4_io_pipe_phv_out_data_296; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_297 = pipe4_io_pipe_phv_out_data_297; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_298 = pipe4_io_pipe_phv_out_data_298; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_299 = pipe4_io_pipe_phv_out_data_299; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_300 = pipe4_io_pipe_phv_out_data_300; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_301 = pipe4_io_pipe_phv_out_data_301; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_302 = pipe4_io_pipe_phv_out_data_302; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_303 = pipe4_io_pipe_phv_out_data_303; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_304 = pipe4_io_pipe_phv_out_data_304; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_305 = pipe4_io_pipe_phv_out_data_305; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_306 = pipe4_io_pipe_phv_out_data_306; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_307 = pipe4_io_pipe_phv_out_data_307; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_308 = pipe4_io_pipe_phv_out_data_308; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_309 = pipe4_io_pipe_phv_out_data_309; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_310 = pipe4_io_pipe_phv_out_data_310; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_311 = pipe4_io_pipe_phv_out_data_311; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_312 = pipe4_io_pipe_phv_out_data_312; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_313 = pipe4_io_pipe_phv_out_data_313; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_314 = pipe4_io_pipe_phv_out_data_314; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_315 = pipe4_io_pipe_phv_out_data_315; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_316 = pipe4_io_pipe_phv_out_data_316; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_317 = pipe4_io_pipe_phv_out_data_317; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_318 = pipe4_io_pipe_phv_out_data_318; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_319 = pipe4_io_pipe_phv_out_data_319; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_320 = pipe4_io_pipe_phv_out_data_320; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_321 = pipe4_io_pipe_phv_out_data_321; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_322 = pipe4_io_pipe_phv_out_data_322; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_323 = pipe4_io_pipe_phv_out_data_323; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_324 = pipe4_io_pipe_phv_out_data_324; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_325 = pipe4_io_pipe_phv_out_data_325; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_326 = pipe4_io_pipe_phv_out_data_326; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_327 = pipe4_io_pipe_phv_out_data_327; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_328 = pipe4_io_pipe_phv_out_data_328; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_329 = pipe4_io_pipe_phv_out_data_329; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_330 = pipe4_io_pipe_phv_out_data_330; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_331 = pipe4_io_pipe_phv_out_data_331; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_332 = pipe4_io_pipe_phv_out_data_332; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_333 = pipe4_io_pipe_phv_out_data_333; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_334 = pipe4_io_pipe_phv_out_data_334; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_335 = pipe4_io_pipe_phv_out_data_335; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_336 = pipe4_io_pipe_phv_out_data_336; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_337 = pipe4_io_pipe_phv_out_data_337; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_338 = pipe4_io_pipe_phv_out_data_338; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_339 = pipe4_io_pipe_phv_out_data_339; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_340 = pipe4_io_pipe_phv_out_data_340; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_341 = pipe4_io_pipe_phv_out_data_341; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_342 = pipe4_io_pipe_phv_out_data_342; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_343 = pipe4_io_pipe_phv_out_data_343; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_344 = pipe4_io_pipe_phv_out_data_344; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_345 = pipe4_io_pipe_phv_out_data_345; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_346 = pipe4_io_pipe_phv_out_data_346; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_347 = pipe4_io_pipe_phv_out_data_347; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_348 = pipe4_io_pipe_phv_out_data_348; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_349 = pipe4_io_pipe_phv_out_data_349; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_350 = pipe4_io_pipe_phv_out_data_350; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_351 = pipe4_io_pipe_phv_out_data_351; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_352 = pipe4_io_pipe_phv_out_data_352; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_353 = pipe4_io_pipe_phv_out_data_353; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_354 = pipe4_io_pipe_phv_out_data_354; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_355 = pipe4_io_pipe_phv_out_data_355; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_356 = pipe4_io_pipe_phv_out_data_356; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_357 = pipe4_io_pipe_phv_out_data_357; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_358 = pipe4_io_pipe_phv_out_data_358; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_359 = pipe4_io_pipe_phv_out_data_359; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_360 = pipe4_io_pipe_phv_out_data_360; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_361 = pipe4_io_pipe_phv_out_data_361; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_362 = pipe4_io_pipe_phv_out_data_362; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_363 = pipe4_io_pipe_phv_out_data_363; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_364 = pipe4_io_pipe_phv_out_data_364; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_365 = pipe4_io_pipe_phv_out_data_365; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_366 = pipe4_io_pipe_phv_out_data_366; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_367 = pipe4_io_pipe_phv_out_data_367; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_368 = pipe4_io_pipe_phv_out_data_368; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_369 = pipe4_io_pipe_phv_out_data_369; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_370 = pipe4_io_pipe_phv_out_data_370; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_371 = pipe4_io_pipe_phv_out_data_371; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_372 = pipe4_io_pipe_phv_out_data_372; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_373 = pipe4_io_pipe_phv_out_data_373; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_374 = pipe4_io_pipe_phv_out_data_374; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_375 = pipe4_io_pipe_phv_out_data_375; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_376 = pipe4_io_pipe_phv_out_data_376; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_377 = pipe4_io_pipe_phv_out_data_377; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_378 = pipe4_io_pipe_phv_out_data_378; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_379 = pipe4_io_pipe_phv_out_data_379; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_380 = pipe4_io_pipe_phv_out_data_380; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_381 = pipe4_io_pipe_phv_out_data_381; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_382 = pipe4_io_pipe_phv_out_data_382; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_383 = pipe4_io_pipe_phv_out_data_383; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_384 = pipe4_io_pipe_phv_out_data_384; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_385 = pipe4_io_pipe_phv_out_data_385; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_386 = pipe4_io_pipe_phv_out_data_386; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_387 = pipe4_io_pipe_phv_out_data_387; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_388 = pipe4_io_pipe_phv_out_data_388; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_389 = pipe4_io_pipe_phv_out_data_389; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_390 = pipe4_io_pipe_phv_out_data_390; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_391 = pipe4_io_pipe_phv_out_data_391; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_392 = pipe4_io_pipe_phv_out_data_392; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_393 = pipe4_io_pipe_phv_out_data_393; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_394 = pipe4_io_pipe_phv_out_data_394; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_395 = pipe4_io_pipe_phv_out_data_395; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_396 = pipe4_io_pipe_phv_out_data_396; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_397 = pipe4_io_pipe_phv_out_data_397; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_398 = pipe4_io_pipe_phv_out_data_398; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_399 = pipe4_io_pipe_phv_out_data_399; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_400 = pipe4_io_pipe_phv_out_data_400; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_401 = pipe4_io_pipe_phv_out_data_401; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_402 = pipe4_io_pipe_phv_out_data_402; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_403 = pipe4_io_pipe_phv_out_data_403; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_404 = pipe4_io_pipe_phv_out_data_404; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_405 = pipe4_io_pipe_phv_out_data_405; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_406 = pipe4_io_pipe_phv_out_data_406; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_407 = pipe4_io_pipe_phv_out_data_407; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_408 = pipe4_io_pipe_phv_out_data_408; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_409 = pipe4_io_pipe_phv_out_data_409; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_410 = pipe4_io_pipe_phv_out_data_410; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_411 = pipe4_io_pipe_phv_out_data_411; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_412 = pipe4_io_pipe_phv_out_data_412; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_413 = pipe4_io_pipe_phv_out_data_413; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_414 = pipe4_io_pipe_phv_out_data_414; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_415 = pipe4_io_pipe_phv_out_data_415; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_416 = pipe4_io_pipe_phv_out_data_416; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_417 = pipe4_io_pipe_phv_out_data_417; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_418 = pipe4_io_pipe_phv_out_data_418; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_419 = pipe4_io_pipe_phv_out_data_419; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_420 = pipe4_io_pipe_phv_out_data_420; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_421 = pipe4_io_pipe_phv_out_data_421; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_422 = pipe4_io_pipe_phv_out_data_422; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_423 = pipe4_io_pipe_phv_out_data_423; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_424 = pipe4_io_pipe_phv_out_data_424; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_425 = pipe4_io_pipe_phv_out_data_425; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_426 = pipe4_io_pipe_phv_out_data_426; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_427 = pipe4_io_pipe_phv_out_data_427; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_428 = pipe4_io_pipe_phv_out_data_428; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_429 = pipe4_io_pipe_phv_out_data_429; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_430 = pipe4_io_pipe_phv_out_data_430; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_431 = pipe4_io_pipe_phv_out_data_431; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_432 = pipe4_io_pipe_phv_out_data_432; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_433 = pipe4_io_pipe_phv_out_data_433; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_434 = pipe4_io_pipe_phv_out_data_434; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_435 = pipe4_io_pipe_phv_out_data_435; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_436 = pipe4_io_pipe_phv_out_data_436; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_437 = pipe4_io_pipe_phv_out_data_437; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_438 = pipe4_io_pipe_phv_out_data_438; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_439 = pipe4_io_pipe_phv_out_data_439; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_440 = pipe4_io_pipe_phv_out_data_440; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_441 = pipe4_io_pipe_phv_out_data_441; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_442 = pipe4_io_pipe_phv_out_data_442; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_443 = pipe4_io_pipe_phv_out_data_443; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_444 = pipe4_io_pipe_phv_out_data_444; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_445 = pipe4_io_pipe_phv_out_data_445; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_446 = pipe4_io_pipe_phv_out_data_446; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_447 = pipe4_io_pipe_phv_out_data_447; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_448 = pipe4_io_pipe_phv_out_data_448; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_449 = pipe4_io_pipe_phv_out_data_449; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_450 = pipe4_io_pipe_phv_out_data_450; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_451 = pipe4_io_pipe_phv_out_data_451; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_452 = pipe4_io_pipe_phv_out_data_452; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_453 = pipe4_io_pipe_phv_out_data_453; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_454 = pipe4_io_pipe_phv_out_data_454; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_455 = pipe4_io_pipe_phv_out_data_455; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_456 = pipe4_io_pipe_phv_out_data_456; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_457 = pipe4_io_pipe_phv_out_data_457; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_458 = pipe4_io_pipe_phv_out_data_458; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_459 = pipe4_io_pipe_phv_out_data_459; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_460 = pipe4_io_pipe_phv_out_data_460; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_461 = pipe4_io_pipe_phv_out_data_461; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_462 = pipe4_io_pipe_phv_out_data_462; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_463 = pipe4_io_pipe_phv_out_data_463; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_464 = pipe4_io_pipe_phv_out_data_464; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_465 = pipe4_io_pipe_phv_out_data_465; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_466 = pipe4_io_pipe_phv_out_data_466; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_467 = pipe4_io_pipe_phv_out_data_467; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_468 = pipe4_io_pipe_phv_out_data_468; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_469 = pipe4_io_pipe_phv_out_data_469; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_470 = pipe4_io_pipe_phv_out_data_470; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_471 = pipe4_io_pipe_phv_out_data_471; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_472 = pipe4_io_pipe_phv_out_data_472; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_473 = pipe4_io_pipe_phv_out_data_473; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_474 = pipe4_io_pipe_phv_out_data_474; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_475 = pipe4_io_pipe_phv_out_data_475; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_476 = pipe4_io_pipe_phv_out_data_476; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_477 = pipe4_io_pipe_phv_out_data_477; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_478 = pipe4_io_pipe_phv_out_data_478; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_479 = pipe4_io_pipe_phv_out_data_479; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_480 = pipe4_io_pipe_phv_out_data_480; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_481 = pipe4_io_pipe_phv_out_data_481; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_482 = pipe4_io_pipe_phv_out_data_482; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_483 = pipe4_io_pipe_phv_out_data_483; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_484 = pipe4_io_pipe_phv_out_data_484; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_485 = pipe4_io_pipe_phv_out_data_485; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_486 = pipe4_io_pipe_phv_out_data_486; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_487 = pipe4_io_pipe_phv_out_data_487; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_488 = pipe4_io_pipe_phv_out_data_488; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_489 = pipe4_io_pipe_phv_out_data_489; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_490 = pipe4_io_pipe_phv_out_data_490; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_491 = pipe4_io_pipe_phv_out_data_491; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_492 = pipe4_io_pipe_phv_out_data_492; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_493 = pipe4_io_pipe_phv_out_data_493; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_494 = pipe4_io_pipe_phv_out_data_494; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_495 = pipe4_io_pipe_phv_out_data_495; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_496 = pipe4_io_pipe_phv_out_data_496; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_497 = pipe4_io_pipe_phv_out_data_497; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_498 = pipe4_io_pipe_phv_out_data_498; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_499 = pipe4_io_pipe_phv_out_data_499; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_500 = pipe4_io_pipe_phv_out_data_500; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_501 = pipe4_io_pipe_phv_out_data_501; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_502 = pipe4_io_pipe_phv_out_data_502; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_503 = pipe4_io_pipe_phv_out_data_503; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_504 = pipe4_io_pipe_phv_out_data_504; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_505 = pipe4_io_pipe_phv_out_data_505; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_506 = pipe4_io_pipe_phv_out_data_506; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_507 = pipe4_io_pipe_phv_out_data_507; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_508 = pipe4_io_pipe_phv_out_data_508; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_509 = pipe4_io_pipe_phv_out_data_509; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_510 = pipe4_io_pipe_phv_out_data_510; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_data_511 = pipe4_io_pipe_phv_out_data_511; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_next_processor_id = pipe4_io_pipe_phv_out_next_processor_id; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_next_config_id = pipe4_io_pipe_phv_out_next_config_id; // @[matcher_pisa.scala 359:26]
  assign io_pipe_phv_out_is_valid_processor = pipe4_io_pipe_phv_out_is_valid_processor; // @[matcher_pisa.scala 359:26]
  assign io_hit = pipe4_io_hit; // @[matcher_pisa.scala 360:26]
  assign io_match_value = pipe4_io_match_value; // @[matcher_pisa.scala 361:26]
  assign pipe1_clock = clock;
  assign pipe1_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_96 = io_pipe_phv_in_data_96; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_97 = io_pipe_phv_in_data_97; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_98 = io_pipe_phv_in_data_98; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_99 = io_pipe_phv_in_data_99; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_100 = io_pipe_phv_in_data_100; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_101 = io_pipe_phv_in_data_101; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_102 = io_pipe_phv_in_data_102; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_103 = io_pipe_phv_in_data_103; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_104 = io_pipe_phv_in_data_104; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_105 = io_pipe_phv_in_data_105; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_106 = io_pipe_phv_in_data_106; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_107 = io_pipe_phv_in_data_107; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_108 = io_pipe_phv_in_data_108; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_109 = io_pipe_phv_in_data_109; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_110 = io_pipe_phv_in_data_110; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_111 = io_pipe_phv_in_data_111; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_112 = io_pipe_phv_in_data_112; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_113 = io_pipe_phv_in_data_113; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_114 = io_pipe_phv_in_data_114; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_115 = io_pipe_phv_in_data_115; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_116 = io_pipe_phv_in_data_116; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_117 = io_pipe_phv_in_data_117; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_118 = io_pipe_phv_in_data_118; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_119 = io_pipe_phv_in_data_119; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_120 = io_pipe_phv_in_data_120; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_121 = io_pipe_phv_in_data_121; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_122 = io_pipe_phv_in_data_122; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_123 = io_pipe_phv_in_data_123; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_124 = io_pipe_phv_in_data_124; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_125 = io_pipe_phv_in_data_125; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_126 = io_pipe_phv_in_data_126; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_127 = io_pipe_phv_in_data_127; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_128 = io_pipe_phv_in_data_128; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_129 = io_pipe_phv_in_data_129; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_130 = io_pipe_phv_in_data_130; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_131 = io_pipe_phv_in_data_131; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_132 = io_pipe_phv_in_data_132; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_133 = io_pipe_phv_in_data_133; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_134 = io_pipe_phv_in_data_134; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_135 = io_pipe_phv_in_data_135; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_136 = io_pipe_phv_in_data_136; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_137 = io_pipe_phv_in_data_137; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_138 = io_pipe_phv_in_data_138; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_139 = io_pipe_phv_in_data_139; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_140 = io_pipe_phv_in_data_140; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_141 = io_pipe_phv_in_data_141; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_142 = io_pipe_phv_in_data_142; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_143 = io_pipe_phv_in_data_143; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_144 = io_pipe_phv_in_data_144; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_145 = io_pipe_phv_in_data_145; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_146 = io_pipe_phv_in_data_146; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_147 = io_pipe_phv_in_data_147; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_148 = io_pipe_phv_in_data_148; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_149 = io_pipe_phv_in_data_149; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_150 = io_pipe_phv_in_data_150; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_151 = io_pipe_phv_in_data_151; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_152 = io_pipe_phv_in_data_152; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_153 = io_pipe_phv_in_data_153; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_154 = io_pipe_phv_in_data_154; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_155 = io_pipe_phv_in_data_155; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_156 = io_pipe_phv_in_data_156; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_157 = io_pipe_phv_in_data_157; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_158 = io_pipe_phv_in_data_158; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_159 = io_pipe_phv_in_data_159; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_160 = io_pipe_phv_in_data_160; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_161 = io_pipe_phv_in_data_161; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_162 = io_pipe_phv_in_data_162; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_163 = io_pipe_phv_in_data_163; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_164 = io_pipe_phv_in_data_164; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_165 = io_pipe_phv_in_data_165; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_166 = io_pipe_phv_in_data_166; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_167 = io_pipe_phv_in_data_167; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_168 = io_pipe_phv_in_data_168; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_169 = io_pipe_phv_in_data_169; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_170 = io_pipe_phv_in_data_170; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_171 = io_pipe_phv_in_data_171; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_172 = io_pipe_phv_in_data_172; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_173 = io_pipe_phv_in_data_173; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_174 = io_pipe_phv_in_data_174; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_175 = io_pipe_phv_in_data_175; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_176 = io_pipe_phv_in_data_176; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_177 = io_pipe_phv_in_data_177; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_178 = io_pipe_phv_in_data_178; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_179 = io_pipe_phv_in_data_179; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_180 = io_pipe_phv_in_data_180; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_181 = io_pipe_phv_in_data_181; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_182 = io_pipe_phv_in_data_182; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_183 = io_pipe_phv_in_data_183; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_184 = io_pipe_phv_in_data_184; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_185 = io_pipe_phv_in_data_185; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_186 = io_pipe_phv_in_data_186; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_187 = io_pipe_phv_in_data_187; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_188 = io_pipe_phv_in_data_188; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_189 = io_pipe_phv_in_data_189; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_190 = io_pipe_phv_in_data_190; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_191 = io_pipe_phv_in_data_191; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_192 = io_pipe_phv_in_data_192; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_193 = io_pipe_phv_in_data_193; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_194 = io_pipe_phv_in_data_194; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_195 = io_pipe_phv_in_data_195; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_196 = io_pipe_phv_in_data_196; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_197 = io_pipe_phv_in_data_197; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_198 = io_pipe_phv_in_data_198; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_199 = io_pipe_phv_in_data_199; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_200 = io_pipe_phv_in_data_200; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_201 = io_pipe_phv_in_data_201; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_202 = io_pipe_phv_in_data_202; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_203 = io_pipe_phv_in_data_203; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_204 = io_pipe_phv_in_data_204; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_205 = io_pipe_phv_in_data_205; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_206 = io_pipe_phv_in_data_206; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_207 = io_pipe_phv_in_data_207; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_208 = io_pipe_phv_in_data_208; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_209 = io_pipe_phv_in_data_209; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_210 = io_pipe_phv_in_data_210; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_211 = io_pipe_phv_in_data_211; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_212 = io_pipe_phv_in_data_212; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_213 = io_pipe_phv_in_data_213; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_214 = io_pipe_phv_in_data_214; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_215 = io_pipe_phv_in_data_215; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_216 = io_pipe_phv_in_data_216; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_217 = io_pipe_phv_in_data_217; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_218 = io_pipe_phv_in_data_218; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_219 = io_pipe_phv_in_data_219; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_220 = io_pipe_phv_in_data_220; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_221 = io_pipe_phv_in_data_221; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_222 = io_pipe_phv_in_data_222; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_223 = io_pipe_phv_in_data_223; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_224 = io_pipe_phv_in_data_224; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_225 = io_pipe_phv_in_data_225; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_226 = io_pipe_phv_in_data_226; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_227 = io_pipe_phv_in_data_227; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_228 = io_pipe_phv_in_data_228; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_229 = io_pipe_phv_in_data_229; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_230 = io_pipe_phv_in_data_230; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_231 = io_pipe_phv_in_data_231; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_232 = io_pipe_phv_in_data_232; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_233 = io_pipe_phv_in_data_233; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_234 = io_pipe_phv_in_data_234; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_235 = io_pipe_phv_in_data_235; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_236 = io_pipe_phv_in_data_236; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_237 = io_pipe_phv_in_data_237; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_238 = io_pipe_phv_in_data_238; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_239 = io_pipe_phv_in_data_239; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_240 = io_pipe_phv_in_data_240; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_241 = io_pipe_phv_in_data_241; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_242 = io_pipe_phv_in_data_242; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_243 = io_pipe_phv_in_data_243; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_244 = io_pipe_phv_in_data_244; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_245 = io_pipe_phv_in_data_245; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_246 = io_pipe_phv_in_data_246; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_247 = io_pipe_phv_in_data_247; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_248 = io_pipe_phv_in_data_248; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_249 = io_pipe_phv_in_data_249; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_250 = io_pipe_phv_in_data_250; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_251 = io_pipe_phv_in_data_251; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_252 = io_pipe_phv_in_data_252; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_253 = io_pipe_phv_in_data_253; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_254 = io_pipe_phv_in_data_254; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_255 = io_pipe_phv_in_data_255; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_256 = io_pipe_phv_in_data_256; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_257 = io_pipe_phv_in_data_257; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_258 = io_pipe_phv_in_data_258; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_259 = io_pipe_phv_in_data_259; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_260 = io_pipe_phv_in_data_260; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_261 = io_pipe_phv_in_data_261; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_262 = io_pipe_phv_in_data_262; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_263 = io_pipe_phv_in_data_263; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_264 = io_pipe_phv_in_data_264; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_265 = io_pipe_phv_in_data_265; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_266 = io_pipe_phv_in_data_266; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_267 = io_pipe_phv_in_data_267; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_268 = io_pipe_phv_in_data_268; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_269 = io_pipe_phv_in_data_269; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_270 = io_pipe_phv_in_data_270; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_271 = io_pipe_phv_in_data_271; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_272 = io_pipe_phv_in_data_272; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_273 = io_pipe_phv_in_data_273; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_274 = io_pipe_phv_in_data_274; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_275 = io_pipe_phv_in_data_275; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_276 = io_pipe_phv_in_data_276; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_277 = io_pipe_phv_in_data_277; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_278 = io_pipe_phv_in_data_278; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_279 = io_pipe_phv_in_data_279; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_280 = io_pipe_phv_in_data_280; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_281 = io_pipe_phv_in_data_281; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_282 = io_pipe_phv_in_data_282; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_283 = io_pipe_phv_in_data_283; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_284 = io_pipe_phv_in_data_284; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_285 = io_pipe_phv_in_data_285; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_286 = io_pipe_phv_in_data_286; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_287 = io_pipe_phv_in_data_287; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_288 = io_pipe_phv_in_data_288; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_289 = io_pipe_phv_in_data_289; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_290 = io_pipe_phv_in_data_290; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_291 = io_pipe_phv_in_data_291; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_292 = io_pipe_phv_in_data_292; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_293 = io_pipe_phv_in_data_293; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_294 = io_pipe_phv_in_data_294; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_295 = io_pipe_phv_in_data_295; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_296 = io_pipe_phv_in_data_296; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_297 = io_pipe_phv_in_data_297; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_298 = io_pipe_phv_in_data_298; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_299 = io_pipe_phv_in_data_299; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_300 = io_pipe_phv_in_data_300; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_301 = io_pipe_phv_in_data_301; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_302 = io_pipe_phv_in_data_302; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_303 = io_pipe_phv_in_data_303; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_304 = io_pipe_phv_in_data_304; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_305 = io_pipe_phv_in_data_305; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_306 = io_pipe_phv_in_data_306; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_307 = io_pipe_phv_in_data_307; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_308 = io_pipe_phv_in_data_308; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_309 = io_pipe_phv_in_data_309; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_310 = io_pipe_phv_in_data_310; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_311 = io_pipe_phv_in_data_311; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_312 = io_pipe_phv_in_data_312; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_313 = io_pipe_phv_in_data_313; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_314 = io_pipe_phv_in_data_314; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_315 = io_pipe_phv_in_data_315; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_316 = io_pipe_phv_in_data_316; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_317 = io_pipe_phv_in_data_317; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_318 = io_pipe_phv_in_data_318; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_319 = io_pipe_phv_in_data_319; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_320 = io_pipe_phv_in_data_320; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_321 = io_pipe_phv_in_data_321; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_322 = io_pipe_phv_in_data_322; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_323 = io_pipe_phv_in_data_323; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_324 = io_pipe_phv_in_data_324; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_325 = io_pipe_phv_in_data_325; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_326 = io_pipe_phv_in_data_326; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_327 = io_pipe_phv_in_data_327; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_328 = io_pipe_phv_in_data_328; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_329 = io_pipe_phv_in_data_329; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_330 = io_pipe_phv_in_data_330; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_331 = io_pipe_phv_in_data_331; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_332 = io_pipe_phv_in_data_332; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_333 = io_pipe_phv_in_data_333; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_334 = io_pipe_phv_in_data_334; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_335 = io_pipe_phv_in_data_335; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_336 = io_pipe_phv_in_data_336; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_337 = io_pipe_phv_in_data_337; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_338 = io_pipe_phv_in_data_338; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_339 = io_pipe_phv_in_data_339; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_340 = io_pipe_phv_in_data_340; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_341 = io_pipe_phv_in_data_341; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_342 = io_pipe_phv_in_data_342; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_343 = io_pipe_phv_in_data_343; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_344 = io_pipe_phv_in_data_344; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_345 = io_pipe_phv_in_data_345; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_346 = io_pipe_phv_in_data_346; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_347 = io_pipe_phv_in_data_347; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_348 = io_pipe_phv_in_data_348; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_349 = io_pipe_phv_in_data_349; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_350 = io_pipe_phv_in_data_350; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_351 = io_pipe_phv_in_data_351; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_352 = io_pipe_phv_in_data_352; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_353 = io_pipe_phv_in_data_353; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_354 = io_pipe_phv_in_data_354; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_355 = io_pipe_phv_in_data_355; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_356 = io_pipe_phv_in_data_356; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_357 = io_pipe_phv_in_data_357; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_358 = io_pipe_phv_in_data_358; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_359 = io_pipe_phv_in_data_359; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_360 = io_pipe_phv_in_data_360; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_361 = io_pipe_phv_in_data_361; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_362 = io_pipe_phv_in_data_362; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_363 = io_pipe_phv_in_data_363; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_364 = io_pipe_phv_in_data_364; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_365 = io_pipe_phv_in_data_365; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_366 = io_pipe_phv_in_data_366; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_367 = io_pipe_phv_in_data_367; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_368 = io_pipe_phv_in_data_368; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_369 = io_pipe_phv_in_data_369; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_370 = io_pipe_phv_in_data_370; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_371 = io_pipe_phv_in_data_371; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_372 = io_pipe_phv_in_data_372; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_373 = io_pipe_phv_in_data_373; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_374 = io_pipe_phv_in_data_374; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_375 = io_pipe_phv_in_data_375; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_376 = io_pipe_phv_in_data_376; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_377 = io_pipe_phv_in_data_377; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_378 = io_pipe_phv_in_data_378; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_379 = io_pipe_phv_in_data_379; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_380 = io_pipe_phv_in_data_380; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_381 = io_pipe_phv_in_data_381; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_382 = io_pipe_phv_in_data_382; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_383 = io_pipe_phv_in_data_383; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_384 = io_pipe_phv_in_data_384; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_385 = io_pipe_phv_in_data_385; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_386 = io_pipe_phv_in_data_386; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_387 = io_pipe_phv_in_data_387; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_388 = io_pipe_phv_in_data_388; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_389 = io_pipe_phv_in_data_389; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_390 = io_pipe_phv_in_data_390; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_391 = io_pipe_phv_in_data_391; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_392 = io_pipe_phv_in_data_392; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_393 = io_pipe_phv_in_data_393; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_394 = io_pipe_phv_in_data_394; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_395 = io_pipe_phv_in_data_395; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_396 = io_pipe_phv_in_data_396; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_397 = io_pipe_phv_in_data_397; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_398 = io_pipe_phv_in_data_398; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_399 = io_pipe_phv_in_data_399; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_400 = io_pipe_phv_in_data_400; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_401 = io_pipe_phv_in_data_401; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_402 = io_pipe_phv_in_data_402; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_403 = io_pipe_phv_in_data_403; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_404 = io_pipe_phv_in_data_404; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_405 = io_pipe_phv_in_data_405; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_406 = io_pipe_phv_in_data_406; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_407 = io_pipe_phv_in_data_407; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_408 = io_pipe_phv_in_data_408; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_409 = io_pipe_phv_in_data_409; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_410 = io_pipe_phv_in_data_410; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_411 = io_pipe_phv_in_data_411; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_412 = io_pipe_phv_in_data_412; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_413 = io_pipe_phv_in_data_413; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_414 = io_pipe_phv_in_data_414; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_415 = io_pipe_phv_in_data_415; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_416 = io_pipe_phv_in_data_416; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_417 = io_pipe_phv_in_data_417; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_418 = io_pipe_phv_in_data_418; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_419 = io_pipe_phv_in_data_419; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_420 = io_pipe_phv_in_data_420; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_421 = io_pipe_phv_in_data_421; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_422 = io_pipe_phv_in_data_422; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_423 = io_pipe_phv_in_data_423; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_424 = io_pipe_phv_in_data_424; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_425 = io_pipe_phv_in_data_425; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_426 = io_pipe_phv_in_data_426; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_427 = io_pipe_phv_in_data_427; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_428 = io_pipe_phv_in_data_428; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_429 = io_pipe_phv_in_data_429; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_430 = io_pipe_phv_in_data_430; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_431 = io_pipe_phv_in_data_431; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_432 = io_pipe_phv_in_data_432; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_433 = io_pipe_phv_in_data_433; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_434 = io_pipe_phv_in_data_434; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_435 = io_pipe_phv_in_data_435; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_436 = io_pipe_phv_in_data_436; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_437 = io_pipe_phv_in_data_437; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_438 = io_pipe_phv_in_data_438; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_439 = io_pipe_phv_in_data_439; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_440 = io_pipe_phv_in_data_440; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_441 = io_pipe_phv_in_data_441; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_442 = io_pipe_phv_in_data_442; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_443 = io_pipe_phv_in_data_443; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_444 = io_pipe_phv_in_data_444; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_445 = io_pipe_phv_in_data_445; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_446 = io_pipe_phv_in_data_446; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_447 = io_pipe_phv_in_data_447; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_448 = io_pipe_phv_in_data_448; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_449 = io_pipe_phv_in_data_449; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_450 = io_pipe_phv_in_data_450; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_451 = io_pipe_phv_in_data_451; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_452 = io_pipe_phv_in_data_452; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_453 = io_pipe_phv_in_data_453; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_454 = io_pipe_phv_in_data_454; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_455 = io_pipe_phv_in_data_455; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_456 = io_pipe_phv_in_data_456; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_457 = io_pipe_phv_in_data_457; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_458 = io_pipe_phv_in_data_458; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_459 = io_pipe_phv_in_data_459; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_460 = io_pipe_phv_in_data_460; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_461 = io_pipe_phv_in_data_461; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_462 = io_pipe_phv_in_data_462; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_463 = io_pipe_phv_in_data_463; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_464 = io_pipe_phv_in_data_464; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_465 = io_pipe_phv_in_data_465; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_466 = io_pipe_phv_in_data_466; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_467 = io_pipe_phv_in_data_467; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_468 = io_pipe_phv_in_data_468; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_469 = io_pipe_phv_in_data_469; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_470 = io_pipe_phv_in_data_470; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_471 = io_pipe_phv_in_data_471; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_472 = io_pipe_phv_in_data_472; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_473 = io_pipe_phv_in_data_473; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_474 = io_pipe_phv_in_data_474; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_475 = io_pipe_phv_in_data_475; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_476 = io_pipe_phv_in_data_476; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_477 = io_pipe_phv_in_data_477; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_478 = io_pipe_phv_in_data_478; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_479 = io_pipe_phv_in_data_479; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_480 = io_pipe_phv_in_data_480; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_481 = io_pipe_phv_in_data_481; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_482 = io_pipe_phv_in_data_482; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_483 = io_pipe_phv_in_data_483; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_484 = io_pipe_phv_in_data_484; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_485 = io_pipe_phv_in_data_485; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_486 = io_pipe_phv_in_data_486; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_487 = io_pipe_phv_in_data_487; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_488 = io_pipe_phv_in_data_488; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_489 = io_pipe_phv_in_data_489; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_490 = io_pipe_phv_in_data_490; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_491 = io_pipe_phv_in_data_491; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_492 = io_pipe_phv_in_data_492; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_493 = io_pipe_phv_in_data_493; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_494 = io_pipe_phv_in_data_494; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_495 = io_pipe_phv_in_data_495; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_496 = io_pipe_phv_in_data_496; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_497 = io_pipe_phv_in_data_497; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_498 = io_pipe_phv_in_data_498; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_499 = io_pipe_phv_in_data_499; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_500 = io_pipe_phv_in_data_500; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_501 = io_pipe_phv_in_data_501; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_502 = io_pipe_phv_in_data_502; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_503 = io_pipe_phv_in_data_503; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_504 = io_pipe_phv_in_data_504; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_505 = io_pipe_phv_in_data_505; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_506 = io_pipe_phv_in_data_506; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_507 = io_pipe_phv_in_data_507; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_508 = io_pipe_phv_in_data_508; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_509 = io_pipe_phv_in_data_509; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_510 = io_pipe_phv_in_data_510; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_data_511 = io_pipe_phv_in_data_511; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_next_processor_id = io_pipe_phv_in_next_processor_id; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_next_config_id = io_pipe_phv_in_next_config_id; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_pipe_phv_in_is_valid_processor = io_pipe_phv_in_is_valid_processor; // @[matcher_pisa.scala 338:26]
  assign pipe1_io_key_config_0_field_config_0 = key_config_0_field_config_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_config_1 = key_config_0_field_config_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_config_2 = key_config_0_field_config_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_config_3 = key_config_0_field_config_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_config_4 = key_config_0_field_config_4; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_config_5 = key_config_0_field_config_5; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_0_0 = key_config_0_field_mask_0_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_0_1 = key_config_0_field_mask_0_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_0_2 = key_config_0_field_mask_0_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_0_3 = key_config_0_field_mask_0_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_1_0 = key_config_0_field_mask_1_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_1_1 = key_config_0_field_mask_1_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_1_2 = key_config_0_field_mask_1_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_1_3 = key_config_0_field_mask_1_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_2_0 = key_config_0_field_mask_2_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_2_1 = key_config_0_field_mask_2_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_2_2 = key_config_0_field_mask_2_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_2_3 = key_config_0_field_mask_2_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_3_0 = key_config_0_field_mask_3_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_3_1 = key_config_0_field_mask_3_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_3_2 = key_config_0_field_mask_3_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_3_3 = key_config_0_field_mask_3_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_4_0 = key_config_0_field_mask_4_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_4_1 = key_config_0_field_mask_4_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_4_2 = key_config_0_field_mask_4_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_4_3 = key_config_0_field_mask_4_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_5_0 = key_config_0_field_mask_5_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_5_1 = key_config_0_field_mask_5_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_5_2 = key_config_0_field_mask_5_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_mask_5_3 = key_config_0_field_mask_5_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_0_0 = key_config_0_field_id_0_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_0_1 = key_config_0_field_id_0_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_0_2 = key_config_0_field_id_0_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_0_3 = key_config_0_field_id_0_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_1_0 = key_config_0_field_id_1_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_1_1 = key_config_0_field_id_1_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_1_2 = key_config_0_field_id_1_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_1_3 = key_config_0_field_id_1_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_2_0 = key_config_0_field_id_2_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_2_1 = key_config_0_field_id_2_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_2_2 = key_config_0_field_id_2_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_2_3 = key_config_0_field_id_2_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_3_0 = key_config_0_field_id_3_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_3_1 = key_config_0_field_id_3_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_3_2 = key_config_0_field_id_3_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_3_3 = key_config_0_field_id_3_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_4_0 = key_config_0_field_id_4_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_4_1 = key_config_0_field_id_4_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_4_2 = key_config_0_field_id_4_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_4_3 = key_config_0_field_id_4_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_5_0 = key_config_0_field_id_5_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_5_1 = key_config_0_field_id_5_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_5_2 = key_config_0_field_id_5_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_0_field_id_5_3 = key_config_0_field_id_5_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_config_0 = key_config_1_field_config_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_config_1 = key_config_1_field_config_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_config_2 = key_config_1_field_config_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_config_3 = key_config_1_field_config_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_config_4 = key_config_1_field_config_4; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_config_5 = key_config_1_field_config_5; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_0_0 = key_config_1_field_mask_0_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_0_1 = key_config_1_field_mask_0_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_0_2 = key_config_1_field_mask_0_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_0_3 = key_config_1_field_mask_0_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_1_0 = key_config_1_field_mask_1_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_1_1 = key_config_1_field_mask_1_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_1_2 = key_config_1_field_mask_1_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_1_3 = key_config_1_field_mask_1_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_2_0 = key_config_1_field_mask_2_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_2_1 = key_config_1_field_mask_2_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_2_2 = key_config_1_field_mask_2_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_2_3 = key_config_1_field_mask_2_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_3_0 = key_config_1_field_mask_3_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_3_1 = key_config_1_field_mask_3_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_3_2 = key_config_1_field_mask_3_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_3_3 = key_config_1_field_mask_3_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_4_0 = key_config_1_field_mask_4_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_4_1 = key_config_1_field_mask_4_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_4_2 = key_config_1_field_mask_4_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_4_3 = key_config_1_field_mask_4_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_5_0 = key_config_1_field_mask_5_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_5_1 = key_config_1_field_mask_5_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_5_2 = key_config_1_field_mask_5_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_mask_5_3 = key_config_1_field_mask_5_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_0_0 = key_config_1_field_id_0_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_0_1 = key_config_1_field_id_0_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_0_2 = key_config_1_field_id_0_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_0_3 = key_config_1_field_id_0_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_1_0 = key_config_1_field_id_1_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_1_1 = key_config_1_field_id_1_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_1_2 = key_config_1_field_id_1_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_1_3 = key_config_1_field_id_1_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_2_0 = key_config_1_field_id_2_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_2_1 = key_config_1_field_id_2_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_2_2 = key_config_1_field_id_2_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_2_3 = key_config_1_field_id_2_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_3_0 = key_config_1_field_id_3_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_3_1 = key_config_1_field_id_3_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_3_2 = key_config_1_field_id_3_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_3_3 = key_config_1_field_id_3_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_4_0 = key_config_1_field_id_4_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_4_1 = key_config_1_field_id_4_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_4_2 = key_config_1_field_id_4_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_4_3 = key_config_1_field_id_4_3; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_5_0 = key_config_1_field_id_5_0; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_5_1 = key_config_1_field_id_5_1; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_5_2 = key_config_1_field_id_5_2; // @[matcher_pisa.scala 339:26]
  assign pipe1_io_key_config_1_field_id_5_3 = key_config_1_field_id_5_3; // @[matcher_pisa.scala 339:26]
  assign pipe2_clock = clock;
  assign pipe2_io_pipe_phv_in_data_0 = pipe1_io_pipe_phv_out_data_0; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_1 = pipe1_io_pipe_phv_out_data_1; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_2 = pipe1_io_pipe_phv_out_data_2; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_3 = pipe1_io_pipe_phv_out_data_3; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_4 = pipe1_io_pipe_phv_out_data_4; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_5 = pipe1_io_pipe_phv_out_data_5; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_6 = pipe1_io_pipe_phv_out_data_6; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_7 = pipe1_io_pipe_phv_out_data_7; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_8 = pipe1_io_pipe_phv_out_data_8; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_9 = pipe1_io_pipe_phv_out_data_9; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_10 = pipe1_io_pipe_phv_out_data_10; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_11 = pipe1_io_pipe_phv_out_data_11; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_12 = pipe1_io_pipe_phv_out_data_12; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_13 = pipe1_io_pipe_phv_out_data_13; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_14 = pipe1_io_pipe_phv_out_data_14; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_15 = pipe1_io_pipe_phv_out_data_15; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_16 = pipe1_io_pipe_phv_out_data_16; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_17 = pipe1_io_pipe_phv_out_data_17; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_18 = pipe1_io_pipe_phv_out_data_18; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_19 = pipe1_io_pipe_phv_out_data_19; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_20 = pipe1_io_pipe_phv_out_data_20; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_21 = pipe1_io_pipe_phv_out_data_21; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_22 = pipe1_io_pipe_phv_out_data_22; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_23 = pipe1_io_pipe_phv_out_data_23; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_24 = pipe1_io_pipe_phv_out_data_24; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_25 = pipe1_io_pipe_phv_out_data_25; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_26 = pipe1_io_pipe_phv_out_data_26; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_27 = pipe1_io_pipe_phv_out_data_27; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_28 = pipe1_io_pipe_phv_out_data_28; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_29 = pipe1_io_pipe_phv_out_data_29; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_30 = pipe1_io_pipe_phv_out_data_30; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_31 = pipe1_io_pipe_phv_out_data_31; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_32 = pipe1_io_pipe_phv_out_data_32; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_33 = pipe1_io_pipe_phv_out_data_33; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_34 = pipe1_io_pipe_phv_out_data_34; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_35 = pipe1_io_pipe_phv_out_data_35; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_36 = pipe1_io_pipe_phv_out_data_36; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_37 = pipe1_io_pipe_phv_out_data_37; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_38 = pipe1_io_pipe_phv_out_data_38; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_39 = pipe1_io_pipe_phv_out_data_39; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_40 = pipe1_io_pipe_phv_out_data_40; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_41 = pipe1_io_pipe_phv_out_data_41; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_42 = pipe1_io_pipe_phv_out_data_42; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_43 = pipe1_io_pipe_phv_out_data_43; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_44 = pipe1_io_pipe_phv_out_data_44; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_45 = pipe1_io_pipe_phv_out_data_45; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_46 = pipe1_io_pipe_phv_out_data_46; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_47 = pipe1_io_pipe_phv_out_data_47; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_48 = pipe1_io_pipe_phv_out_data_48; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_49 = pipe1_io_pipe_phv_out_data_49; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_50 = pipe1_io_pipe_phv_out_data_50; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_51 = pipe1_io_pipe_phv_out_data_51; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_52 = pipe1_io_pipe_phv_out_data_52; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_53 = pipe1_io_pipe_phv_out_data_53; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_54 = pipe1_io_pipe_phv_out_data_54; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_55 = pipe1_io_pipe_phv_out_data_55; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_56 = pipe1_io_pipe_phv_out_data_56; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_57 = pipe1_io_pipe_phv_out_data_57; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_58 = pipe1_io_pipe_phv_out_data_58; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_59 = pipe1_io_pipe_phv_out_data_59; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_60 = pipe1_io_pipe_phv_out_data_60; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_61 = pipe1_io_pipe_phv_out_data_61; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_62 = pipe1_io_pipe_phv_out_data_62; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_63 = pipe1_io_pipe_phv_out_data_63; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_64 = pipe1_io_pipe_phv_out_data_64; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_65 = pipe1_io_pipe_phv_out_data_65; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_66 = pipe1_io_pipe_phv_out_data_66; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_67 = pipe1_io_pipe_phv_out_data_67; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_68 = pipe1_io_pipe_phv_out_data_68; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_69 = pipe1_io_pipe_phv_out_data_69; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_70 = pipe1_io_pipe_phv_out_data_70; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_71 = pipe1_io_pipe_phv_out_data_71; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_72 = pipe1_io_pipe_phv_out_data_72; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_73 = pipe1_io_pipe_phv_out_data_73; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_74 = pipe1_io_pipe_phv_out_data_74; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_75 = pipe1_io_pipe_phv_out_data_75; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_76 = pipe1_io_pipe_phv_out_data_76; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_77 = pipe1_io_pipe_phv_out_data_77; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_78 = pipe1_io_pipe_phv_out_data_78; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_79 = pipe1_io_pipe_phv_out_data_79; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_80 = pipe1_io_pipe_phv_out_data_80; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_81 = pipe1_io_pipe_phv_out_data_81; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_82 = pipe1_io_pipe_phv_out_data_82; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_83 = pipe1_io_pipe_phv_out_data_83; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_84 = pipe1_io_pipe_phv_out_data_84; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_85 = pipe1_io_pipe_phv_out_data_85; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_86 = pipe1_io_pipe_phv_out_data_86; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_87 = pipe1_io_pipe_phv_out_data_87; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_88 = pipe1_io_pipe_phv_out_data_88; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_89 = pipe1_io_pipe_phv_out_data_89; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_90 = pipe1_io_pipe_phv_out_data_90; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_91 = pipe1_io_pipe_phv_out_data_91; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_92 = pipe1_io_pipe_phv_out_data_92; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_93 = pipe1_io_pipe_phv_out_data_93; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_94 = pipe1_io_pipe_phv_out_data_94; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_95 = pipe1_io_pipe_phv_out_data_95; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_96 = pipe1_io_pipe_phv_out_data_96; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_97 = pipe1_io_pipe_phv_out_data_97; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_98 = pipe1_io_pipe_phv_out_data_98; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_99 = pipe1_io_pipe_phv_out_data_99; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_100 = pipe1_io_pipe_phv_out_data_100; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_101 = pipe1_io_pipe_phv_out_data_101; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_102 = pipe1_io_pipe_phv_out_data_102; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_103 = pipe1_io_pipe_phv_out_data_103; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_104 = pipe1_io_pipe_phv_out_data_104; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_105 = pipe1_io_pipe_phv_out_data_105; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_106 = pipe1_io_pipe_phv_out_data_106; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_107 = pipe1_io_pipe_phv_out_data_107; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_108 = pipe1_io_pipe_phv_out_data_108; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_109 = pipe1_io_pipe_phv_out_data_109; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_110 = pipe1_io_pipe_phv_out_data_110; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_111 = pipe1_io_pipe_phv_out_data_111; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_112 = pipe1_io_pipe_phv_out_data_112; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_113 = pipe1_io_pipe_phv_out_data_113; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_114 = pipe1_io_pipe_phv_out_data_114; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_115 = pipe1_io_pipe_phv_out_data_115; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_116 = pipe1_io_pipe_phv_out_data_116; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_117 = pipe1_io_pipe_phv_out_data_117; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_118 = pipe1_io_pipe_phv_out_data_118; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_119 = pipe1_io_pipe_phv_out_data_119; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_120 = pipe1_io_pipe_phv_out_data_120; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_121 = pipe1_io_pipe_phv_out_data_121; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_122 = pipe1_io_pipe_phv_out_data_122; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_123 = pipe1_io_pipe_phv_out_data_123; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_124 = pipe1_io_pipe_phv_out_data_124; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_125 = pipe1_io_pipe_phv_out_data_125; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_126 = pipe1_io_pipe_phv_out_data_126; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_127 = pipe1_io_pipe_phv_out_data_127; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_128 = pipe1_io_pipe_phv_out_data_128; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_129 = pipe1_io_pipe_phv_out_data_129; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_130 = pipe1_io_pipe_phv_out_data_130; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_131 = pipe1_io_pipe_phv_out_data_131; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_132 = pipe1_io_pipe_phv_out_data_132; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_133 = pipe1_io_pipe_phv_out_data_133; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_134 = pipe1_io_pipe_phv_out_data_134; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_135 = pipe1_io_pipe_phv_out_data_135; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_136 = pipe1_io_pipe_phv_out_data_136; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_137 = pipe1_io_pipe_phv_out_data_137; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_138 = pipe1_io_pipe_phv_out_data_138; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_139 = pipe1_io_pipe_phv_out_data_139; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_140 = pipe1_io_pipe_phv_out_data_140; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_141 = pipe1_io_pipe_phv_out_data_141; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_142 = pipe1_io_pipe_phv_out_data_142; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_143 = pipe1_io_pipe_phv_out_data_143; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_144 = pipe1_io_pipe_phv_out_data_144; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_145 = pipe1_io_pipe_phv_out_data_145; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_146 = pipe1_io_pipe_phv_out_data_146; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_147 = pipe1_io_pipe_phv_out_data_147; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_148 = pipe1_io_pipe_phv_out_data_148; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_149 = pipe1_io_pipe_phv_out_data_149; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_150 = pipe1_io_pipe_phv_out_data_150; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_151 = pipe1_io_pipe_phv_out_data_151; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_152 = pipe1_io_pipe_phv_out_data_152; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_153 = pipe1_io_pipe_phv_out_data_153; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_154 = pipe1_io_pipe_phv_out_data_154; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_155 = pipe1_io_pipe_phv_out_data_155; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_156 = pipe1_io_pipe_phv_out_data_156; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_157 = pipe1_io_pipe_phv_out_data_157; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_158 = pipe1_io_pipe_phv_out_data_158; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_159 = pipe1_io_pipe_phv_out_data_159; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_160 = pipe1_io_pipe_phv_out_data_160; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_161 = pipe1_io_pipe_phv_out_data_161; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_162 = pipe1_io_pipe_phv_out_data_162; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_163 = pipe1_io_pipe_phv_out_data_163; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_164 = pipe1_io_pipe_phv_out_data_164; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_165 = pipe1_io_pipe_phv_out_data_165; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_166 = pipe1_io_pipe_phv_out_data_166; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_167 = pipe1_io_pipe_phv_out_data_167; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_168 = pipe1_io_pipe_phv_out_data_168; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_169 = pipe1_io_pipe_phv_out_data_169; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_170 = pipe1_io_pipe_phv_out_data_170; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_171 = pipe1_io_pipe_phv_out_data_171; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_172 = pipe1_io_pipe_phv_out_data_172; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_173 = pipe1_io_pipe_phv_out_data_173; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_174 = pipe1_io_pipe_phv_out_data_174; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_175 = pipe1_io_pipe_phv_out_data_175; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_176 = pipe1_io_pipe_phv_out_data_176; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_177 = pipe1_io_pipe_phv_out_data_177; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_178 = pipe1_io_pipe_phv_out_data_178; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_179 = pipe1_io_pipe_phv_out_data_179; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_180 = pipe1_io_pipe_phv_out_data_180; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_181 = pipe1_io_pipe_phv_out_data_181; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_182 = pipe1_io_pipe_phv_out_data_182; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_183 = pipe1_io_pipe_phv_out_data_183; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_184 = pipe1_io_pipe_phv_out_data_184; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_185 = pipe1_io_pipe_phv_out_data_185; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_186 = pipe1_io_pipe_phv_out_data_186; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_187 = pipe1_io_pipe_phv_out_data_187; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_188 = pipe1_io_pipe_phv_out_data_188; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_189 = pipe1_io_pipe_phv_out_data_189; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_190 = pipe1_io_pipe_phv_out_data_190; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_191 = pipe1_io_pipe_phv_out_data_191; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_192 = pipe1_io_pipe_phv_out_data_192; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_193 = pipe1_io_pipe_phv_out_data_193; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_194 = pipe1_io_pipe_phv_out_data_194; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_195 = pipe1_io_pipe_phv_out_data_195; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_196 = pipe1_io_pipe_phv_out_data_196; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_197 = pipe1_io_pipe_phv_out_data_197; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_198 = pipe1_io_pipe_phv_out_data_198; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_199 = pipe1_io_pipe_phv_out_data_199; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_200 = pipe1_io_pipe_phv_out_data_200; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_201 = pipe1_io_pipe_phv_out_data_201; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_202 = pipe1_io_pipe_phv_out_data_202; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_203 = pipe1_io_pipe_phv_out_data_203; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_204 = pipe1_io_pipe_phv_out_data_204; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_205 = pipe1_io_pipe_phv_out_data_205; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_206 = pipe1_io_pipe_phv_out_data_206; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_207 = pipe1_io_pipe_phv_out_data_207; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_208 = pipe1_io_pipe_phv_out_data_208; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_209 = pipe1_io_pipe_phv_out_data_209; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_210 = pipe1_io_pipe_phv_out_data_210; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_211 = pipe1_io_pipe_phv_out_data_211; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_212 = pipe1_io_pipe_phv_out_data_212; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_213 = pipe1_io_pipe_phv_out_data_213; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_214 = pipe1_io_pipe_phv_out_data_214; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_215 = pipe1_io_pipe_phv_out_data_215; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_216 = pipe1_io_pipe_phv_out_data_216; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_217 = pipe1_io_pipe_phv_out_data_217; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_218 = pipe1_io_pipe_phv_out_data_218; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_219 = pipe1_io_pipe_phv_out_data_219; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_220 = pipe1_io_pipe_phv_out_data_220; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_221 = pipe1_io_pipe_phv_out_data_221; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_222 = pipe1_io_pipe_phv_out_data_222; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_223 = pipe1_io_pipe_phv_out_data_223; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_224 = pipe1_io_pipe_phv_out_data_224; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_225 = pipe1_io_pipe_phv_out_data_225; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_226 = pipe1_io_pipe_phv_out_data_226; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_227 = pipe1_io_pipe_phv_out_data_227; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_228 = pipe1_io_pipe_phv_out_data_228; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_229 = pipe1_io_pipe_phv_out_data_229; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_230 = pipe1_io_pipe_phv_out_data_230; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_231 = pipe1_io_pipe_phv_out_data_231; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_232 = pipe1_io_pipe_phv_out_data_232; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_233 = pipe1_io_pipe_phv_out_data_233; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_234 = pipe1_io_pipe_phv_out_data_234; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_235 = pipe1_io_pipe_phv_out_data_235; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_236 = pipe1_io_pipe_phv_out_data_236; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_237 = pipe1_io_pipe_phv_out_data_237; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_238 = pipe1_io_pipe_phv_out_data_238; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_239 = pipe1_io_pipe_phv_out_data_239; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_240 = pipe1_io_pipe_phv_out_data_240; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_241 = pipe1_io_pipe_phv_out_data_241; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_242 = pipe1_io_pipe_phv_out_data_242; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_243 = pipe1_io_pipe_phv_out_data_243; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_244 = pipe1_io_pipe_phv_out_data_244; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_245 = pipe1_io_pipe_phv_out_data_245; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_246 = pipe1_io_pipe_phv_out_data_246; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_247 = pipe1_io_pipe_phv_out_data_247; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_248 = pipe1_io_pipe_phv_out_data_248; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_249 = pipe1_io_pipe_phv_out_data_249; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_250 = pipe1_io_pipe_phv_out_data_250; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_251 = pipe1_io_pipe_phv_out_data_251; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_252 = pipe1_io_pipe_phv_out_data_252; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_253 = pipe1_io_pipe_phv_out_data_253; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_254 = pipe1_io_pipe_phv_out_data_254; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_255 = pipe1_io_pipe_phv_out_data_255; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_256 = pipe1_io_pipe_phv_out_data_256; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_257 = pipe1_io_pipe_phv_out_data_257; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_258 = pipe1_io_pipe_phv_out_data_258; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_259 = pipe1_io_pipe_phv_out_data_259; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_260 = pipe1_io_pipe_phv_out_data_260; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_261 = pipe1_io_pipe_phv_out_data_261; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_262 = pipe1_io_pipe_phv_out_data_262; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_263 = pipe1_io_pipe_phv_out_data_263; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_264 = pipe1_io_pipe_phv_out_data_264; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_265 = pipe1_io_pipe_phv_out_data_265; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_266 = pipe1_io_pipe_phv_out_data_266; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_267 = pipe1_io_pipe_phv_out_data_267; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_268 = pipe1_io_pipe_phv_out_data_268; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_269 = pipe1_io_pipe_phv_out_data_269; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_270 = pipe1_io_pipe_phv_out_data_270; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_271 = pipe1_io_pipe_phv_out_data_271; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_272 = pipe1_io_pipe_phv_out_data_272; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_273 = pipe1_io_pipe_phv_out_data_273; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_274 = pipe1_io_pipe_phv_out_data_274; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_275 = pipe1_io_pipe_phv_out_data_275; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_276 = pipe1_io_pipe_phv_out_data_276; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_277 = pipe1_io_pipe_phv_out_data_277; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_278 = pipe1_io_pipe_phv_out_data_278; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_279 = pipe1_io_pipe_phv_out_data_279; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_280 = pipe1_io_pipe_phv_out_data_280; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_281 = pipe1_io_pipe_phv_out_data_281; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_282 = pipe1_io_pipe_phv_out_data_282; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_283 = pipe1_io_pipe_phv_out_data_283; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_284 = pipe1_io_pipe_phv_out_data_284; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_285 = pipe1_io_pipe_phv_out_data_285; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_286 = pipe1_io_pipe_phv_out_data_286; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_287 = pipe1_io_pipe_phv_out_data_287; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_288 = pipe1_io_pipe_phv_out_data_288; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_289 = pipe1_io_pipe_phv_out_data_289; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_290 = pipe1_io_pipe_phv_out_data_290; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_291 = pipe1_io_pipe_phv_out_data_291; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_292 = pipe1_io_pipe_phv_out_data_292; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_293 = pipe1_io_pipe_phv_out_data_293; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_294 = pipe1_io_pipe_phv_out_data_294; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_295 = pipe1_io_pipe_phv_out_data_295; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_296 = pipe1_io_pipe_phv_out_data_296; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_297 = pipe1_io_pipe_phv_out_data_297; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_298 = pipe1_io_pipe_phv_out_data_298; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_299 = pipe1_io_pipe_phv_out_data_299; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_300 = pipe1_io_pipe_phv_out_data_300; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_301 = pipe1_io_pipe_phv_out_data_301; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_302 = pipe1_io_pipe_phv_out_data_302; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_303 = pipe1_io_pipe_phv_out_data_303; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_304 = pipe1_io_pipe_phv_out_data_304; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_305 = pipe1_io_pipe_phv_out_data_305; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_306 = pipe1_io_pipe_phv_out_data_306; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_307 = pipe1_io_pipe_phv_out_data_307; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_308 = pipe1_io_pipe_phv_out_data_308; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_309 = pipe1_io_pipe_phv_out_data_309; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_310 = pipe1_io_pipe_phv_out_data_310; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_311 = pipe1_io_pipe_phv_out_data_311; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_312 = pipe1_io_pipe_phv_out_data_312; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_313 = pipe1_io_pipe_phv_out_data_313; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_314 = pipe1_io_pipe_phv_out_data_314; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_315 = pipe1_io_pipe_phv_out_data_315; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_316 = pipe1_io_pipe_phv_out_data_316; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_317 = pipe1_io_pipe_phv_out_data_317; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_318 = pipe1_io_pipe_phv_out_data_318; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_319 = pipe1_io_pipe_phv_out_data_319; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_320 = pipe1_io_pipe_phv_out_data_320; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_321 = pipe1_io_pipe_phv_out_data_321; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_322 = pipe1_io_pipe_phv_out_data_322; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_323 = pipe1_io_pipe_phv_out_data_323; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_324 = pipe1_io_pipe_phv_out_data_324; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_325 = pipe1_io_pipe_phv_out_data_325; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_326 = pipe1_io_pipe_phv_out_data_326; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_327 = pipe1_io_pipe_phv_out_data_327; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_328 = pipe1_io_pipe_phv_out_data_328; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_329 = pipe1_io_pipe_phv_out_data_329; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_330 = pipe1_io_pipe_phv_out_data_330; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_331 = pipe1_io_pipe_phv_out_data_331; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_332 = pipe1_io_pipe_phv_out_data_332; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_333 = pipe1_io_pipe_phv_out_data_333; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_334 = pipe1_io_pipe_phv_out_data_334; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_335 = pipe1_io_pipe_phv_out_data_335; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_336 = pipe1_io_pipe_phv_out_data_336; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_337 = pipe1_io_pipe_phv_out_data_337; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_338 = pipe1_io_pipe_phv_out_data_338; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_339 = pipe1_io_pipe_phv_out_data_339; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_340 = pipe1_io_pipe_phv_out_data_340; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_341 = pipe1_io_pipe_phv_out_data_341; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_342 = pipe1_io_pipe_phv_out_data_342; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_343 = pipe1_io_pipe_phv_out_data_343; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_344 = pipe1_io_pipe_phv_out_data_344; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_345 = pipe1_io_pipe_phv_out_data_345; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_346 = pipe1_io_pipe_phv_out_data_346; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_347 = pipe1_io_pipe_phv_out_data_347; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_348 = pipe1_io_pipe_phv_out_data_348; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_349 = pipe1_io_pipe_phv_out_data_349; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_350 = pipe1_io_pipe_phv_out_data_350; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_351 = pipe1_io_pipe_phv_out_data_351; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_352 = pipe1_io_pipe_phv_out_data_352; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_353 = pipe1_io_pipe_phv_out_data_353; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_354 = pipe1_io_pipe_phv_out_data_354; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_355 = pipe1_io_pipe_phv_out_data_355; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_356 = pipe1_io_pipe_phv_out_data_356; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_357 = pipe1_io_pipe_phv_out_data_357; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_358 = pipe1_io_pipe_phv_out_data_358; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_359 = pipe1_io_pipe_phv_out_data_359; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_360 = pipe1_io_pipe_phv_out_data_360; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_361 = pipe1_io_pipe_phv_out_data_361; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_362 = pipe1_io_pipe_phv_out_data_362; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_363 = pipe1_io_pipe_phv_out_data_363; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_364 = pipe1_io_pipe_phv_out_data_364; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_365 = pipe1_io_pipe_phv_out_data_365; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_366 = pipe1_io_pipe_phv_out_data_366; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_367 = pipe1_io_pipe_phv_out_data_367; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_368 = pipe1_io_pipe_phv_out_data_368; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_369 = pipe1_io_pipe_phv_out_data_369; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_370 = pipe1_io_pipe_phv_out_data_370; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_371 = pipe1_io_pipe_phv_out_data_371; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_372 = pipe1_io_pipe_phv_out_data_372; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_373 = pipe1_io_pipe_phv_out_data_373; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_374 = pipe1_io_pipe_phv_out_data_374; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_375 = pipe1_io_pipe_phv_out_data_375; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_376 = pipe1_io_pipe_phv_out_data_376; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_377 = pipe1_io_pipe_phv_out_data_377; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_378 = pipe1_io_pipe_phv_out_data_378; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_379 = pipe1_io_pipe_phv_out_data_379; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_380 = pipe1_io_pipe_phv_out_data_380; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_381 = pipe1_io_pipe_phv_out_data_381; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_382 = pipe1_io_pipe_phv_out_data_382; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_383 = pipe1_io_pipe_phv_out_data_383; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_384 = pipe1_io_pipe_phv_out_data_384; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_385 = pipe1_io_pipe_phv_out_data_385; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_386 = pipe1_io_pipe_phv_out_data_386; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_387 = pipe1_io_pipe_phv_out_data_387; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_388 = pipe1_io_pipe_phv_out_data_388; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_389 = pipe1_io_pipe_phv_out_data_389; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_390 = pipe1_io_pipe_phv_out_data_390; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_391 = pipe1_io_pipe_phv_out_data_391; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_392 = pipe1_io_pipe_phv_out_data_392; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_393 = pipe1_io_pipe_phv_out_data_393; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_394 = pipe1_io_pipe_phv_out_data_394; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_395 = pipe1_io_pipe_phv_out_data_395; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_396 = pipe1_io_pipe_phv_out_data_396; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_397 = pipe1_io_pipe_phv_out_data_397; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_398 = pipe1_io_pipe_phv_out_data_398; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_399 = pipe1_io_pipe_phv_out_data_399; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_400 = pipe1_io_pipe_phv_out_data_400; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_401 = pipe1_io_pipe_phv_out_data_401; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_402 = pipe1_io_pipe_phv_out_data_402; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_403 = pipe1_io_pipe_phv_out_data_403; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_404 = pipe1_io_pipe_phv_out_data_404; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_405 = pipe1_io_pipe_phv_out_data_405; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_406 = pipe1_io_pipe_phv_out_data_406; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_407 = pipe1_io_pipe_phv_out_data_407; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_408 = pipe1_io_pipe_phv_out_data_408; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_409 = pipe1_io_pipe_phv_out_data_409; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_410 = pipe1_io_pipe_phv_out_data_410; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_411 = pipe1_io_pipe_phv_out_data_411; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_412 = pipe1_io_pipe_phv_out_data_412; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_413 = pipe1_io_pipe_phv_out_data_413; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_414 = pipe1_io_pipe_phv_out_data_414; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_415 = pipe1_io_pipe_phv_out_data_415; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_416 = pipe1_io_pipe_phv_out_data_416; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_417 = pipe1_io_pipe_phv_out_data_417; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_418 = pipe1_io_pipe_phv_out_data_418; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_419 = pipe1_io_pipe_phv_out_data_419; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_420 = pipe1_io_pipe_phv_out_data_420; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_421 = pipe1_io_pipe_phv_out_data_421; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_422 = pipe1_io_pipe_phv_out_data_422; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_423 = pipe1_io_pipe_phv_out_data_423; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_424 = pipe1_io_pipe_phv_out_data_424; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_425 = pipe1_io_pipe_phv_out_data_425; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_426 = pipe1_io_pipe_phv_out_data_426; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_427 = pipe1_io_pipe_phv_out_data_427; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_428 = pipe1_io_pipe_phv_out_data_428; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_429 = pipe1_io_pipe_phv_out_data_429; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_430 = pipe1_io_pipe_phv_out_data_430; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_431 = pipe1_io_pipe_phv_out_data_431; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_432 = pipe1_io_pipe_phv_out_data_432; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_433 = pipe1_io_pipe_phv_out_data_433; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_434 = pipe1_io_pipe_phv_out_data_434; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_435 = pipe1_io_pipe_phv_out_data_435; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_436 = pipe1_io_pipe_phv_out_data_436; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_437 = pipe1_io_pipe_phv_out_data_437; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_438 = pipe1_io_pipe_phv_out_data_438; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_439 = pipe1_io_pipe_phv_out_data_439; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_440 = pipe1_io_pipe_phv_out_data_440; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_441 = pipe1_io_pipe_phv_out_data_441; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_442 = pipe1_io_pipe_phv_out_data_442; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_443 = pipe1_io_pipe_phv_out_data_443; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_444 = pipe1_io_pipe_phv_out_data_444; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_445 = pipe1_io_pipe_phv_out_data_445; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_446 = pipe1_io_pipe_phv_out_data_446; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_447 = pipe1_io_pipe_phv_out_data_447; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_448 = pipe1_io_pipe_phv_out_data_448; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_449 = pipe1_io_pipe_phv_out_data_449; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_450 = pipe1_io_pipe_phv_out_data_450; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_451 = pipe1_io_pipe_phv_out_data_451; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_452 = pipe1_io_pipe_phv_out_data_452; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_453 = pipe1_io_pipe_phv_out_data_453; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_454 = pipe1_io_pipe_phv_out_data_454; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_455 = pipe1_io_pipe_phv_out_data_455; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_456 = pipe1_io_pipe_phv_out_data_456; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_457 = pipe1_io_pipe_phv_out_data_457; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_458 = pipe1_io_pipe_phv_out_data_458; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_459 = pipe1_io_pipe_phv_out_data_459; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_460 = pipe1_io_pipe_phv_out_data_460; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_461 = pipe1_io_pipe_phv_out_data_461; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_462 = pipe1_io_pipe_phv_out_data_462; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_463 = pipe1_io_pipe_phv_out_data_463; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_464 = pipe1_io_pipe_phv_out_data_464; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_465 = pipe1_io_pipe_phv_out_data_465; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_466 = pipe1_io_pipe_phv_out_data_466; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_467 = pipe1_io_pipe_phv_out_data_467; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_468 = pipe1_io_pipe_phv_out_data_468; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_469 = pipe1_io_pipe_phv_out_data_469; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_470 = pipe1_io_pipe_phv_out_data_470; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_471 = pipe1_io_pipe_phv_out_data_471; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_472 = pipe1_io_pipe_phv_out_data_472; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_473 = pipe1_io_pipe_phv_out_data_473; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_474 = pipe1_io_pipe_phv_out_data_474; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_475 = pipe1_io_pipe_phv_out_data_475; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_476 = pipe1_io_pipe_phv_out_data_476; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_477 = pipe1_io_pipe_phv_out_data_477; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_478 = pipe1_io_pipe_phv_out_data_478; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_479 = pipe1_io_pipe_phv_out_data_479; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_480 = pipe1_io_pipe_phv_out_data_480; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_481 = pipe1_io_pipe_phv_out_data_481; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_482 = pipe1_io_pipe_phv_out_data_482; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_483 = pipe1_io_pipe_phv_out_data_483; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_484 = pipe1_io_pipe_phv_out_data_484; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_485 = pipe1_io_pipe_phv_out_data_485; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_486 = pipe1_io_pipe_phv_out_data_486; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_487 = pipe1_io_pipe_phv_out_data_487; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_488 = pipe1_io_pipe_phv_out_data_488; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_489 = pipe1_io_pipe_phv_out_data_489; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_490 = pipe1_io_pipe_phv_out_data_490; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_491 = pipe1_io_pipe_phv_out_data_491; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_492 = pipe1_io_pipe_phv_out_data_492; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_493 = pipe1_io_pipe_phv_out_data_493; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_494 = pipe1_io_pipe_phv_out_data_494; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_495 = pipe1_io_pipe_phv_out_data_495; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_496 = pipe1_io_pipe_phv_out_data_496; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_497 = pipe1_io_pipe_phv_out_data_497; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_498 = pipe1_io_pipe_phv_out_data_498; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_499 = pipe1_io_pipe_phv_out_data_499; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_500 = pipe1_io_pipe_phv_out_data_500; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_501 = pipe1_io_pipe_phv_out_data_501; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_502 = pipe1_io_pipe_phv_out_data_502; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_503 = pipe1_io_pipe_phv_out_data_503; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_504 = pipe1_io_pipe_phv_out_data_504; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_505 = pipe1_io_pipe_phv_out_data_505; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_506 = pipe1_io_pipe_phv_out_data_506; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_507 = pipe1_io_pipe_phv_out_data_507; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_508 = pipe1_io_pipe_phv_out_data_508; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_509 = pipe1_io_pipe_phv_out_data_509; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_510 = pipe1_io_pipe_phv_out_data_510; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_data_511 = pipe1_io_pipe_phv_out_data_511; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_next_processor_id = pipe1_io_pipe_phv_out_next_processor_id; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_next_config_id = pipe1_io_pipe_phv_out_next_config_id; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_pipe_phv_in_is_valid_processor = pipe1_io_pipe_phv_out_is_valid_processor; // @[matcher_pisa.scala 341:26]
  assign pipe2_io_mod_hash_depth_mod = io_mod_en; // @[matcher_pisa.scala 342:33]
  assign pipe2_io_mod_config_id = io_mod_config_id; // @[matcher_pisa.scala 343:28]
  assign pipe2_io_mod_hash_depth = io_mod_table_mod_table_depth[3:0]; // @[matcher_pisa.scala 344:29]
  assign pipe2_io_key_in = pipe1_io_match_key; // @[matcher_pisa.scala 345:26]
  assign pipe3_clock = clock;
  assign pipe3_io_pipe_phv_in_data_0 = pipe2_io_pipe_phv_out_data_0; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_1 = pipe2_io_pipe_phv_out_data_1; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_2 = pipe2_io_pipe_phv_out_data_2; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_3 = pipe2_io_pipe_phv_out_data_3; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_4 = pipe2_io_pipe_phv_out_data_4; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_5 = pipe2_io_pipe_phv_out_data_5; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_6 = pipe2_io_pipe_phv_out_data_6; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_7 = pipe2_io_pipe_phv_out_data_7; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_8 = pipe2_io_pipe_phv_out_data_8; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_9 = pipe2_io_pipe_phv_out_data_9; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_10 = pipe2_io_pipe_phv_out_data_10; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_11 = pipe2_io_pipe_phv_out_data_11; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_12 = pipe2_io_pipe_phv_out_data_12; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_13 = pipe2_io_pipe_phv_out_data_13; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_14 = pipe2_io_pipe_phv_out_data_14; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_15 = pipe2_io_pipe_phv_out_data_15; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_16 = pipe2_io_pipe_phv_out_data_16; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_17 = pipe2_io_pipe_phv_out_data_17; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_18 = pipe2_io_pipe_phv_out_data_18; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_19 = pipe2_io_pipe_phv_out_data_19; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_20 = pipe2_io_pipe_phv_out_data_20; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_21 = pipe2_io_pipe_phv_out_data_21; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_22 = pipe2_io_pipe_phv_out_data_22; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_23 = pipe2_io_pipe_phv_out_data_23; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_24 = pipe2_io_pipe_phv_out_data_24; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_25 = pipe2_io_pipe_phv_out_data_25; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_26 = pipe2_io_pipe_phv_out_data_26; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_27 = pipe2_io_pipe_phv_out_data_27; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_28 = pipe2_io_pipe_phv_out_data_28; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_29 = pipe2_io_pipe_phv_out_data_29; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_30 = pipe2_io_pipe_phv_out_data_30; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_31 = pipe2_io_pipe_phv_out_data_31; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_32 = pipe2_io_pipe_phv_out_data_32; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_33 = pipe2_io_pipe_phv_out_data_33; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_34 = pipe2_io_pipe_phv_out_data_34; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_35 = pipe2_io_pipe_phv_out_data_35; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_36 = pipe2_io_pipe_phv_out_data_36; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_37 = pipe2_io_pipe_phv_out_data_37; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_38 = pipe2_io_pipe_phv_out_data_38; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_39 = pipe2_io_pipe_phv_out_data_39; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_40 = pipe2_io_pipe_phv_out_data_40; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_41 = pipe2_io_pipe_phv_out_data_41; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_42 = pipe2_io_pipe_phv_out_data_42; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_43 = pipe2_io_pipe_phv_out_data_43; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_44 = pipe2_io_pipe_phv_out_data_44; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_45 = pipe2_io_pipe_phv_out_data_45; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_46 = pipe2_io_pipe_phv_out_data_46; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_47 = pipe2_io_pipe_phv_out_data_47; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_48 = pipe2_io_pipe_phv_out_data_48; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_49 = pipe2_io_pipe_phv_out_data_49; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_50 = pipe2_io_pipe_phv_out_data_50; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_51 = pipe2_io_pipe_phv_out_data_51; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_52 = pipe2_io_pipe_phv_out_data_52; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_53 = pipe2_io_pipe_phv_out_data_53; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_54 = pipe2_io_pipe_phv_out_data_54; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_55 = pipe2_io_pipe_phv_out_data_55; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_56 = pipe2_io_pipe_phv_out_data_56; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_57 = pipe2_io_pipe_phv_out_data_57; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_58 = pipe2_io_pipe_phv_out_data_58; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_59 = pipe2_io_pipe_phv_out_data_59; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_60 = pipe2_io_pipe_phv_out_data_60; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_61 = pipe2_io_pipe_phv_out_data_61; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_62 = pipe2_io_pipe_phv_out_data_62; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_63 = pipe2_io_pipe_phv_out_data_63; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_64 = pipe2_io_pipe_phv_out_data_64; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_65 = pipe2_io_pipe_phv_out_data_65; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_66 = pipe2_io_pipe_phv_out_data_66; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_67 = pipe2_io_pipe_phv_out_data_67; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_68 = pipe2_io_pipe_phv_out_data_68; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_69 = pipe2_io_pipe_phv_out_data_69; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_70 = pipe2_io_pipe_phv_out_data_70; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_71 = pipe2_io_pipe_phv_out_data_71; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_72 = pipe2_io_pipe_phv_out_data_72; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_73 = pipe2_io_pipe_phv_out_data_73; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_74 = pipe2_io_pipe_phv_out_data_74; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_75 = pipe2_io_pipe_phv_out_data_75; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_76 = pipe2_io_pipe_phv_out_data_76; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_77 = pipe2_io_pipe_phv_out_data_77; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_78 = pipe2_io_pipe_phv_out_data_78; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_79 = pipe2_io_pipe_phv_out_data_79; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_80 = pipe2_io_pipe_phv_out_data_80; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_81 = pipe2_io_pipe_phv_out_data_81; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_82 = pipe2_io_pipe_phv_out_data_82; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_83 = pipe2_io_pipe_phv_out_data_83; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_84 = pipe2_io_pipe_phv_out_data_84; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_85 = pipe2_io_pipe_phv_out_data_85; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_86 = pipe2_io_pipe_phv_out_data_86; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_87 = pipe2_io_pipe_phv_out_data_87; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_88 = pipe2_io_pipe_phv_out_data_88; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_89 = pipe2_io_pipe_phv_out_data_89; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_90 = pipe2_io_pipe_phv_out_data_90; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_91 = pipe2_io_pipe_phv_out_data_91; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_92 = pipe2_io_pipe_phv_out_data_92; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_93 = pipe2_io_pipe_phv_out_data_93; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_94 = pipe2_io_pipe_phv_out_data_94; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_95 = pipe2_io_pipe_phv_out_data_95; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_96 = pipe2_io_pipe_phv_out_data_96; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_97 = pipe2_io_pipe_phv_out_data_97; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_98 = pipe2_io_pipe_phv_out_data_98; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_99 = pipe2_io_pipe_phv_out_data_99; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_100 = pipe2_io_pipe_phv_out_data_100; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_101 = pipe2_io_pipe_phv_out_data_101; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_102 = pipe2_io_pipe_phv_out_data_102; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_103 = pipe2_io_pipe_phv_out_data_103; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_104 = pipe2_io_pipe_phv_out_data_104; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_105 = pipe2_io_pipe_phv_out_data_105; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_106 = pipe2_io_pipe_phv_out_data_106; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_107 = pipe2_io_pipe_phv_out_data_107; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_108 = pipe2_io_pipe_phv_out_data_108; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_109 = pipe2_io_pipe_phv_out_data_109; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_110 = pipe2_io_pipe_phv_out_data_110; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_111 = pipe2_io_pipe_phv_out_data_111; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_112 = pipe2_io_pipe_phv_out_data_112; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_113 = pipe2_io_pipe_phv_out_data_113; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_114 = pipe2_io_pipe_phv_out_data_114; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_115 = pipe2_io_pipe_phv_out_data_115; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_116 = pipe2_io_pipe_phv_out_data_116; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_117 = pipe2_io_pipe_phv_out_data_117; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_118 = pipe2_io_pipe_phv_out_data_118; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_119 = pipe2_io_pipe_phv_out_data_119; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_120 = pipe2_io_pipe_phv_out_data_120; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_121 = pipe2_io_pipe_phv_out_data_121; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_122 = pipe2_io_pipe_phv_out_data_122; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_123 = pipe2_io_pipe_phv_out_data_123; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_124 = pipe2_io_pipe_phv_out_data_124; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_125 = pipe2_io_pipe_phv_out_data_125; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_126 = pipe2_io_pipe_phv_out_data_126; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_127 = pipe2_io_pipe_phv_out_data_127; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_128 = pipe2_io_pipe_phv_out_data_128; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_129 = pipe2_io_pipe_phv_out_data_129; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_130 = pipe2_io_pipe_phv_out_data_130; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_131 = pipe2_io_pipe_phv_out_data_131; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_132 = pipe2_io_pipe_phv_out_data_132; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_133 = pipe2_io_pipe_phv_out_data_133; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_134 = pipe2_io_pipe_phv_out_data_134; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_135 = pipe2_io_pipe_phv_out_data_135; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_136 = pipe2_io_pipe_phv_out_data_136; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_137 = pipe2_io_pipe_phv_out_data_137; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_138 = pipe2_io_pipe_phv_out_data_138; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_139 = pipe2_io_pipe_phv_out_data_139; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_140 = pipe2_io_pipe_phv_out_data_140; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_141 = pipe2_io_pipe_phv_out_data_141; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_142 = pipe2_io_pipe_phv_out_data_142; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_143 = pipe2_io_pipe_phv_out_data_143; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_144 = pipe2_io_pipe_phv_out_data_144; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_145 = pipe2_io_pipe_phv_out_data_145; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_146 = pipe2_io_pipe_phv_out_data_146; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_147 = pipe2_io_pipe_phv_out_data_147; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_148 = pipe2_io_pipe_phv_out_data_148; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_149 = pipe2_io_pipe_phv_out_data_149; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_150 = pipe2_io_pipe_phv_out_data_150; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_151 = pipe2_io_pipe_phv_out_data_151; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_152 = pipe2_io_pipe_phv_out_data_152; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_153 = pipe2_io_pipe_phv_out_data_153; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_154 = pipe2_io_pipe_phv_out_data_154; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_155 = pipe2_io_pipe_phv_out_data_155; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_156 = pipe2_io_pipe_phv_out_data_156; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_157 = pipe2_io_pipe_phv_out_data_157; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_158 = pipe2_io_pipe_phv_out_data_158; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_159 = pipe2_io_pipe_phv_out_data_159; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_160 = pipe2_io_pipe_phv_out_data_160; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_161 = pipe2_io_pipe_phv_out_data_161; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_162 = pipe2_io_pipe_phv_out_data_162; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_163 = pipe2_io_pipe_phv_out_data_163; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_164 = pipe2_io_pipe_phv_out_data_164; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_165 = pipe2_io_pipe_phv_out_data_165; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_166 = pipe2_io_pipe_phv_out_data_166; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_167 = pipe2_io_pipe_phv_out_data_167; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_168 = pipe2_io_pipe_phv_out_data_168; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_169 = pipe2_io_pipe_phv_out_data_169; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_170 = pipe2_io_pipe_phv_out_data_170; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_171 = pipe2_io_pipe_phv_out_data_171; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_172 = pipe2_io_pipe_phv_out_data_172; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_173 = pipe2_io_pipe_phv_out_data_173; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_174 = pipe2_io_pipe_phv_out_data_174; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_175 = pipe2_io_pipe_phv_out_data_175; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_176 = pipe2_io_pipe_phv_out_data_176; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_177 = pipe2_io_pipe_phv_out_data_177; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_178 = pipe2_io_pipe_phv_out_data_178; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_179 = pipe2_io_pipe_phv_out_data_179; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_180 = pipe2_io_pipe_phv_out_data_180; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_181 = pipe2_io_pipe_phv_out_data_181; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_182 = pipe2_io_pipe_phv_out_data_182; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_183 = pipe2_io_pipe_phv_out_data_183; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_184 = pipe2_io_pipe_phv_out_data_184; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_185 = pipe2_io_pipe_phv_out_data_185; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_186 = pipe2_io_pipe_phv_out_data_186; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_187 = pipe2_io_pipe_phv_out_data_187; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_188 = pipe2_io_pipe_phv_out_data_188; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_189 = pipe2_io_pipe_phv_out_data_189; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_190 = pipe2_io_pipe_phv_out_data_190; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_191 = pipe2_io_pipe_phv_out_data_191; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_192 = pipe2_io_pipe_phv_out_data_192; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_193 = pipe2_io_pipe_phv_out_data_193; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_194 = pipe2_io_pipe_phv_out_data_194; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_195 = pipe2_io_pipe_phv_out_data_195; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_196 = pipe2_io_pipe_phv_out_data_196; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_197 = pipe2_io_pipe_phv_out_data_197; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_198 = pipe2_io_pipe_phv_out_data_198; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_199 = pipe2_io_pipe_phv_out_data_199; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_200 = pipe2_io_pipe_phv_out_data_200; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_201 = pipe2_io_pipe_phv_out_data_201; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_202 = pipe2_io_pipe_phv_out_data_202; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_203 = pipe2_io_pipe_phv_out_data_203; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_204 = pipe2_io_pipe_phv_out_data_204; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_205 = pipe2_io_pipe_phv_out_data_205; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_206 = pipe2_io_pipe_phv_out_data_206; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_207 = pipe2_io_pipe_phv_out_data_207; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_208 = pipe2_io_pipe_phv_out_data_208; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_209 = pipe2_io_pipe_phv_out_data_209; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_210 = pipe2_io_pipe_phv_out_data_210; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_211 = pipe2_io_pipe_phv_out_data_211; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_212 = pipe2_io_pipe_phv_out_data_212; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_213 = pipe2_io_pipe_phv_out_data_213; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_214 = pipe2_io_pipe_phv_out_data_214; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_215 = pipe2_io_pipe_phv_out_data_215; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_216 = pipe2_io_pipe_phv_out_data_216; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_217 = pipe2_io_pipe_phv_out_data_217; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_218 = pipe2_io_pipe_phv_out_data_218; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_219 = pipe2_io_pipe_phv_out_data_219; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_220 = pipe2_io_pipe_phv_out_data_220; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_221 = pipe2_io_pipe_phv_out_data_221; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_222 = pipe2_io_pipe_phv_out_data_222; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_223 = pipe2_io_pipe_phv_out_data_223; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_224 = pipe2_io_pipe_phv_out_data_224; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_225 = pipe2_io_pipe_phv_out_data_225; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_226 = pipe2_io_pipe_phv_out_data_226; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_227 = pipe2_io_pipe_phv_out_data_227; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_228 = pipe2_io_pipe_phv_out_data_228; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_229 = pipe2_io_pipe_phv_out_data_229; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_230 = pipe2_io_pipe_phv_out_data_230; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_231 = pipe2_io_pipe_phv_out_data_231; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_232 = pipe2_io_pipe_phv_out_data_232; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_233 = pipe2_io_pipe_phv_out_data_233; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_234 = pipe2_io_pipe_phv_out_data_234; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_235 = pipe2_io_pipe_phv_out_data_235; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_236 = pipe2_io_pipe_phv_out_data_236; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_237 = pipe2_io_pipe_phv_out_data_237; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_238 = pipe2_io_pipe_phv_out_data_238; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_239 = pipe2_io_pipe_phv_out_data_239; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_240 = pipe2_io_pipe_phv_out_data_240; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_241 = pipe2_io_pipe_phv_out_data_241; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_242 = pipe2_io_pipe_phv_out_data_242; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_243 = pipe2_io_pipe_phv_out_data_243; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_244 = pipe2_io_pipe_phv_out_data_244; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_245 = pipe2_io_pipe_phv_out_data_245; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_246 = pipe2_io_pipe_phv_out_data_246; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_247 = pipe2_io_pipe_phv_out_data_247; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_248 = pipe2_io_pipe_phv_out_data_248; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_249 = pipe2_io_pipe_phv_out_data_249; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_250 = pipe2_io_pipe_phv_out_data_250; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_251 = pipe2_io_pipe_phv_out_data_251; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_252 = pipe2_io_pipe_phv_out_data_252; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_253 = pipe2_io_pipe_phv_out_data_253; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_254 = pipe2_io_pipe_phv_out_data_254; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_255 = pipe2_io_pipe_phv_out_data_255; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_256 = pipe2_io_pipe_phv_out_data_256; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_257 = pipe2_io_pipe_phv_out_data_257; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_258 = pipe2_io_pipe_phv_out_data_258; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_259 = pipe2_io_pipe_phv_out_data_259; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_260 = pipe2_io_pipe_phv_out_data_260; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_261 = pipe2_io_pipe_phv_out_data_261; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_262 = pipe2_io_pipe_phv_out_data_262; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_263 = pipe2_io_pipe_phv_out_data_263; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_264 = pipe2_io_pipe_phv_out_data_264; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_265 = pipe2_io_pipe_phv_out_data_265; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_266 = pipe2_io_pipe_phv_out_data_266; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_267 = pipe2_io_pipe_phv_out_data_267; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_268 = pipe2_io_pipe_phv_out_data_268; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_269 = pipe2_io_pipe_phv_out_data_269; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_270 = pipe2_io_pipe_phv_out_data_270; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_271 = pipe2_io_pipe_phv_out_data_271; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_272 = pipe2_io_pipe_phv_out_data_272; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_273 = pipe2_io_pipe_phv_out_data_273; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_274 = pipe2_io_pipe_phv_out_data_274; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_275 = pipe2_io_pipe_phv_out_data_275; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_276 = pipe2_io_pipe_phv_out_data_276; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_277 = pipe2_io_pipe_phv_out_data_277; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_278 = pipe2_io_pipe_phv_out_data_278; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_279 = pipe2_io_pipe_phv_out_data_279; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_280 = pipe2_io_pipe_phv_out_data_280; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_281 = pipe2_io_pipe_phv_out_data_281; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_282 = pipe2_io_pipe_phv_out_data_282; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_283 = pipe2_io_pipe_phv_out_data_283; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_284 = pipe2_io_pipe_phv_out_data_284; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_285 = pipe2_io_pipe_phv_out_data_285; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_286 = pipe2_io_pipe_phv_out_data_286; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_287 = pipe2_io_pipe_phv_out_data_287; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_288 = pipe2_io_pipe_phv_out_data_288; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_289 = pipe2_io_pipe_phv_out_data_289; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_290 = pipe2_io_pipe_phv_out_data_290; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_291 = pipe2_io_pipe_phv_out_data_291; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_292 = pipe2_io_pipe_phv_out_data_292; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_293 = pipe2_io_pipe_phv_out_data_293; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_294 = pipe2_io_pipe_phv_out_data_294; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_295 = pipe2_io_pipe_phv_out_data_295; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_296 = pipe2_io_pipe_phv_out_data_296; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_297 = pipe2_io_pipe_phv_out_data_297; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_298 = pipe2_io_pipe_phv_out_data_298; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_299 = pipe2_io_pipe_phv_out_data_299; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_300 = pipe2_io_pipe_phv_out_data_300; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_301 = pipe2_io_pipe_phv_out_data_301; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_302 = pipe2_io_pipe_phv_out_data_302; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_303 = pipe2_io_pipe_phv_out_data_303; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_304 = pipe2_io_pipe_phv_out_data_304; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_305 = pipe2_io_pipe_phv_out_data_305; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_306 = pipe2_io_pipe_phv_out_data_306; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_307 = pipe2_io_pipe_phv_out_data_307; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_308 = pipe2_io_pipe_phv_out_data_308; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_309 = pipe2_io_pipe_phv_out_data_309; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_310 = pipe2_io_pipe_phv_out_data_310; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_311 = pipe2_io_pipe_phv_out_data_311; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_312 = pipe2_io_pipe_phv_out_data_312; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_313 = pipe2_io_pipe_phv_out_data_313; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_314 = pipe2_io_pipe_phv_out_data_314; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_315 = pipe2_io_pipe_phv_out_data_315; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_316 = pipe2_io_pipe_phv_out_data_316; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_317 = pipe2_io_pipe_phv_out_data_317; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_318 = pipe2_io_pipe_phv_out_data_318; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_319 = pipe2_io_pipe_phv_out_data_319; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_320 = pipe2_io_pipe_phv_out_data_320; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_321 = pipe2_io_pipe_phv_out_data_321; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_322 = pipe2_io_pipe_phv_out_data_322; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_323 = pipe2_io_pipe_phv_out_data_323; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_324 = pipe2_io_pipe_phv_out_data_324; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_325 = pipe2_io_pipe_phv_out_data_325; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_326 = pipe2_io_pipe_phv_out_data_326; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_327 = pipe2_io_pipe_phv_out_data_327; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_328 = pipe2_io_pipe_phv_out_data_328; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_329 = pipe2_io_pipe_phv_out_data_329; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_330 = pipe2_io_pipe_phv_out_data_330; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_331 = pipe2_io_pipe_phv_out_data_331; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_332 = pipe2_io_pipe_phv_out_data_332; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_333 = pipe2_io_pipe_phv_out_data_333; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_334 = pipe2_io_pipe_phv_out_data_334; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_335 = pipe2_io_pipe_phv_out_data_335; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_336 = pipe2_io_pipe_phv_out_data_336; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_337 = pipe2_io_pipe_phv_out_data_337; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_338 = pipe2_io_pipe_phv_out_data_338; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_339 = pipe2_io_pipe_phv_out_data_339; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_340 = pipe2_io_pipe_phv_out_data_340; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_341 = pipe2_io_pipe_phv_out_data_341; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_342 = pipe2_io_pipe_phv_out_data_342; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_343 = pipe2_io_pipe_phv_out_data_343; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_344 = pipe2_io_pipe_phv_out_data_344; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_345 = pipe2_io_pipe_phv_out_data_345; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_346 = pipe2_io_pipe_phv_out_data_346; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_347 = pipe2_io_pipe_phv_out_data_347; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_348 = pipe2_io_pipe_phv_out_data_348; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_349 = pipe2_io_pipe_phv_out_data_349; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_350 = pipe2_io_pipe_phv_out_data_350; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_351 = pipe2_io_pipe_phv_out_data_351; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_352 = pipe2_io_pipe_phv_out_data_352; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_353 = pipe2_io_pipe_phv_out_data_353; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_354 = pipe2_io_pipe_phv_out_data_354; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_355 = pipe2_io_pipe_phv_out_data_355; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_356 = pipe2_io_pipe_phv_out_data_356; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_357 = pipe2_io_pipe_phv_out_data_357; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_358 = pipe2_io_pipe_phv_out_data_358; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_359 = pipe2_io_pipe_phv_out_data_359; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_360 = pipe2_io_pipe_phv_out_data_360; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_361 = pipe2_io_pipe_phv_out_data_361; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_362 = pipe2_io_pipe_phv_out_data_362; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_363 = pipe2_io_pipe_phv_out_data_363; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_364 = pipe2_io_pipe_phv_out_data_364; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_365 = pipe2_io_pipe_phv_out_data_365; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_366 = pipe2_io_pipe_phv_out_data_366; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_367 = pipe2_io_pipe_phv_out_data_367; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_368 = pipe2_io_pipe_phv_out_data_368; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_369 = pipe2_io_pipe_phv_out_data_369; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_370 = pipe2_io_pipe_phv_out_data_370; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_371 = pipe2_io_pipe_phv_out_data_371; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_372 = pipe2_io_pipe_phv_out_data_372; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_373 = pipe2_io_pipe_phv_out_data_373; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_374 = pipe2_io_pipe_phv_out_data_374; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_375 = pipe2_io_pipe_phv_out_data_375; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_376 = pipe2_io_pipe_phv_out_data_376; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_377 = pipe2_io_pipe_phv_out_data_377; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_378 = pipe2_io_pipe_phv_out_data_378; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_379 = pipe2_io_pipe_phv_out_data_379; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_380 = pipe2_io_pipe_phv_out_data_380; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_381 = pipe2_io_pipe_phv_out_data_381; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_382 = pipe2_io_pipe_phv_out_data_382; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_383 = pipe2_io_pipe_phv_out_data_383; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_384 = pipe2_io_pipe_phv_out_data_384; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_385 = pipe2_io_pipe_phv_out_data_385; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_386 = pipe2_io_pipe_phv_out_data_386; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_387 = pipe2_io_pipe_phv_out_data_387; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_388 = pipe2_io_pipe_phv_out_data_388; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_389 = pipe2_io_pipe_phv_out_data_389; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_390 = pipe2_io_pipe_phv_out_data_390; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_391 = pipe2_io_pipe_phv_out_data_391; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_392 = pipe2_io_pipe_phv_out_data_392; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_393 = pipe2_io_pipe_phv_out_data_393; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_394 = pipe2_io_pipe_phv_out_data_394; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_395 = pipe2_io_pipe_phv_out_data_395; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_396 = pipe2_io_pipe_phv_out_data_396; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_397 = pipe2_io_pipe_phv_out_data_397; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_398 = pipe2_io_pipe_phv_out_data_398; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_399 = pipe2_io_pipe_phv_out_data_399; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_400 = pipe2_io_pipe_phv_out_data_400; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_401 = pipe2_io_pipe_phv_out_data_401; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_402 = pipe2_io_pipe_phv_out_data_402; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_403 = pipe2_io_pipe_phv_out_data_403; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_404 = pipe2_io_pipe_phv_out_data_404; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_405 = pipe2_io_pipe_phv_out_data_405; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_406 = pipe2_io_pipe_phv_out_data_406; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_407 = pipe2_io_pipe_phv_out_data_407; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_408 = pipe2_io_pipe_phv_out_data_408; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_409 = pipe2_io_pipe_phv_out_data_409; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_410 = pipe2_io_pipe_phv_out_data_410; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_411 = pipe2_io_pipe_phv_out_data_411; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_412 = pipe2_io_pipe_phv_out_data_412; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_413 = pipe2_io_pipe_phv_out_data_413; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_414 = pipe2_io_pipe_phv_out_data_414; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_415 = pipe2_io_pipe_phv_out_data_415; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_416 = pipe2_io_pipe_phv_out_data_416; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_417 = pipe2_io_pipe_phv_out_data_417; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_418 = pipe2_io_pipe_phv_out_data_418; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_419 = pipe2_io_pipe_phv_out_data_419; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_420 = pipe2_io_pipe_phv_out_data_420; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_421 = pipe2_io_pipe_phv_out_data_421; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_422 = pipe2_io_pipe_phv_out_data_422; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_423 = pipe2_io_pipe_phv_out_data_423; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_424 = pipe2_io_pipe_phv_out_data_424; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_425 = pipe2_io_pipe_phv_out_data_425; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_426 = pipe2_io_pipe_phv_out_data_426; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_427 = pipe2_io_pipe_phv_out_data_427; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_428 = pipe2_io_pipe_phv_out_data_428; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_429 = pipe2_io_pipe_phv_out_data_429; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_430 = pipe2_io_pipe_phv_out_data_430; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_431 = pipe2_io_pipe_phv_out_data_431; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_432 = pipe2_io_pipe_phv_out_data_432; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_433 = pipe2_io_pipe_phv_out_data_433; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_434 = pipe2_io_pipe_phv_out_data_434; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_435 = pipe2_io_pipe_phv_out_data_435; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_436 = pipe2_io_pipe_phv_out_data_436; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_437 = pipe2_io_pipe_phv_out_data_437; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_438 = pipe2_io_pipe_phv_out_data_438; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_439 = pipe2_io_pipe_phv_out_data_439; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_440 = pipe2_io_pipe_phv_out_data_440; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_441 = pipe2_io_pipe_phv_out_data_441; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_442 = pipe2_io_pipe_phv_out_data_442; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_443 = pipe2_io_pipe_phv_out_data_443; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_444 = pipe2_io_pipe_phv_out_data_444; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_445 = pipe2_io_pipe_phv_out_data_445; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_446 = pipe2_io_pipe_phv_out_data_446; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_447 = pipe2_io_pipe_phv_out_data_447; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_448 = pipe2_io_pipe_phv_out_data_448; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_449 = pipe2_io_pipe_phv_out_data_449; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_450 = pipe2_io_pipe_phv_out_data_450; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_451 = pipe2_io_pipe_phv_out_data_451; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_452 = pipe2_io_pipe_phv_out_data_452; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_453 = pipe2_io_pipe_phv_out_data_453; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_454 = pipe2_io_pipe_phv_out_data_454; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_455 = pipe2_io_pipe_phv_out_data_455; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_456 = pipe2_io_pipe_phv_out_data_456; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_457 = pipe2_io_pipe_phv_out_data_457; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_458 = pipe2_io_pipe_phv_out_data_458; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_459 = pipe2_io_pipe_phv_out_data_459; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_460 = pipe2_io_pipe_phv_out_data_460; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_461 = pipe2_io_pipe_phv_out_data_461; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_462 = pipe2_io_pipe_phv_out_data_462; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_463 = pipe2_io_pipe_phv_out_data_463; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_464 = pipe2_io_pipe_phv_out_data_464; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_465 = pipe2_io_pipe_phv_out_data_465; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_466 = pipe2_io_pipe_phv_out_data_466; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_467 = pipe2_io_pipe_phv_out_data_467; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_468 = pipe2_io_pipe_phv_out_data_468; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_469 = pipe2_io_pipe_phv_out_data_469; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_470 = pipe2_io_pipe_phv_out_data_470; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_471 = pipe2_io_pipe_phv_out_data_471; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_472 = pipe2_io_pipe_phv_out_data_472; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_473 = pipe2_io_pipe_phv_out_data_473; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_474 = pipe2_io_pipe_phv_out_data_474; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_475 = pipe2_io_pipe_phv_out_data_475; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_476 = pipe2_io_pipe_phv_out_data_476; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_477 = pipe2_io_pipe_phv_out_data_477; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_478 = pipe2_io_pipe_phv_out_data_478; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_479 = pipe2_io_pipe_phv_out_data_479; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_480 = pipe2_io_pipe_phv_out_data_480; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_481 = pipe2_io_pipe_phv_out_data_481; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_482 = pipe2_io_pipe_phv_out_data_482; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_483 = pipe2_io_pipe_phv_out_data_483; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_484 = pipe2_io_pipe_phv_out_data_484; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_485 = pipe2_io_pipe_phv_out_data_485; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_486 = pipe2_io_pipe_phv_out_data_486; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_487 = pipe2_io_pipe_phv_out_data_487; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_488 = pipe2_io_pipe_phv_out_data_488; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_489 = pipe2_io_pipe_phv_out_data_489; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_490 = pipe2_io_pipe_phv_out_data_490; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_491 = pipe2_io_pipe_phv_out_data_491; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_492 = pipe2_io_pipe_phv_out_data_492; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_493 = pipe2_io_pipe_phv_out_data_493; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_494 = pipe2_io_pipe_phv_out_data_494; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_495 = pipe2_io_pipe_phv_out_data_495; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_496 = pipe2_io_pipe_phv_out_data_496; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_497 = pipe2_io_pipe_phv_out_data_497; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_498 = pipe2_io_pipe_phv_out_data_498; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_499 = pipe2_io_pipe_phv_out_data_499; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_500 = pipe2_io_pipe_phv_out_data_500; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_501 = pipe2_io_pipe_phv_out_data_501; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_502 = pipe2_io_pipe_phv_out_data_502; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_503 = pipe2_io_pipe_phv_out_data_503; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_504 = pipe2_io_pipe_phv_out_data_504; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_505 = pipe2_io_pipe_phv_out_data_505; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_506 = pipe2_io_pipe_phv_out_data_506; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_507 = pipe2_io_pipe_phv_out_data_507; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_508 = pipe2_io_pipe_phv_out_data_508; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_509 = pipe2_io_pipe_phv_out_data_509; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_510 = pipe2_io_pipe_phv_out_data_510; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_data_511 = pipe2_io_pipe_phv_out_data_511; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_next_processor_id = pipe2_io_pipe_phv_out_next_processor_id; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_next_config_id = pipe2_io_pipe_phv_out_next_config_id; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_pipe_phv_in_is_valid_processor = pipe2_io_pipe_phv_out_is_valid_processor; // @[matcher_pisa.scala 347:26]
  assign pipe3_io_table_config_0_table_depth = table_config_0_table_depth; // @[matcher_pisa.scala 348:27]
  assign pipe3_io_table_config_0_table_width = table_config_0_table_width; // @[matcher_pisa.scala 348:27]
  assign pipe3_io_table_config_1_table_depth = table_config_1_table_depth; // @[matcher_pisa.scala 348:27]
  assign pipe3_io_table_config_1_table_width = table_config_1_table_width; // @[matcher_pisa.scala 348:27]
  assign pipe3_io_key_in = pipe2_io_key_out; // @[matcher_pisa.scala 349:26]
  assign pipe3_io_addr_in = pipe2_io_hash_val; // @[matcher_pisa.scala 350:26]
  assign pipe3_io_cs_in = pipe2_io_hash_val_cs; // @[matcher_pisa.scala 351:26]
  assign pipe3_io_w_en = io_mod_w_en; // @[matcher_pisa.scala 352:26]
  assign pipe3_io_w_sram_id = io_mod_w_sram_id; // @[matcher_pisa.scala 352:26]
  assign pipe3_io_w_addr = io_mod_w_addr; // @[matcher_pisa.scala 352:26]
  assign pipe3_io_w_data = io_mod_w_data; // @[matcher_pisa.scala 352:26]
  assign pipe4_clock = clock;
  assign pipe4_io_pipe_phv_in_data_0 = pipe3_io_pipe_phv_out_data_0; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_1 = pipe3_io_pipe_phv_out_data_1; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_2 = pipe3_io_pipe_phv_out_data_2; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_3 = pipe3_io_pipe_phv_out_data_3; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_4 = pipe3_io_pipe_phv_out_data_4; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_5 = pipe3_io_pipe_phv_out_data_5; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_6 = pipe3_io_pipe_phv_out_data_6; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_7 = pipe3_io_pipe_phv_out_data_7; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_8 = pipe3_io_pipe_phv_out_data_8; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_9 = pipe3_io_pipe_phv_out_data_9; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_10 = pipe3_io_pipe_phv_out_data_10; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_11 = pipe3_io_pipe_phv_out_data_11; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_12 = pipe3_io_pipe_phv_out_data_12; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_13 = pipe3_io_pipe_phv_out_data_13; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_14 = pipe3_io_pipe_phv_out_data_14; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_15 = pipe3_io_pipe_phv_out_data_15; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_16 = pipe3_io_pipe_phv_out_data_16; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_17 = pipe3_io_pipe_phv_out_data_17; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_18 = pipe3_io_pipe_phv_out_data_18; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_19 = pipe3_io_pipe_phv_out_data_19; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_20 = pipe3_io_pipe_phv_out_data_20; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_21 = pipe3_io_pipe_phv_out_data_21; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_22 = pipe3_io_pipe_phv_out_data_22; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_23 = pipe3_io_pipe_phv_out_data_23; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_24 = pipe3_io_pipe_phv_out_data_24; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_25 = pipe3_io_pipe_phv_out_data_25; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_26 = pipe3_io_pipe_phv_out_data_26; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_27 = pipe3_io_pipe_phv_out_data_27; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_28 = pipe3_io_pipe_phv_out_data_28; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_29 = pipe3_io_pipe_phv_out_data_29; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_30 = pipe3_io_pipe_phv_out_data_30; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_31 = pipe3_io_pipe_phv_out_data_31; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_32 = pipe3_io_pipe_phv_out_data_32; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_33 = pipe3_io_pipe_phv_out_data_33; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_34 = pipe3_io_pipe_phv_out_data_34; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_35 = pipe3_io_pipe_phv_out_data_35; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_36 = pipe3_io_pipe_phv_out_data_36; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_37 = pipe3_io_pipe_phv_out_data_37; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_38 = pipe3_io_pipe_phv_out_data_38; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_39 = pipe3_io_pipe_phv_out_data_39; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_40 = pipe3_io_pipe_phv_out_data_40; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_41 = pipe3_io_pipe_phv_out_data_41; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_42 = pipe3_io_pipe_phv_out_data_42; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_43 = pipe3_io_pipe_phv_out_data_43; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_44 = pipe3_io_pipe_phv_out_data_44; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_45 = pipe3_io_pipe_phv_out_data_45; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_46 = pipe3_io_pipe_phv_out_data_46; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_47 = pipe3_io_pipe_phv_out_data_47; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_48 = pipe3_io_pipe_phv_out_data_48; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_49 = pipe3_io_pipe_phv_out_data_49; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_50 = pipe3_io_pipe_phv_out_data_50; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_51 = pipe3_io_pipe_phv_out_data_51; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_52 = pipe3_io_pipe_phv_out_data_52; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_53 = pipe3_io_pipe_phv_out_data_53; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_54 = pipe3_io_pipe_phv_out_data_54; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_55 = pipe3_io_pipe_phv_out_data_55; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_56 = pipe3_io_pipe_phv_out_data_56; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_57 = pipe3_io_pipe_phv_out_data_57; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_58 = pipe3_io_pipe_phv_out_data_58; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_59 = pipe3_io_pipe_phv_out_data_59; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_60 = pipe3_io_pipe_phv_out_data_60; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_61 = pipe3_io_pipe_phv_out_data_61; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_62 = pipe3_io_pipe_phv_out_data_62; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_63 = pipe3_io_pipe_phv_out_data_63; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_64 = pipe3_io_pipe_phv_out_data_64; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_65 = pipe3_io_pipe_phv_out_data_65; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_66 = pipe3_io_pipe_phv_out_data_66; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_67 = pipe3_io_pipe_phv_out_data_67; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_68 = pipe3_io_pipe_phv_out_data_68; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_69 = pipe3_io_pipe_phv_out_data_69; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_70 = pipe3_io_pipe_phv_out_data_70; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_71 = pipe3_io_pipe_phv_out_data_71; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_72 = pipe3_io_pipe_phv_out_data_72; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_73 = pipe3_io_pipe_phv_out_data_73; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_74 = pipe3_io_pipe_phv_out_data_74; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_75 = pipe3_io_pipe_phv_out_data_75; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_76 = pipe3_io_pipe_phv_out_data_76; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_77 = pipe3_io_pipe_phv_out_data_77; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_78 = pipe3_io_pipe_phv_out_data_78; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_79 = pipe3_io_pipe_phv_out_data_79; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_80 = pipe3_io_pipe_phv_out_data_80; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_81 = pipe3_io_pipe_phv_out_data_81; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_82 = pipe3_io_pipe_phv_out_data_82; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_83 = pipe3_io_pipe_phv_out_data_83; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_84 = pipe3_io_pipe_phv_out_data_84; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_85 = pipe3_io_pipe_phv_out_data_85; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_86 = pipe3_io_pipe_phv_out_data_86; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_87 = pipe3_io_pipe_phv_out_data_87; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_88 = pipe3_io_pipe_phv_out_data_88; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_89 = pipe3_io_pipe_phv_out_data_89; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_90 = pipe3_io_pipe_phv_out_data_90; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_91 = pipe3_io_pipe_phv_out_data_91; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_92 = pipe3_io_pipe_phv_out_data_92; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_93 = pipe3_io_pipe_phv_out_data_93; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_94 = pipe3_io_pipe_phv_out_data_94; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_95 = pipe3_io_pipe_phv_out_data_95; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_96 = pipe3_io_pipe_phv_out_data_96; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_97 = pipe3_io_pipe_phv_out_data_97; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_98 = pipe3_io_pipe_phv_out_data_98; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_99 = pipe3_io_pipe_phv_out_data_99; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_100 = pipe3_io_pipe_phv_out_data_100; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_101 = pipe3_io_pipe_phv_out_data_101; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_102 = pipe3_io_pipe_phv_out_data_102; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_103 = pipe3_io_pipe_phv_out_data_103; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_104 = pipe3_io_pipe_phv_out_data_104; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_105 = pipe3_io_pipe_phv_out_data_105; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_106 = pipe3_io_pipe_phv_out_data_106; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_107 = pipe3_io_pipe_phv_out_data_107; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_108 = pipe3_io_pipe_phv_out_data_108; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_109 = pipe3_io_pipe_phv_out_data_109; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_110 = pipe3_io_pipe_phv_out_data_110; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_111 = pipe3_io_pipe_phv_out_data_111; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_112 = pipe3_io_pipe_phv_out_data_112; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_113 = pipe3_io_pipe_phv_out_data_113; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_114 = pipe3_io_pipe_phv_out_data_114; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_115 = pipe3_io_pipe_phv_out_data_115; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_116 = pipe3_io_pipe_phv_out_data_116; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_117 = pipe3_io_pipe_phv_out_data_117; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_118 = pipe3_io_pipe_phv_out_data_118; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_119 = pipe3_io_pipe_phv_out_data_119; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_120 = pipe3_io_pipe_phv_out_data_120; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_121 = pipe3_io_pipe_phv_out_data_121; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_122 = pipe3_io_pipe_phv_out_data_122; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_123 = pipe3_io_pipe_phv_out_data_123; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_124 = pipe3_io_pipe_phv_out_data_124; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_125 = pipe3_io_pipe_phv_out_data_125; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_126 = pipe3_io_pipe_phv_out_data_126; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_127 = pipe3_io_pipe_phv_out_data_127; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_128 = pipe3_io_pipe_phv_out_data_128; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_129 = pipe3_io_pipe_phv_out_data_129; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_130 = pipe3_io_pipe_phv_out_data_130; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_131 = pipe3_io_pipe_phv_out_data_131; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_132 = pipe3_io_pipe_phv_out_data_132; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_133 = pipe3_io_pipe_phv_out_data_133; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_134 = pipe3_io_pipe_phv_out_data_134; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_135 = pipe3_io_pipe_phv_out_data_135; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_136 = pipe3_io_pipe_phv_out_data_136; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_137 = pipe3_io_pipe_phv_out_data_137; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_138 = pipe3_io_pipe_phv_out_data_138; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_139 = pipe3_io_pipe_phv_out_data_139; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_140 = pipe3_io_pipe_phv_out_data_140; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_141 = pipe3_io_pipe_phv_out_data_141; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_142 = pipe3_io_pipe_phv_out_data_142; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_143 = pipe3_io_pipe_phv_out_data_143; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_144 = pipe3_io_pipe_phv_out_data_144; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_145 = pipe3_io_pipe_phv_out_data_145; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_146 = pipe3_io_pipe_phv_out_data_146; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_147 = pipe3_io_pipe_phv_out_data_147; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_148 = pipe3_io_pipe_phv_out_data_148; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_149 = pipe3_io_pipe_phv_out_data_149; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_150 = pipe3_io_pipe_phv_out_data_150; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_151 = pipe3_io_pipe_phv_out_data_151; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_152 = pipe3_io_pipe_phv_out_data_152; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_153 = pipe3_io_pipe_phv_out_data_153; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_154 = pipe3_io_pipe_phv_out_data_154; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_155 = pipe3_io_pipe_phv_out_data_155; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_156 = pipe3_io_pipe_phv_out_data_156; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_157 = pipe3_io_pipe_phv_out_data_157; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_158 = pipe3_io_pipe_phv_out_data_158; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_159 = pipe3_io_pipe_phv_out_data_159; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_160 = pipe3_io_pipe_phv_out_data_160; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_161 = pipe3_io_pipe_phv_out_data_161; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_162 = pipe3_io_pipe_phv_out_data_162; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_163 = pipe3_io_pipe_phv_out_data_163; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_164 = pipe3_io_pipe_phv_out_data_164; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_165 = pipe3_io_pipe_phv_out_data_165; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_166 = pipe3_io_pipe_phv_out_data_166; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_167 = pipe3_io_pipe_phv_out_data_167; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_168 = pipe3_io_pipe_phv_out_data_168; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_169 = pipe3_io_pipe_phv_out_data_169; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_170 = pipe3_io_pipe_phv_out_data_170; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_171 = pipe3_io_pipe_phv_out_data_171; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_172 = pipe3_io_pipe_phv_out_data_172; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_173 = pipe3_io_pipe_phv_out_data_173; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_174 = pipe3_io_pipe_phv_out_data_174; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_175 = pipe3_io_pipe_phv_out_data_175; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_176 = pipe3_io_pipe_phv_out_data_176; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_177 = pipe3_io_pipe_phv_out_data_177; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_178 = pipe3_io_pipe_phv_out_data_178; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_179 = pipe3_io_pipe_phv_out_data_179; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_180 = pipe3_io_pipe_phv_out_data_180; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_181 = pipe3_io_pipe_phv_out_data_181; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_182 = pipe3_io_pipe_phv_out_data_182; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_183 = pipe3_io_pipe_phv_out_data_183; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_184 = pipe3_io_pipe_phv_out_data_184; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_185 = pipe3_io_pipe_phv_out_data_185; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_186 = pipe3_io_pipe_phv_out_data_186; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_187 = pipe3_io_pipe_phv_out_data_187; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_188 = pipe3_io_pipe_phv_out_data_188; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_189 = pipe3_io_pipe_phv_out_data_189; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_190 = pipe3_io_pipe_phv_out_data_190; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_191 = pipe3_io_pipe_phv_out_data_191; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_192 = pipe3_io_pipe_phv_out_data_192; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_193 = pipe3_io_pipe_phv_out_data_193; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_194 = pipe3_io_pipe_phv_out_data_194; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_195 = pipe3_io_pipe_phv_out_data_195; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_196 = pipe3_io_pipe_phv_out_data_196; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_197 = pipe3_io_pipe_phv_out_data_197; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_198 = pipe3_io_pipe_phv_out_data_198; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_199 = pipe3_io_pipe_phv_out_data_199; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_200 = pipe3_io_pipe_phv_out_data_200; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_201 = pipe3_io_pipe_phv_out_data_201; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_202 = pipe3_io_pipe_phv_out_data_202; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_203 = pipe3_io_pipe_phv_out_data_203; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_204 = pipe3_io_pipe_phv_out_data_204; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_205 = pipe3_io_pipe_phv_out_data_205; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_206 = pipe3_io_pipe_phv_out_data_206; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_207 = pipe3_io_pipe_phv_out_data_207; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_208 = pipe3_io_pipe_phv_out_data_208; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_209 = pipe3_io_pipe_phv_out_data_209; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_210 = pipe3_io_pipe_phv_out_data_210; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_211 = pipe3_io_pipe_phv_out_data_211; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_212 = pipe3_io_pipe_phv_out_data_212; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_213 = pipe3_io_pipe_phv_out_data_213; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_214 = pipe3_io_pipe_phv_out_data_214; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_215 = pipe3_io_pipe_phv_out_data_215; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_216 = pipe3_io_pipe_phv_out_data_216; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_217 = pipe3_io_pipe_phv_out_data_217; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_218 = pipe3_io_pipe_phv_out_data_218; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_219 = pipe3_io_pipe_phv_out_data_219; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_220 = pipe3_io_pipe_phv_out_data_220; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_221 = pipe3_io_pipe_phv_out_data_221; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_222 = pipe3_io_pipe_phv_out_data_222; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_223 = pipe3_io_pipe_phv_out_data_223; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_224 = pipe3_io_pipe_phv_out_data_224; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_225 = pipe3_io_pipe_phv_out_data_225; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_226 = pipe3_io_pipe_phv_out_data_226; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_227 = pipe3_io_pipe_phv_out_data_227; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_228 = pipe3_io_pipe_phv_out_data_228; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_229 = pipe3_io_pipe_phv_out_data_229; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_230 = pipe3_io_pipe_phv_out_data_230; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_231 = pipe3_io_pipe_phv_out_data_231; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_232 = pipe3_io_pipe_phv_out_data_232; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_233 = pipe3_io_pipe_phv_out_data_233; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_234 = pipe3_io_pipe_phv_out_data_234; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_235 = pipe3_io_pipe_phv_out_data_235; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_236 = pipe3_io_pipe_phv_out_data_236; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_237 = pipe3_io_pipe_phv_out_data_237; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_238 = pipe3_io_pipe_phv_out_data_238; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_239 = pipe3_io_pipe_phv_out_data_239; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_240 = pipe3_io_pipe_phv_out_data_240; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_241 = pipe3_io_pipe_phv_out_data_241; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_242 = pipe3_io_pipe_phv_out_data_242; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_243 = pipe3_io_pipe_phv_out_data_243; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_244 = pipe3_io_pipe_phv_out_data_244; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_245 = pipe3_io_pipe_phv_out_data_245; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_246 = pipe3_io_pipe_phv_out_data_246; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_247 = pipe3_io_pipe_phv_out_data_247; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_248 = pipe3_io_pipe_phv_out_data_248; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_249 = pipe3_io_pipe_phv_out_data_249; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_250 = pipe3_io_pipe_phv_out_data_250; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_251 = pipe3_io_pipe_phv_out_data_251; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_252 = pipe3_io_pipe_phv_out_data_252; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_253 = pipe3_io_pipe_phv_out_data_253; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_254 = pipe3_io_pipe_phv_out_data_254; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_255 = pipe3_io_pipe_phv_out_data_255; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_256 = pipe3_io_pipe_phv_out_data_256; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_257 = pipe3_io_pipe_phv_out_data_257; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_258 = pipe3_io_pipe_phv_out_data_258; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_259 = pipe3_io_pipe_phv_out_data_259; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_260 = pipe3_io_pipe_phv_out_data_260; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_261 = pipe3_io_pipe_phv_out_data_261; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_262 = pipe3_io_pipe_phv_out_data_262; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_263 = pipe3_io_pipe_phv_out_data_263; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_264 = pipe3_io_pipe_phv_out_data_264; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_265 = pipe3_io_pipe_phv_out_data_265; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_266 = pipe3_io_pipe_phv_out_data_266; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_267 = pipe3_io_pipe_phv_out_data_267; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_268 = pipe3_io_pipe_phv_out_data_268; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_269 = pipe3_io_pipe_phv_out_data_269; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_270 = pipe3_io_pipe_phv_out_data_270; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_271 = pipe3_io_pipe_phv_out_data_271; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_272 = pipe3_io_pipe_phv_out_data_272; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_273 = pipe3_io_pipe_phv_out_data_273; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_274 = pipe3_io_pipe_phv_out_data_274; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_275 = pipe3_io_pipe_phv_out_data_275; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_276 = pipe3_io_pipe_phv_out_data_276; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_277 = pipe3_io_pipe_phv_out_data_277; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_278 = pipe3_io_pipe_phv_out_data_278; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_279 = pipe3_io_pipe_phv_out_data_279; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_280 = pipe3_io_pipe_phv_out_data_280; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_281 = pipe3_io_pipe_phv_out_data_281; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_282 = pipe3_io_pipe_phv_out_data_282; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_283 = pipe3_io_pipe_phv_out_data_283; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_284 = pipe3_io_pipe_phv_out_data_284; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_285 = pipe3_io_pipe_phv_out_data_285; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_286 = pipe3_io_pipe_phv_out_data_286; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_287 = pipe3_io_pipe_phv_out_data_287; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_288 = pipe3_io_pipe_phv_out_data_288; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_289 = pipe3_io_pipe_phv_out_data_289; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_290 = pipe3_io_pipe_phv_out_data_290; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_291 = pipe3_io_pipe_phv_out_data_291; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_292 = pipe3_io_pipe_phv_out_data_292; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_293 = pipe3_io_pipe_phv_out_data_293; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_294 = pipe3_io_pipe_phv_out_data_294; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_295 = pipe3_io_pipe_phv_out_data_295; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_296 = pipe3_io_pipe_phv_out_data_296; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_297 = pipe3_io_pipe_phv_out_data_297; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_298 = pipe3_io_pipe_phv_out_data_298; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_299 = pipe3_io_pipe_phv_out_data_299; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_300 = pipe3_io_pipe_phv_out_data_300; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_301 = pipe3_io_pipe_phv_out_data_301; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_302 = pipe3_io_pipe_phv_out_data_302; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_303 = pipe3_io_pipe_phv_out_data_303; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_304 = pipe3_io_pipe_phv_out_data_304; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_305 = pipe3_io_pipe_phv_out_data_305; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_306 = pipe3_io_pipe_phv_out_data_306; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_307 = pipe3_io_pipe_phv_out_data_307; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_308 = pipe3_io_pipe_phv_out_data_308; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_309 = pipe3_io_pipe_phv_out_data_309; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_310 = pipe3_io_pipe_phv_out_data_310; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_311 = pipe3_io_pipe_phv_out_data_311; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_312 = pipe3_io_pipe_phv_out_data_312; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_313 = pipe3_io_pipe_phv_out_data_313; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_314 = pipe3_io_pipe_phv_out_data_314; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_315 = pipe3_io_pipe_phv_out_data_315; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_316 = pipe3_io_pipe_phv_out_data_316; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_317 = pipe3_io_pipe_phv_out_data_317; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_318 = pipe3_io_pipe_phv_out_data_318; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_319 = pipe3_io_pipe_phv_out_data_319; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_320 = pipe3_io_pipe_phv_out_data_320; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_321 = pipe3_io_pipe_phv_out_data_321; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_322 = pipe3_io_pipe_phv_out_data_322; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_323 = pipe3_io_pipe_phv_out_data_323; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_324 = pipe3_io_pipe_phv_out_data_324; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_325 = pipe3_io_pipe_phv_out_data_325; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_326 = pipe3_io_pipe_phv_out_data_326; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_327 = pipe3_io_pipe_phv_out_data_327; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_328 = pipe3_io_pipe_phv_out_data_328; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_329 = pipe3_io_pipe_phv_out_data_329; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_330 = pipe3_io_pipe_phv_out_data_330; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_331 = pipe3_io_pipe_phv_out_data_331; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_332 = pipe3_io_pipe_phv_out_data_332; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_333 = pipe3_io_pipe_phv_out_data_333; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_334 = pipe3_io_pipe_phv_out_data_334; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_335 = pipe3_io_pipe_phv_out_data_335; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_336 = pipe3_io_pipe_phv_out_data_336; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_337 = pipe3_io_pipe_phv_out_data_337; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_338 = pipe3_io_pipe_phv_out_data_338; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_339 = pipe3_io_pipe_phv_out_data_339; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_340 = pipe3_io_pipe_phv_out_data_340; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_341 = pipe3_io_pipe_phv_out_data_341; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_342 = pipe3_io_pipe_phv_out_data_342; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_343 = pipe3_io_pipe_phv_out_data_343; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_344 = pipe3_io_pipe_phv_out_data_344; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_345 = pipe3_io_pipe_phv_out_data_345; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_346 = pipe3_io_pipe_phv_out_data_346; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_347 = pipe3_io_pipe_phv_out_data_347; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_348 = pipe3_io_pipe_phv_out_data_348; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_349 = pipe3_io_pipe_phv_out_data_349; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_350 = pipe3_io_pipe_phv_out_data_350; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_351 = pipe3_io_pipe_phv_out_data_351; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_352 = pipe3_io_pipe_phv_out_data_352; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_353 = pipe3_io_pipe_phv_out_data_353; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_354 = pipe3_io_pipe_phv_out_data_354; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_355 = pipe3_io_pipe_phv_out_data_355; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_356 = pipe3_io_pipe_phv_out_data_356; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_357 = pipe3_io_pipe_phv_out_data_357; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_358 = pipe3_io_pipe_phv_out_data_358; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_359 = pipe3_io_pipe_phv_out_data_359; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_360 = pipe3_io_pipe_phv_out_data_360; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_361 = pipe3_io_pipe_phv_out_data_361; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_362 = pipe3_io_pipe_phv_out_data_362; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_363 = pipe3_io_pipe_phv_out_data_363; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_364 = pipe3_io_pipe_phv_out_data_364; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_365 = pipe3_io_pipe_phv_out_data_365; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_366 = pipe3_io_pipe_phv_out_data_366; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_367 = pipe3_io_pipe_phv_out_data_367; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_368 = pipe3_io_pipe_phv_out_data_368; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_369 = pipe3_io_pipe_phv_out_data_369; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_370 = pipe3_io_pipe_phv_out_data_370; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_371 = pipe3_io_pipe_phv_out_data_371; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_372 = pipe3_io_pipe_phv_out_data_372; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_373 = pipe3_io_pipe_phv_out_data_373; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_374 = pipe3_io_pipe_phv_out_data_374; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_375 = pipe3_io_pipe_phv_out_data_375; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_376 = pipe3_io_pipe_phv_out_data_376; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_377 = pipe3_io_pipe_phv_out_data_377; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_378 = pipe3_io_pipe_phv_out_data_378; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_379 = pipe3_io_pipe_phv_out_data_379; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_380 = pipe3_io_pipe_phv_out_data_380; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_381 = pipe3_io_pipe_phv_out_data_381; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_382 = pipe3_io_pipe_phv_out_data_382; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_383 = pipe3_io_pipe_phv_out_data_383; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_384 = pipe3_io_pipe_phv_out_data_384; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_385 = pipe3_io_pipe_phv_out_data_385; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_386 = pipe3_io_pipe_phv_out_data_386; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_387 = pipe3_io_pipe_phv_out_data_387; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_388 = pipe3_io_pipe_phv_out_data_388; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_389 = pipe3_io_pipe_phv_out_data_389; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_390 = pipe3_io_pipe_phv_out_data_390; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_391 = pipe3_io_pipe_phv_out_data_391; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_392 = pipe3_io_pipe_phv_out_data_392; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_393 = pipe3_io_pipe_phv_out_data_393; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_394 = pipe3_io_pipe_phv_out_data_394; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_395 = pipe3_io_pipe_phv_out_data_395; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_396 = pipe3_io_pipe_phv_out_data_396; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_397 = pipe3_io_pipe_phv_out_data_397; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_398 = pipe3_io_pipe_phv_out_data_398; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_399 = pipe3_io_pipe_phv_out_data_399; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_400 = pipe3_io_pipe_phv_out_data_400; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_401 = pipe3_io_pipe_phv_out_data_401; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_402 = pipe3_io_pipe_phv_out_data_402; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_403 = pipe3_io_pipe_phv_out_data_403; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_404 = pipe3_io_pipe_phv_out_data_404; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_405 = pipe3_io_pipe_phv_out_data_405; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_406 = pipe3_io_pipe_phv_out_data_406; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_407 = pipe3_io_pipe_phv_out_data_407; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_408 = pipe3_io_pipe_phv_out_data_408; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_409 = pipe3_io_pipe_phv_out_data_409; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_410 = pipe3_io_pipe_phv_out_data_410; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_411 = pipe3_io_pipe_phv_out_data_411; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_412 = pipe3_io_pipe_phv_out_data_412; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_413 = pipe3_io_pipe_phv_out_data_413; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_414 = pipe3_io_pipe_phv_out_data_414; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_415 = pipe3_io_pipe_phv_out_data_415; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_416 = pipe3_io_pipe_phv_out_data_416; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_417 = pipe3_io_pipe_phv_out_data_417; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_418 = pipe3_io_pipe_phv_out_data_418; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_419 = pipe3_io_pipe_phv_out_data_419; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_420 = pipe3_io_pipe_phv_out_data_420; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_421 = pipe3_io_pipe_phv_out_data_421; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_422 = pipe3_io_pipe_phv_out_data_422; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_423 = pipe3_io_pipe_phv_out_data_423; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_424 = pipe3_io_pipe_phv_out_data_424; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_425 = pipe3_io_pipe_phv_out_data_425; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_426 = pipe3_io_pipe_phv_out_data_426; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_427 = pipe3_io_pipe_phv_out_data_427; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_428 = pipe3_io_pipe_phv_out_data_428; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_429 = pipe3_io_pipe_phv_out_data_429; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_430 = pipe3_io_pipe_phv_out_data_430; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_431 = pipe3_io_pipe_phv_out_data_431; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_432 = pipe3_io_pipe_phv_out_data_432; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_433 = pipe3_io_pipe_phv_out_data_433; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_434 = pipe3_io_pipe_phv_out_data_434; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_435 = pipe3_io_pipe_phv_out_data_435; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_436 = pipe3_io_pipe_phv_out_data_436; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_437 = pipe3_io_pipe_phv_out_data_437; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_438 = pipe3_io_pipe_phv_out_data_438; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_439 = pipe3_io_pipe_phv_out_data_439; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_440 = pipe3_io_pipe_phv_out_data_440; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_441 = pipe3_io_pipe_phv_out_data_441; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_442 = pipe3_io_pipe_phv_out_data_442; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_443 = pipe3_io_pipe_phv_out_data_443; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_444 = pipe3_io_pipe_phv_out_data_444; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_445 = pipe3_io_pipe_phv_out_data_445; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_446 = pipe3_io_pipe_phv_out_data_446; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_447 = pipe3_io_pipe_phv_out_data_447; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_448 = pipe3_io_pipe_phv_out_data_448; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_449 = pipe3_io_pipe_phv_out_data_449; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_450 = pipe3_io_pipe_phv_out_data_450; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_451 = pipe3_io_pipe_phv_out_data_451; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_452 = pipe3_io_pipe_phv_out_data_452; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_453 = pipe3_io_pipe_phv_out_data_453; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_454 = pipe3_io_pipe_phv_out_data_454; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_455 = pipe3_io_pipe_phv_out_data_455; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_456 = pipe3_io_pipe_phv_out_data_456; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_457 = pipe3_io_pipe_phv_out_data_457; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_458 = pipe3_io_pipe_phv_out_data_458; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_459 = pipe3_io_pipe_phv_out_data_459; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_460 = pipe3_io_pipe_phv_out_data_460; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_461 = pipe3_io_pipe_phv_out_data_461; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_462 = pipe3_io_pipe_phv_out_data_462; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_463 = pipe3_io_pipe_phv_out_data_463; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_464 = pipe3_io_pipe_phv_out_data_464; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_465 = pipe3_io_pipe_phv_out_data_465; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_466 = pipe3_io_pipe_phv_out_data_466; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_467 = pipe3_io_pipe_phv_out_data_467; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_468 = pipe3_io_pipe_phv_out_data_468; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_469 = pipe3_io_pipe_phv_out_data_469; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_470 = pipe3_io_pipe_phv_out_data_470; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_471 = pipe3_io_pipe_phv_out_data_471; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_472 = pipe3_io_pipe_phv_out_data_472; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_473 = pipe3_io_pipe_phv_out_data_473; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_474 = pipe3_io_pipe_phv_out_data_474; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_475 = pipe3_io_pipe_phv_out_data_475; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_476 = pipe3_io_pipe_phv_out_data_476; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_477 = pipe3_io_pipe_phv_out_data_477; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_478 = pipe3_io_pipe_phv_out_data_478; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_479 = pipe3_io_pipe_phv_out_data_479; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_480 = pipe3_io_pipe_phv_out_data_480; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_481 = pipe3_io_pipe_phv_out_data_481; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_482 = pipe3_io_pipe_phv_out_data_482; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_483 = pipe3_io_pipe_phv_out_data_483; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_484 = pipe3_io_pipe_phv_out_data_484; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_485 = pipe3_io_pipe_phv_out_data_485; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_486 = pipe3_io_pipe_phv_out_data_486; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_487 = pipe3_io_pipe_phv_out_data_487; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_488 = pipe3_io_pipe_phv_out_data_488; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_489 = pipe3_io_pipe_phv_out_data_489; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_490 = pipe3_io_pipe_phv_out_data_490; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_491 = pipe3_io_pipe_phv_out_data_491; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_492 = pipe3_io_pipe_phv_out_data_492; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_493 = pipe3_io_pipe_phv_out_data_493; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_494 = pipe3_io_pipe_phv_out_data_494; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_495 = pipe3_io_pipe_phv_out_data_495; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_496 = pipe3_io_pipe_phv_out_data_496; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_497 = pipe3_io_pipe_phv_out_data_497; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_498 = pipe3_io_pipe_phv_out_data_498; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_499 = pipe3_io_pipe_phv_out_data_499; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_500 = pipe3_io_pipe_phv_out_data_500; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_501 = pipe3_io_pipe_phv_out_data_501; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_502 = pipe3_io_pipe_phv_out_data_502; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_503 = pipe3_io_pipe_phv_out_data_503; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_504 = pipe3_io_pipe_phv_out_data_504; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_505 = pipe3_io_pipe_phv_out_data_505; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_506 = pipe3_io_pipe_phv_out_data_506; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_507 = pipe3_io_pipe_phv_out_data_507; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_508 = pipe3_io_pipe_phv_out_data_508; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_509 = pipe3_io_pipe_phv_out_data_509; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_510 = pipe3_io_pipe_phv_out_data_510; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_data_511 = pipe3_io_pipe_phv_out_data_511; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_next_processor_id = pipe3_io_pipe_phv_out_next_processor_id; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_next_config_id = pipe3_io_pipe_phv_out_next_config_id; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_pipe_phv_in_is_valid_processor = pipe3_io_pipe_phv_out_is_valid_processor; // @[matcher_pisa.scala 354:26]
  assign pipe4_io_key_config_0_field_config_0 = key_config_0_field_config_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_config_1 = key_config_0_field_config_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_config_2 = key_config_0_field_config_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_config_3 = key_config_0_field_config_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_config_4 = key_config_0_field_config_4; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_config_5 = key_config_0_field_config_5; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_0_0 = key_config_0_field_mask_0_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_0_1 = key_config_0_field_mask_0_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_0_2 = key_config_0_field_mask_0_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_0_3 = key_config_0_field_mask_0_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_1_0 = key_config_0_field_mask_1_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_1_1 = key_config_0_field_mask_1_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_1_2 = key_config_0_field_mask_1_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_1_3 = key_config_0_field_mask_1_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_2_0 = key_config_0_field_mask_2_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_2_1 = key_config_0_field_mask_2_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_2_2 = key_config_0_field_mask_2_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_2_3 = key_config_0_field_mask_2_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_3_0 = key_config_0_field_mask_3_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_3_1 = key_config_0_field_mask_3_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_3_2 = key_config_0_field_mask_3_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_3_3 = key_config_0_field_mask_3_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_4_0 = key_config_0_field_mask_4_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_4_1 = key_config_0_field_mask_4_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_4_2 = key_config_0_field_mask_4_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_4_3 = key_config_0_field_mask_4_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_5_0 = key_config_0_field_mask_5_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_5_1 = key_config_0_field_mask_5_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_5_2 = key_config_0_field_mask_5_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_0_field_mask_5_3 = key_config_0_field_mask_5_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_config_0 = key_config_1_field_config_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_config_1 = key_config_1_field_config_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_config_2 = key_config_1_field_config_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_config_3 = key_config_1_field_config_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_config_4 = key_config_1_field_config_4; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_config_5 = key_config_1_field_config_5; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_0_0 = key_config_1_field_mask_0_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_0_1 = key_config_1_field_mask_0_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_0_2 = key_config_1_field_mask_0_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_0_3 = key_config_1_field_mask_0_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_1_0 = key_config_1_field_mask_1_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_1_1 = key_config_1_field_mask_1_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_1_2 = key_config_1_field_mask_1_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_1_3 = key_config_1_field_mask_1_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_2_0 = key_config_1_field_mask_2_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_2_1 = key_config_1_field_mask_2_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_2_2 = key_config_1_field_mask_2_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_2_3 = key_config_1_field_mask_2_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_3_0 = key_config_1_field_mask_3_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_3_1 = key_config_1_field_mask_3_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_3_2 = key_config_1_field_mask_3_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_3_3 = key_config_1_field_mask_3_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_4_0 = key_config_1_field_mask_4_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_4_1 = key_config_1_field_mask_4_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_4_2 = key_config_1_field_mask_4_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_4_3 = key_config_1_field_mask_4_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_5_0 = key_config_1_field_mask_5_0; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_5_1 = key_config_1_field_mask_5_1; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_5_2 = key_config_1_field_mask_5_2; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_config_1_field_mask_5_3 = key_config_1_field_mask_5_3; // @[matcher_pisa.scala 357:26]
  assign pipe4_io_key_in = pipe3_io_key_out; // @[matcher_pisa.scala 355:26]
  assign pipe4_io_data_in = pipe3_io_data_out; // @[matcher_pisa.scala 356:26]
  always @(posedge clock) begin
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (~io_mod_config_id & 3'h0 == io_mod_key_mod_group_index) begin // @[matcher_pisa.scala 74:83]
          key_config_0_field_config_0 <= io_mod_key_mod_group_config; // @[matcher_pisa.scala 74:83]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (~io_mod_config_id & 3'h1 == io_mod_key_mod_group_index) begin // @[matcher_pisa.scala 74:83]
          key_config_0_field_config_1 <= io_mod_key_mod_group_config; // @[matcher_pisa.scala 74:83]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (~io_mod_config_id & 3'h2 == io_mod_key_mod_group_index) begin // @[matcher_pisa.scala 74:83]
          key_config_0_field_config_2 <= io_mod_key_mod_group_config; // @[matcher_pisa.scala 74:83]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (~io_mod_config_id & 3'h3 == io_mod_key_mod_group_index) begin // @[matcher_pisa.scala 74:83]
          key_config_0_field_config_3 <= io_mod_key_mod_group_config; // @[matcher_pisa.scala 74:83]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (~io_mod_config_id & 3'h4 == io_mod_key_mod_group_index) begin // @[matcher_pisa.scala 74:83]
          key_config_0_field_config_4 <= io_mod_key_mod_group_config; // @[matcher_pisa.scala 74:83]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (~io_mod_config_id & 3'h5 == io_mod_key_mod_group_index) begin // @[matcher_pisa.scala 74:83]
          key_config_0_field_config_5 <= io_mod_key_mod_group_config; // @[matcher_pisa.scala 74:83]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_339) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_0_0 <= io_mod_key_mod_group_mask_0; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_339) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_0_1 <= io_mod_key_mod_group_mask_1; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_339) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_0_2 <= io_mod_key_mod_group_mask_2; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_339) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_0_3 <= io_mod_key_mod_group_mask_3; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_341) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_1_0 <= io_mod_key_mod_group_mask_0; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_341) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_1_1 <= io_mod_key_mod_group_mask_1; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_341) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_1_2 <= io_mod_key_mod_group_mask_2; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_341) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_1_3 <= io_mod_key_mod_group_mask_3; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_343) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_2_0 <= io_mod_key_mod_group_mask_0; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_343) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_2_1 <= io_mod_key_mod_group_mask_1; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_343) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_2_2 <= io_mod_key_mod_group_mask_2; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_343) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_2_3 <= io_mod_key_mod_group_mask_3; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_345) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_3_0 <= io_mod_key_mod_group_mask_0; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_345) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_3_1 <= io_mod_key_mod_group_mask_1; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_345) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_3_2 <= io_mod_key_mod_group_mask_2; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_345) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_3_3 <= io_mod_key_mod_group_mask_3; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_347) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_4_0 <= io_mod_key_mod_group_mask_0; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_347) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_4_1 <= io_mod_key_mod_group_mask_1; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_347) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_4_2 <= io_mod_key_mod_group_mask_2; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_347) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_4_3 <= io_mod_key_mod_group_mask_3; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_349) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_5_0 <= io_mod_key_mod_group_mask_0; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_349) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_5_1 <= io_mod_key_mod_group_mask_1; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_349) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_5_2 <= io_mod_key_mod_group_mask_2; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_349) begin // @[matcher_pisa.scala 76:81]
          key_config_0_field_mask_5_3 <= io_mod_key_mod_group_mask_3; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_339) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_0_0 <= io_mod_key_mod_group_id_0; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_339) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_0_1 <= io_mod_key_mod_group_id_1; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_339) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_0_2 <= io_mod_key_mod_group_id_2; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_339) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_0_3 <= io_mod_key_mod_group_id_3; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_341) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_1_0 <= io_mod_key_mod_group_id_0; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_341) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_1_1 <= io_mod_key_mod_group_id_1; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_341) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_1_2 <= io_mod_key_mod_group_id_2; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_341) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_1_3 <= io_mod_key_mod_group_id_3; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_343) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_2_0 <= io_mod_key_mod_group_id_0; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_343) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_2_1 <= io_mod_key_mod_group_id_1; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_343) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_2_2 <= io_mod_key_mod_group_id_2; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_343) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_2_3 <= io_mod_key_mod_group_id_3; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_345) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_3_0 <= io_mod_key_mod_group_id_0; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_345) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_3_1 <= io_mod_key_mod_group_id_1; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_345) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_3_2 <= io_mod_key_mod_group_id_2; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_345) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_3_3 <= io_mod_key_mod_group_id_3; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_347) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_4_0 <= io_mod_key_mod_group_id_0; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_347) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_4_1 <= io_mod_key_mod_group_id_1; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_347) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_4_2 <= io_mod_key_mod_group_id_2; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_347) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_4_3 <= io_mod_key_mod_group_id_3; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_349) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_5_0 <= io_mod_key_mod_group_id_0; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_349) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_5_1 <= io_mod_key_mod_group_id_1; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_349) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_5_2 <= io_mod_key_mod_group_id_2; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (_GEN_338 & _GEN_349) begin // @[matcher_pisa.scala 75:79]
          key_config_0_field_id_5_3 <= io_mod_key_mod_group_id_3; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & 3'h0 == io_mod_key_mod_group_index) begin // @[matcher_pisa.scala 74:83]
          key_config_1_field_config_0 <= io_mod_key_mod_group_config; // @[matcher_pisa.scala 74:83]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & 3'h1 == io_mod_key_mod_group_index) begin // @[matcher_pisa.scala 74:83]
          key_config_1_field_config_1 <= io_mod_key_mod_group_config; // @[matcher_pisa.scala 74:83]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & 3'h2 == io_mod_key_mod_group_index) begin // @[matcher_pisa.scala 74:83]
          key_config_1_field_config_2 <= io_mod_key_mod_group_config; // @[matcher_pisa.scala 74:83]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & 3'h3 == io_mod_key_mod_group_index) begin // @[matcher_pisa.scala 74:83]
          key_config_1_field_config_3 <= io_mod_key_mod_group_config; // @[matcher_pisa.scala 74:83]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & 3'h4 == io_mod_key_mod_group_index) begin // @[matcher_pisa.scala 74:83]
          key_config_1_field_config_4 <= io_mod_key_mod_group_config; // @[matcher_pisa.scala 74:83]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & 3'h5 == io_mod_key_mod_group_index) begin // @[matcher_pisa.scala 74:83]
          key_config_1_field_config_5 <= io_mod_key_mod_group_config; // @[matcher_pisa.scala 74:83]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_339) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_0_0 <= io_mod_key_mod_group_mask_0; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_339) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_0_1 <= io_mod_key_mod_group_mask_1; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_339) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_0_2 <= io_mod_key_mod_group_mask_2; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_339) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_0_3 <= io_mod_key_mod_group_mask_3; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_341) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_1_0 <= io_mod_key_mod_group_mask_0; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_341) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_1_1 <= io_mod_key_mod_group_mask_1; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_341) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_1_2 <= io_mod_key_mod_group_mask_2; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_341) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_1_3 <= io_mod_key_mod_group_mask_3; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_343) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_2_0 <= io_mod_key_mod_group_mask_0; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_343) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_2_1 <= io_mod_key_mod_group_mask_1; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_343) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_2_2 <= io_mod_key_mod_group_mask_2; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_343) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_2_3 <= io_mod_key_mod_group_mask_3; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_345) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_3_0 <= io_mod_key_mod_group_mask_0; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_345) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_3_1 <= io_mod_key_mod_group_mask_1; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_345) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_3_2 <= io_mod_key_mod_group_mask_2; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_345) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_3_3 <= io_mod_key_mod_group_mask_3; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_347) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_4_0 <= io_mod_key_mod_group_mask_0; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_347) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_4_1 <= io_mod_key_mod_group_mask_1; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_347) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_4_2 <= io_mod_key_mod_group_mask_2; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_347) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_4_3 <= io_mod_key_mod_group_mask_3; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_349) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_5_0 <= io_mod_key_mod_group_mask_0; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_349) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_5_1 <= io_mod_key_mod_group_mask_1; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_349) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_5_2 <= io_mod_key_mod_group_mask_2; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_349) begin // @[matcher_pisa.scala 76:81]
          key_config_1_field_mask_5_3 <= io_mod_key_mod_group_mask_3; // @[matcher_pisa.scala 76:81]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_339) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_0_0 <= io_mod_key_mod_group_id_0; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_339) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_0_1 <= io_mod_key_mod_group_id_1; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_339) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_0_2 <= io_mod_key_mod_group_id_2; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_339) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_0_3 <= io_mod_key_mod_group_id_3; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_341) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_1_0 <= io_mod_key_mod_group_id_0; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_341) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_1_1 <= io_mod_key_mod_group_id_1; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_341) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_1_2 <= io_mod_key_mod_group_id_2; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_341) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_1_3 <= io_mod_key_mod_group_id_3; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_343) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_2_0 <= io_mod_key_mod_group_id_0; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_343) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_2_1 <= io_mod_key_mod_group_id_1; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_343) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_2_2 <= io_mod_key_mod_group_id_2; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_343) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_2_3 <= io_mod_key_mod_group_id_3; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_345) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_3_0 <= io_mod_key_mod_group_id_0; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_345) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_3_1 <= io_mod_key_mod_group_id_1; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_345) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_3_2 <= io_mod_key_mod_group_id_2; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_345) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_3_3 <= io_mod_key_mod_group_id_3; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_347) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_4_0 <= io_mod_key_mod_group_id_0; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_347) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_4_1 <= io_mod_key_mod_group_id_1; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_347) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_4_2 <= io_mod_key_mod_group_id_2; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_347) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_4_3 <= io_mod_key_mod_group_id_3; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_349) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_5_0 <= io_mod_key_mod_group_id_0; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_349) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_5_1 <= io_mod_key_mod_group_id_1; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_349) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_5_2 <= io_mod_key_mod_group_id_2; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_key_mod_en) begin // @[matcher_pisa.scala 73:34]
        if (io_mod_config_id & _GEN_349) begin // @[matcher_pisa.scala 75:79]
          key_config_1_field_id_5_3 <= io_mod_key_mod_group_id_3; // @[matcher_pisa.scala 75:79]
        end
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (~io_mod_config_id) begin // @[matcher_pisa.scala 79:40]
        table_config_0_table_depth <= io_mod_table_mod_table_depth; // @[matcher_pisa.scala 79:40]
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (~io_mod_config_id) begin // @[matcher_pisa.scala 79:40]
        table_config_0_table_width <= io_mod_table_mod_table_width; // @[matcher_pisa.scala 79:40]
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_config_id) begin // @[matcher_pisa.scala 79:40]
        table_config_1_table_depth <= io_mod_table_mod_table_depth; // @[matcher_pisa.scala 79:40]
      end
    end
    if (io_mod_en) begin // @[matcher_pisa.scala 72:22]
      if (io_mod_config_id) begin // @[matcher_pisa.scala 79:40]
        table_config_1_table_width <= io_mod_table_mod_table_width; // @[matcher_pisa.scala 79:40]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  key_config_0_field_config_0 = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  key_config_0_field_config_1 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  key_config_0_field_config_2 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  key_config_0_field_config_3 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  key_config_0_field_config_4 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  key_config_0_field_config_5 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  key_config_0_field_mask_0_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  key_config_0_field_mask_0_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  key_config_0_field_mask_0_2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  key_config_0_field_mask_0_3 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  key_config_0_field_mask_1_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  key_config_0_field_mask_1_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  key_config_0_field_mask_1_2 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  key_config_0_field_mask_1_3 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  key_config_0_field_mask_2_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  key_config_0_field_mask_2_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  key_config_0_field_mask_2_2 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  key_config_0_field_mask_2_3 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  key_config_0_field_mask_3_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  key_config_0_field_mask_3_1 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  key_config_0_field_mask_3_2 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  key_config_0_field_mask_3_3 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  key_config_0_field_mask_4_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  key_config_0_field_mask_4_1 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  key_config_0_field_mask_4_2 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  key_config_0_field_mask_4_3 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  key_config_0_field_mask_5_0 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  key_config_0_field_mask_5_1 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  key_config_0_field_mask_5_2 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  key_config_0_field_mask_5_3 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  key_config_0_field_id_0_0 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  key_config_0_field_id_0_1 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  key_config_0_field_id_0_2 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  key_config_0_field_id_0_3 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  key_config_0_field_id_1_0 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  key_config_0_field_id_1_1 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  key_config_0_field_id_1_2 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  key_config_0_field_id_1_3 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  key_config_0_field_id_2_0 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  key_config_0_field_id_2_1 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  key_config_0_field_id_2_2 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  key_config_0_field_id_2_3 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  key_config_0_field_id_3_0 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  key_config_0_field_id_3_1 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  key_config_0_field_id_3_2 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  key_config_0_field_id_3_3 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  key_config_0_field_id_4_0 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  key_config_0_field_id_4_1 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  key_config_0_field_id_4_2 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  key_config_0_field_id_4_3 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  key_config_0_field_id_5_0 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  key_config_0_field_id_5_1 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  key_config_0_field_id_5_2 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  key_config_0_field_id_5_3 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  key_config_1_field_config_0 = _RAND_54[1:0];
  _RAND_55 = {1{`RANDOM}};
  key_config_1_field_config_1 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  key_config_1_field_config_2 = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  key_config_1_field_config_3 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  key_config_1_field_config_4 = _RAND_58[1:0];
  _RAND_59 = {1{`RANDOM}};
  key_config_1_field_config_5 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  key_config_1_field_mask_0_0 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  key_config_1_field_mask_0_1 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  key_config_1_field_mask_0_2 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  key_config_1_field_mask_0_3 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  key_config_1_field_mask_1_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  key_config_1_field_mask_1_1 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  key_config_1_field_mask_1_2 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  key_config_1_field_mask_1_3 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  key_config_1_field_mask_2_0 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  key_config_1_field_mask_2_1 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  key_config_1_field_mask_2_2 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  key_config_1_field_mask_2_3 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  key_config_1_field_mask_3_0 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  key_config_1_field_mask_3_1 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  key_config_1_field_mask_3_2 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  key_config_1_field_mask_3_3 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  key_config_1_field_mask_4_0 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  key_config_1_field_mask_4_1 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  key_config_1_field_mask_4_2 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  key_config_1_field_mask_4_3 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  key_config_1_field_mask_5_0 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  key_config_1_field_mask_5_1 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  key_config_1_field_mask_5_2 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  key_config_1_field_mask_5_3 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  key_config_1_field_id_0_0 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  key_config_1_field_id_0_1 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  key_config_1_field_id_0_2 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  key_config_1_field_id_0_3 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  key_config_1_field_id_1_0 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  key_config_1_field_id_1_1 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  key_config_1_field_id_1_2 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  key_config_1_field_id_1_3 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  key_config_1_field_id_2_0 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  key_config_1_field_id_2_1 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  key_config_1_field_id_2_2 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  key_config_1_field_id_2_3 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  key_config_1_field_id_3_0 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  key_config_1_field_id_3_1 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  key_config_1_field_id_3_2 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  key_config_1_field_id_3_3 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  key_config_1_field_id_4_0 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  key_config_1_field_id_4_1 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  key_config_1_field_id_4_2 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  key_config_1_field_id_4_3 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  key_config_1_field_id_5_0 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  key_config_1_field_id_5_1 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  key_config_1_field_id_5_2 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  key_config_1_field_id_5_3 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  table_config_0_table_depth = _RAND_108[4:0];
  _RAND_109 = {1{`RANDOM}};
  table_config_0_table_width = _RAND_109[4:0];
  _RAND_110 = {1{`RANDOM}};
  table_config_1_table_depth = _RAND_110[4:0];
  _RAND_111 = {1{`RANDOM}};
  table_config_1_table_width = _RAND_111[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
