module MatchResult(
  input          clock,
  input  [7:0]   io_pipe_phv_in_data_0,
  input  [7:0]   io_pipe_phv_in_data_1,
  input  [7:0]   io_pipe_phv_in_data_2,
  input  [7:0]   io_pipe_phv_in_data_3,
  input  [7:0]   io_pipe_phv_in_data_4,
  input  [7:0]   io_pipe_phv_in_data_5,
  input  [7:0]   io_pipe_phv_in_data_6,
  input  [7:0]   io_pipe_phv_in_data_7,
  input  [7:0]   io_pipe_phv_in_data_8,
  input  [7:0]   io_pipe_phv_in_data_9,
  input  [7:0]   io_pipe_phv_in_data_10,
  input  [7:0]   io_pipe_phv_in_data_11,
  input  [7:0]   io_pipe_phv_in_data_12,
  input  [7:0]   io_pipe_phv_in_data_13,
  input  [7:0]   io_pipe_phv_in_data_14,
  input  [7:0]   io_pipe_phv_in_data_15,
  input  [7:0]   io_pipe_phv_in_data_16,
  input  [7:0]   io_pipe_phv_in_data_17,
  input  [7:0]   io_pipe_phv_in_data_18,
  input  [7:0]   io_pipe_phv_in_data_19,
  input  [7:0]   io_pipe_phv_in_data_20,
  input  [7:0]   io_pipe_phv_in_data_21,
  input  [7:0]   io_pipe_phv_in_data_22,
  input  [7:0]   io_pipe_phv_in_data_23,
  input  [7:0]   io_pipe_phv_in_data_24,
  input  [7:0]   io_pipe_phv_in_data_25,
  input  [7:0]   io_pipe_phv_in_data_26,
  input  [7:0]   io_pipe_phv_in_data_27,
  input  [7:0]   io_pipe_phv_in_data_28,
  input  [7:0]   io_pipe_phv_in_data_29,
  input  [7:0]   io_pipe_phv_in_data_30,
  input  [7:0]   io_pipe_phv_in_data_31,
  input  [7:0]   io_pipe_phv_in_data_32,
  input  [7:0]   io_pipe_phv_in_data_33,
  input  [7:0]   io_pipe_phv_in_data_34,
  input  [7:0]   io_pipe_phv_in_data_35,
  input  [7:0]   io_pipe_phv_in_data_36,
  input  [7:0]   io_pipe_phv_in_data_37,
  input  [7:0]   io_pipe_phv_in_data_38,
  input  [7:0]   io_pipe_phv_in_data_39,
  input  [7:0]   io_pipe_phv_in_data_40,
  input  [7:0]   io_pipe_phv_in_data_41,
  input  [7:0]   io_pipe_phv_in_data_42,
  input  [7:0]   io_pipe_phv_in_data_43,
  input  [7:0]   io_pipe_phv_in_data_44,
  input  [7:0]   io_pipe_phv_in_data_45,
  input  [7:0]   io_pipe_phv_in_data_46,
  input  [7:0]   io_pipe_phv_in_data_47,
  input  [7:0]   io_pipe_phv_in_data_48,
  input  [7:0]   io_pipe_phv_in_data_49,
  input  [7:0]   io_pipe_phv_in_data_50,
  input  [7:0]   io_pipe_phv_in_data_51,
  input  [7:0]   io_pipe_phv_in_data_52,
  input  [7:0]   io_pipe_phv_in_data_53,
  input  [7:0]   io_pipe_phv_in_data_54,
  input  [7:0]   io_pipe_phv_in_data_55,
  input  [7:0]   io_pipe_phv_in_data_56,
  input  [7:0]   io_pipe_phv_in_data_57,
  input  [7:0]   io_pipe_phv_in_data_58,
  input  [7:0]   io_pipe_phv_in_data_59,
  input  [7:0]   io_pipe_phv_in_data_60,
  input  [7:0]   io_pipe_phv_in_data_61,
  input  [7:0]   io_pipe_phv_in_data_62,
  input  [7:0]   io_pipe_phv_in_data_63,
  input  [7:0]   io_pipe_phv_in_data_64,
  input  [7:0]   io_pipe_phv_in_data_65,
  input  [7:0]   io_pipe_phv_in_data_66,
  input  [7:0]   io_pipe_phv_in_data_67,
  input  [7:0]   io_pipe_phv_in_data_68,
  input  [7:0]   io_pipe_phv_in_data_69,
  input  [7:0]   io_pipe_phv_in_data_70,
  input  [7:0]   io_pipe_phv_in_data_71,
  input  [7:0]   io_pipe_phv_in_data_72,
  input  [7:0]   io_pipe_phv_in_data_73,
  input  [7:0]   io_pipe_phv_in_data_74,
  input  [7:0]   io_pipe_phv_in_data_75,
  input  [7:0]   io_pipe_phv_in_data_76,
  input  [7:0]   io_pipe_phv_in_data_77,
  input  [7:0]   io_pipe_phv_in_data_78,
  input  [7:0]   io_pipe_phv_in_data_79,
  input  [7:0]   io_pipe_phv_in_data_80,
  input  [7:0]   io_pipe_phv_in_data_81,
  input  [7:0]   io_pipe_phv_in_data_82,
  input  [7:0]   io_pipe_phv_in_data_83,
  input  [7:0]   io_pipe_phv_in_data_84,
  input  [7:0]   io_pipe_phv_in_data_85,
  input  [7:0]   io_pipe_phv_in_data_86,
  input  [7:0]   io_pipe_phv_in_data_87,
  input  [7:0]   io_pipe_phv_in_data_88,
  input  [7:0]   io_pipe_phv_in_data_89,
  input  [7:0]   io_pipe_phv_in_data_90,
  input  [7:0]   io_pipe_phv_in_data_91,
  input  [7:0]   io_pipe_phv_in_data_92,
  input  [7:0]   io_pipe_phv_in_data_93,
  input  [7:0]   io_pipe_phv_in_data_94,
  input  [7:0]   io_pipe_phv_in_data_95,
  input  [7:0]   io_pipe_phv_in_data_96,
  input  [7:0]   io_pipe_phv_in_data_97,
  input  [7:0]   io_pipe_phv_in_data_98,
  input  [7:0]   io_pipe_phv_in_data_99,
  input  [7:0]   io_pipe_phv_in_data_100,
  input  [7:0]   io_pipe_phv_in_data_101,
  input  [7:0]   io_pipe_phv_in_data_102,
  input  [7:0]   io_pipe_phv_in_data_103,
  input  [7:0]   io_pipe_phv_in_data_104,
  input  [7:0]   io_pipe_phv_in_data_105,
  input  [7:0]   io_pipe_phv_in_data_106,
  input  [7:0]   io_pipe_phv_in_data_107,
  input  [7:0]   io_pipe_phv_in_data_108,
  input  [7:0]   io_pipe_phv_in_data_109,
  input  [7:0]   io_pipe_phv_in_data_110,
  input  [7:0]   io_pipe_phv_in_data_111,
  input  [7:0]   io_pipe_phv_in_data_112,
  input  [7:0]   io_pipe_phv_in_data_113,
  input  [7:0]   io_pipe_phv_in_data_114,
  input  [7:0]   io_pipe_phv_in_data_115,
  input  [7:0]   io_pipe_phv_in_data_116,
  input  [7:0]   io_pipe_phv_in_data_117,
  input  [7:0]   io_pipe_phv_in_data_118,
  input  [7:0]   io_pipe_phv_in_data_119,
  input  [7:0]   io_pipe_phv_in_data_120,
  input  [7:0]   io_pipe_phv_in_data_121,
  input  [7:0]   io_pipe_phv_in_data_122,
  input  [7:0]   io_pipe_phv_in_data_123,
  input  [7:0]   io_pipe_phv_in_data_124,
  input  [7:0]   io_pipe_phv_in_data_125,
  input  [7:0]   io_pipe_phv_in_data_126,
  input  [7:0]   io_pipe_phv_in_data_127,
  input  [7:0]   io_pipe_phv_in_data_128,
  input  [7:0]   io_pipe_phv_in_data_129,
  input  [7:0]   io_pipe_phv_in_data_130,
  input  [7:0]   io_pipe_phv_in_data_131,
  input  [7:0]   io_pipe_phv_in_data_132,
  input  [7:0]   io_pipe_phv_in_data_133,
  input  [7:0]   io_pipe_phv_in_data_134,
  input  [7:0]   io_pipe_phv_in_data_135,
  input  [7:0]   io_pipe_phv_in_data_136,
  input  [7:0]   io_pipe_phv_in_data_137,
  input  [7:0]   io_pipe_phv_in_data_138,
  input  [7:0]   io_pipe_phv_in_data_139,
  input  [7:0]   io_pipe_phv_in_data_140,
  input  [7:0]   io_pipe_phv_in_data_141,
  input  [7:0]   io_pipe_phv_in_data_142,
  input  [7:0]   io_pipe_phv_in_data_143,
  input  [7:0]   io_pipe_phv_in_data_144,
  input  [7:0]   io_pipe_phv_in_data_145,
  input  [7:0]   io_pipe_phv_in_data_146,
  input  [7:0]   io_pipe_phv_in_data_147,
  input  [7:0]   io_pipe_phv_in_data_148,
  input  [7:0]   io_pipe_phv_in_data_149,
  input  [7:0]   io_pipe_phv_in_data_150,
  input  [7:0]   io_pipe_phv_in_data_151,
  input  [7:0]   io_pipe_phv_in_data_152,
  input  [7:0]   io_pipe_phv_in_data_153,
  input  [7:0]   io_pipe_phv_in_data_154,
  input  [7:0]   io_pipe_phv_in_data_155,
  input  [7:0]   io_pipe_phv_in_data_156,
  input  [7:0]   io_pipe_phv_in_data_157,
  input  [7:0]   io_pipe_phv_in_data_158,
  input  [7:0]   io_pipe_phv_in_data_159,
  input  [7:0]   io_pipe_phv_in_data_160,
  input  [7:0]   io_pipe_phv_in_data_161,
  input  [7:0]   io_pipe_phv_in_data_162,
  input  [7:0]   io_pipe_phv_in_data_163,
  input  [7:0]   io_pipe_phv_in_data_164,
  input  [7:0]   io_pipe_phv_in_data_165,
  input  [7:0]   io_pipe_phv_in_data_166,
  input  [7:0]   io_pipe_phv_in_data_167,
  input  [7:0]   io_pipe_phv_in_data_168,
  input  [7:0]   io_pipe_phv_in_data_169,
  input  [7:0]   io_pipe_phv_in_data_170,
  input  [7:0]   io_pipe_phv_in_data_171,
  input  [7:0]   io_pipe_phv_in_data_172,
  input  [7:0]   io_pipe_phv_in_data_173,
  input  [7:0]   io_pipe_phv_in_data_174,
  input  [7:0]   io_pipe_phv_in_data_175,
  input  [7:0]   io_pipe_phv_in_data_176,
  input  [7:0]   io_pipe_phv_in_data_177,
  input  [7:0]   io_pipe_phv_in_data_178,
  input  [7:0]   io_pipe_phv_in_data_179,
  input  [7:0]   io_pipe_phv_in_data_180,
  input  [7:0]   io_pipe_phv_in_data_181,
  input  [7:0]   io_pipe_phv_in_data_182,
  input  [7:0]   io_pipe_phv_in_data_183,
  input  [7:0]   io_pipe_phv_in_data_184,
  input  [7:0]   io_pipe_phv_in_data_185,
  input  [7:0]   io_pipe_phv_in_data_186,
  input  [7:0]   io_pipe_phv_in_data_187,
  input  [7:0]   io_pipe_phv_in_data_188,
  input  [7:0]   io_pipe_phv_in_data_189,
  input  [7:0]   io_pipe_phv_in_data_190,
  input  [7:0]   io_pipe_phv_in_data_191,
  input  [7:0]   io_pipe_phv_in_data_192,
  input  [7:0]   io_pipe_phv_in_data_193,
  input  [7:0]   io_pipe_phv_in_data_194,
  input  [7:0]   io_pipe_phv_in_data_195,
  input  [7:0]   io_pipe_phv_in_data_196,
  input  [7:0]   io_pipe_phv_in_data_197,
  input  [7:0]   io_pipe_phv_in_data_198,
  input  [7:0]   io_pipe_phv_in_data_199,
  input  [7:0]   io_pipe_phv_in_data_200,
  input  [7:0]   io_pipe_phv_in_data_201,
  input  [7:0]   io_pipe_phv_in_data_202,
  input  [7:0]   io_pipe_phv_in_data_203,
  input  [7:0]   io_pipe_phv_in_data_204,
  input  [7:0]   io_pipe_phv_in_data_205,
  input  [7:0]   io_pipe_phv_in_data_206,
  input  [7:0]   io_pipe_phv_in_data_207,
  input  [7:0]   io_pipe_phv_in_data_208,
  input  [7:0]   io_pipe_phv_in_data_209,
  input  [7:0]   io_pipe_phv_in_data_210,
  input  [7:0]   io_pipe_phv_in_data_211,
  input  [7:0]   io_pipe_phv_in_data_212,
  input  [7:0]   io_pipe_phv_in_data_213,
  input  [7:0]   io_pipe_phv_in_data_214,
  input  [7:0]   io_pipe_phv_in_data_215,
  input  [7:0]   io_pipe_phv_in_data_216,
  input  [7:0]   io_pipe_phv_in_data_217,
  input  [7:0]   io_pipe_phv_in_data_218,
  input  [7:0]   io_pipe_phv_in_data_219,
  input  [7:0]   io_pipe_phv_in_data_220,
  input  [7:0]   io_pipe_phv_in_data_221,
  input  [7:0]   io_pipe_phv_in_data_222,
  input  [7:0]   io_pipe_phv_in_data_223,
  input  [7:0]   io_pipe_phv_in_data_224,
  input  [7:0]   io_pipe_phv_in_data_225,
  input  [7:0]   io_pipe_phv_in_data_226,
  input  [7:0]   io_pipe_phv_in_data_227,
  input  [7:0]   io_pipe_phv_in_data_228,
  input  [7:0]   io_pipe_phv_in_data_229,
  input  [7:0]   io_pipe_phv_in_data_230,
  input  [7:0]   io_pipe_phv_in_data_231,
  input  [7:0]   io_pipe_phv_in_data_232,
  input  [7:0]   io_pipe_phv_in_data_233,
  input  [7:0]   io_pipe_phv_in_data_234,
  input  [7:0]   io_pipe_phv_in_data_235,
  input  [7:0]   io_pipe_phv_in_data_236,
  input  [7:0]   io_pipe_phv_in_data_237,
  input  [7:0]   io_pipe_phv_in_data_238,
  input  [7:0]   io_pipe_phv_in_data_239,
  input  [7:0]   io_pipe_phv_in_data_240,
  input  [7:0]   io_pipe_phv_in_data_241,
  input  [7:0]   io_pipe_phv_in_data_242,
  input  [7:0]   io_pipe_phv_in_data_243,
  input  [7:0]   io_pipe_phv_in_data_244,
  input  [7:0]   io_pipe_phv_in_data_245,
  input  [7:0]   io_pipe_phv_in_data_246,
  input  [7:0]   io_pipe_phv_in_data_247,
  input  [7:0]   io_pipe_phv_in_data_248,
  input  [7:0]   io_pipe_phv_in_data_249,
  input  [7:0]   io_pipe_phv_in_data_250,
  input  [7:0]   io_pipe_phv_in_data_251,
  input  [7:0]   io_pipe_phv_in_data_252,
  input  [7:0]   io_pipe_phv_in_data_253,
  input  [7:0]   io_pipe_phv_in_data_254,
  input  [7:0]   io_pipe_phv_in_data_255,
  input  [15:0]  io_pipe_phv_in_header_0,
  input  [15:0]  io_pipe_phv_in_header_1,
  input  [15:0]  io_pipe_phv_in_header_2,
  input  [15:0]  io_pipe_phv_in_header_3,
  input  [15:0]  io_pipe_phv_in_header_4,
  input  [15:0]  io_pipe_phv_in_header_5,
  input  [15:0]  io_pipe_phv_in_header_6,
  input  [15:0]  io_pipe_phv_in_header_7,
  input  [15:0]  io_pipe_phv_in_header_8,
  input  [15:0]  io_pipe_phv_in_header_9,
  input  [15:0]  io_pipe_phv_in_header_10,
  input  [15:0]  io_pipe_phv_in_header_11,
  input  [15:0]  io_pipe_phv_in_header_12,
  input  [15:0]  io_pipe_phv_in_header_13,
  input  [15:0]  io_pipe_phv_in_header_14,
  input  [15:0]  io_pipe_phv_in_header_15,
  input  [7:0]   io_pipe_phv_in_parse_current_state,
  input  [7:0]   io_pipe_phv_in_parse_current_offset,
  input  [15:0]  io_pipe_phv_in_parse_transition_field,
  input  [2:0]   io_pipe_phv_in_next_processor_id,
  input          io_pipe_phv_in_next_config_id,
  input          io_pipe_phv_in_is_valid_processor,
  output [7:0]   io_pipe_phv_out_data_0,
  output [7:0]   io_pipe_phv_out_data_1,
  output [7:0]   io_pipe_phv_out_data_2,
  output [7:0]   io_pipe_phv_out_data_3,
  output [7:0]   io_pipe_phv_out_data_4,
  output [7:0]   io_pipe_phv_out_data_5,
  output [7:0]   io_pipe_phv_out_data_6,
  output [7:0]   io_pipe_phv_out_data_7,
  output [7:0]   io_pipe_phv_out_data_8,
  output [7:0]   io_pipe_phv_out_data_9,
  output [7:0]   io_pipe_phv_out_data_10,
  output [7:0]   io_pipe_phv_out_data_11,
  output [7:0]   io_pipe_phv_out_data_12,
  output [7:0]   io_pipe_phv_out_data_13,
  output [7:0]   io_pipe_phv_out_data_14,
  output [7:0]   io_pipe_phv_out_data_15,
  output [7:0]   io_pipe_phv_out_data_16,
  output [7:0]   io_pipe_phv_out_data_17,
  output [7:0]   io_pipe_phv_out_data_18,
  output [7:0]   io_pipe_phv_out_data_19,
  output [7:0]   io_pipe_phv_out_data_20,
  output [7:0]   io_pipe_phv_out_data_21,
  output [7:0]   io_pipe_phv_out_data_22,
  output [7:0]   io_pipe_phv_out_data_23,
  output [7:0]   io_pipe_phv_out_data_24,
  output [7:0]   io_pipe_phv_out_data_25,
  output [7:0]   io_pipe_phv_out_data_26,
  output [7:0]   io_pipe_phv_out_data_27,
  output [7:0]   io_pipe_phv_out_data_28,
  output [7:0]   io_pipe_phv_out_data_29,
  output [7:0]   io_pipe_phv_out_data_30,
  output [7:0]   io_pipe_phv_out_data_31,
  output [7:0]   io_pipe_phv_out_data_32,
  output [7:0]   io_pipe_phv_out_data_33,
  output [7:0]   io_pipe_phv_out_data_34,
  output [7:0]   io_pipe_phv_out_data_35,
  output [7:0]   io_pipe_phv_out_data_36,
  output [7:0]   io_pipe_phv_out_data_37,
  output [7:0]   io_pipe_phv_out_data_38,
  output [7:0]   io_pipe_phv_out_data_39,
  output [7:0]   io_pipe_phv_out_data_40,
  output [7:0]   io_pipe_phv_out_data_41,
  output [7:0]   io_pipe_phv_out_data_42,
  output [7:0]   io_pipe_phv_out_data_43,
  output [7:0]   io_pipe_phv_out_data_44,
  output [7:0]   io_pipe_phv_out_data_45,
  output [7:0]   io_pipe_phv_out_data_46,
  output [7:0]   io_pipe_phv_out_data_47,
  output [7:0]   io_pipe_phv_out_data_48,
  output [7:0]   io_pipe_phv_out_data_49,
  output [7:0]   io_pipe_phv_out_data_50,
  output [7:0]   io_pipe_phv_out_data_51,
  output [7:0]   io_pipe_phv_out_data_52,
  output [7:0]   io_pipe_phv_out_data_53,
  output [7:0]   io_pipe_phv_out_data_54,
  output [7:0]   io_pipe_phv_out_data_55,
  output [7:0]   io_pipe_phv_out_data_56,
  output [7:0]   io_pipe_phv_out_data_57,
  output [7:0]   io_pipe_phv_out_data_58,
  output [7:0]   io_pipe_phv_out_data_59,
  output [7:0]   io_pipe_phv_out_data_60,
  output [7:0]   io_pipe_phv_out_data_61,
  output [7:0]   io_pipe_phv_out_data_62,
  output [7:0]   io_pipe_phv_out_data_63,
  output [7:0]   io_pipe_phv_out_data_64,
  output [7:0]   io_pipe_phv_out_data_65,
  output [7:0]   io_pipe_phv_out_data_66,
  output [7:0]   io_pipe_phv_out_data_67,
  output [7:0]   io_pipe_phv_out_data_68,
  output [7:0]   io_pipe_phv_out_data_69,
  output [7:0]   io_pipe_phv_out_data_70,
  output [7:0]   io_pipe_phv_out_data_71,
  output [7:0]   io_pipe_phv_out_data_72,
  output [7:0]   io_pipe_phv_out_data_73,
  output [7:0]   io_pipe_phv_out_data_74,
  output [7:0]   io_pipe_phv_out_data_75,
  output [7:0]   io_pipe_phv_out_data_76,
  output [7:0]   io_pipe_phv_out_data_77,
  output [7:0]   io_pipe_phv_out_data_78,
  output [7:0]   io_pipe_phv_out_data_79,
  output [7:0]   io_pipe_phv_out_data_80,
  output [7:0]   io_pipe_phv_out_data_81,
  output [7:0]   io_pipe_phv_out_data_82,
  output [7:0]   io_pipe_phv_out_data_83,
  output [7:0]   io_pipe_phv_out_data_84,
  output [7:0]   io_pipe_phv_out_data_85,
  output [7:0]   io_pipe_phv_out_data_86,
  output [7:0]   io_pipe_phv_out_data_87,
  output [7:0]   io_pipe_phv_out_data_88,
  output [7:0]   io_pipe_phv_out_data_89,
  output [7:0]   io_pipe_phv_out_data_90,
  output [7:0]   io_pipe_phv_out_data_91,
  output [7:0]   io_pipe_phv_out_data_92,
  output [7:0]   io_pipe_phv_out_data_93,
  output [7:0]   io_pipe_phv_out_data_94,
  output [7:0]   io_pipe_phv_out_data_95,
  output [7:0]   io_pipe_phv_out_data_96,
  output [7:0]   io_pipe_phv_out_data_97,
  output [7:0]   io_pipe_phv_out_data_98,
  output [7:0]   io_pipe_phv_out_data_99,
  output [7:0]   io_pipe_phv_out_data_100,
  output [7:0]   io_pipe_phv_out_data_101,
  output [7:0]   io_pipe_phv_out_data_102,
  output [7:0]   io_pipe_phv_out_data_103,
  output [7:0]   io_pipe_phv_out_data_104,
  output [7:0]   io_pipe_phv_out_data_105,
  output [7:0]   io_pipe_phv_out_data_106,
  output [7:0]   io_pipe_phv_out_data_107,
  output [7:0]   io_pipe_phv_out_data_108,
  output [7:0]   io_pipe_phv_out_data_109,
  output [7:0]   io_pipe_phv_out_data_110,
  output [7:0]   io_pipe_phv_out_data_111,
  output [7:0]   io_pipe_phv_out_data_112,
  output [7:0]   io_pipe_phv_out_data_113,
  output [7:0]   io_pipe_phv_out_data_114,
  output [7:0]   io_pipe_phv_out_data_115,
  output [7:0]   io_pipe_phv_out_data_116,
  output [7:0]   io_pipe_phv_out_data_117,
  output [7:0]   io_pipe_phv_out_data_118,
  output [7:0]   io_pipe_phv_out_data_119,
  output [7:0]   io_pipe_phv_out_data_120,
  output [7:0]   io_pipe_phv_out_data_121,
  output [7:0]   io_pipe_phv_out_data_122,
  output [7:0]   io_pipe_phv_out_data_123,
  output [7:0]   io_pipe_phv_out_data_124,
  output [7:0]   io_pipe_phv_out_data_125,
  output [7:0]   io_pipe_phv_out_data_126,
  output [7:0]   io_pipe_phv_out_data_127,
  output [7:0]   io_pipe_phv_out_data_128,
  output [7:0]   io_pipe_phv_out_data_129,
  output [7:0]   io_pipe_phv_out_data_130,
  output [7:0]   io_pipe_phv_out_data_131,
  output [7:0]   io_pipe_phv_out_data_132,
  output [7:0]   io_pipe_phv_out_data_133,
  output [7:0]   io_pipe_phv_out_data_134,
  output [7:0]   io_pipe_phv_out_data_135,
  output [7:0]   io_pipe_phv_out_data_136,
  output [7:0]   io_pipe_phv_out_data_137,
  output [7:0]   io_pipe_phv_out_data_138,
  output [7:0]   io_pipe_phv_out_data_139,
  output [7:0]   io_pipe_phv_out_data_140,
  output [7:0]   io_pipe_phv_out_data_141,
  output [7:0]   io_pipe_phv_out_data_142,
  output [7:0]   io_pipe_phv_out_data_143,
  output [7:0]   io_pipe_phv_out_data_144,
  output [7:0]   io_pipe_phv_out_data_145,
  output [7:0]   io_pipe_phv_out_data_146,
  output [7:0]   io_pipe_phv_out_data_147,
  output [7:0]   io_pipe_phv_out_data_148,
  output [7:0]   io_pipe_phv_out_data_149,
  output [7:0]   io_pipe_phv_out_data_150,
  output [7:0]   io_pipe_phv_out_data_151,
  output [7:0]   io_pipe_phv_out_data_152,
  output [7:0]   io_pipe_phv_out_data_153,
  output [7:0]   io_pipe_phv_out_data_154,
  output [7:0]   io_pipe_phv_out_data_155,
  output [7:0]   io_pipe_phv_out_data_156,
  output [7:0]   io_pipe_phv_out_data_157,
  output [7:0]   io_pipe_phv_out_data_158,
  output [7:0]   io_pipe_phv_out_data_159,
  output [7:0]   io_pipe_phv_out_data_160,
  output [7:0]   io_pipe_phv_out_data_161,
  output [7:0]   io_pipe_phv_out_data_162,
  output [7:0]   io_pipe_phv_out_data_163,
  output [7:0]   io_pipe_phv_out_data_164,
  output [7:0]   io_pipe_phv_out_data_165,
  output [7:0]   io_pipe_phv_out_data_166,
  output [7:0]   io_pipe_phv_out_data_167,
  output [7:0]   io_pipe_phv_out_data_168,
  output [7:0]   io_pipe_phv_out_data_169,
  output [7:0]   io_pipe_phv_out_data_170,
  output [7:0]   io_pipe_phv_out_data_171,
  output [7:0]   io_pipe_phv_out_data_172,
  output [7:0]   io_pipe_phv_out_data_173,
  output [7:0]   io_pipe_phv_out_data_174,
  output [7:0]   io_pipe_phv_out_data_175,
  output [7:0]   io_pipe_phv_out_data_176,
  output [7:0]   io_pipe_phv_out_data_177,
  output [7:0]   io_pipe_phv_out_data_178,
  output [7:0]   io_pipe_phv_out_data_179,
  output [7:0]   io_pipe_phv_out_data_180,
  output [7:0]   io_pipe_phv_out_data_181,
  output [7:0]   io_pipe_phv_out_data_182,
  output [7:0]   io_pipe_phv_out_data_183,
  output [7:0]   io_pipe_phv_out_data_184,
  output [7:0]   io_pipe_phv_out_data_185,
  output [7:0]   io_pipe_phv_out_data_186,
  output [7:0]   io_pipe_phv_out_data_187,
  output [7:0]   io_pipe_phv_out_data_188,
  output [7:0]   io_pipe_phv_out_data_189,
  output [7:0]   io_pipe_phv_out_data_190,
  output [7:0]   io_pipe_phv_out_data_191,
  output [7:0]   io_pipe_phv_out_data_192,
  output [7:0]   io_pipe_phv_out_data_193,
  output [7:0]   io_pipe_phv_out_data_194,
  output [7:0]   io_pipe_phv_out_data_195,
  output [7:0]   io_pipe_phv_out_data_196,
  output [7:0]   io_pipe_phv_out_data_197,
  output [7:0]   io_pipe_phv_out_data_198,
  output [7:0]   io_pipe_phv_out_data_199,
  output [7:0]   io_pipe_phv_out_data_200,
  output [7:0]   io_pipe_phv_out_data_201,
  output [7:0]   io_pipe_phv_out_data_202,
  output [7:0]   io_pipe_phv_out_data_203,
  output [7:0]   io_pipe_phv_out_data_204,
  output [7:0]   io_pipe_phv_out_data_205,
  output [7:0]   io_pipe_phv_out_data_206,
  output [7:0]   io_pipe_phv_out_data_207,
  output [7:0]   io_pipe_phv_out_data_208,
  output [7:0]   io_pipe_phv_out_data_209,
  output [7:0]   io_pipe_phv_out_data_210,
  output [7:0]   io_pipe_phv_out_data_211,
  output [7:0]   io_pipe_phv_out_data_212,
  output [7:0]   io_pipe_phv_out_data_213,
  output [7:0]   io_pipe_phv_out_data_214,
  output [7:0]   io_pipe_phv_out_data_215,
  output [7:0]   io_pipe_phv_out_data_216,
  output [7:0]   io_pipe_phv_out_data_217,
  output [7:0]   io_pipe_phv_out_data_218,
  output [7:0]   io_pipe_phv_out_data_219,
  output [7:0]   io_pipe_phv_out_data_220,
  output [7:0]   io_pipe_phv_out_data_221,
  output [7:0]   io_pipe_phv_out_data_222,
  output [7:0]   io_pipe_phv_out_data_223,
  output [7:0]   io_pipe_phv_out_data_224,
  output [7:0]   io_pipe_phv_out_data_225,
  output [7:0]   io_pipe_phv_out_data_226,
  output [7:0]   io_pipe_phv_out_data_227,
  output [7:0]   io_pipe_phv_out_data_228,
  output [7:0]   io_pipe_phv_out_data_229,
  output [7:0]   io_pipe_phv_out_data_230,
  output [7:0]   io_pipe_phv_out_data_231,
  output [7:0]   io_pipe_phv_out_data_232,
  output [7:0]   io_pipe_phv_out_data_233,
  output [7:0]   io_pipe_phv_out_data_234,
  output [7:0]   io_pipe_phv_out_data_235,
  output [7:0]   io_pipe_phv_out_data_236,
  output [7:0]   io_pipe_phv_out_data_237,
  output [7:0]   io_pipe_phv_out_data_238,
  output [7:0]   io_pipe_phv_out_data_239,
  output [7:0]   io_pipe_phv_out_data_240,
  output [7:0]   io_pipe_phv_out_data_241,
  output [7:0]   io_pipe_phv_out_data_242,
  output [7:0]   io_pipe_phv_out_data_243,
  output [7:0]   io_pipe_phv_out_data_244,
  output [7:0]   io_pipe_phv_out_data_245,
  output [7:0]   io_pipe_phv_out_data_246,
  output [7:0]   io_pipe_phv_out_data_247,
  output [7:0]   io_pipe_phv_out_data_248,
  output [7:0]   io_pipe_phv_out_data_249,
  output [7:0]   io_pipe_phv_out_data_250,
  output [7:0]   io_pipe_phv_out_data_251,
  output [7:0]   io_pipe_phv_out_data_252,
  output [7:0]   io_pipe_phv_out_data_253,
  output [7:0]   io_pipe_phv_out_data_254,
  output [7:0]   io_pipe_phv_out_data_255,
  output [15:0]  io_pipe_phv_out_header_0,
  output [15:0]  io_pipe_phv_out_header_1,
  output [15:0]  io_pipe_phv_out_header_2,
  output [15:0]  io_pipe_phv_out_header_3,
  output [15:0]  io_pipe_phv_out_header_4,
  output [15:0]  io_pipe_phv_out_header_5,
  output [15:0]  io_pipe_phv_out_header_6,
  output [15:0]  io_pipe_phv_out_header_7,
  output [15:0]  io_pipe_phv_out_header_8,
  output [15:0]  io_pipe_phv_out_header_9,
  output [15:0]  io_pipe_phv_out_header_10,
  output [15:0]  io_pipe_phv_out_header_11,
  output [15:0]  io_pipe_phv_out_header_12,
  output [15:0]  io_pipe_phv_out_header_13,
  output [15:0]  io_pipe_phv_out_header_14,
  output [15:0]  io_pipe_phv_out_header_15,
  output [7:0]   io_pipe_phv_out_parse_current_state,
  output [7:0]   io_pipe_phv_out_parse_current_offset,
  output [15:0]  io_pipe_phv_out_parse_transition_field,
  output [2:0]   io_pipe_phv_out_next_processor_id,
  output         io_pipe_phv_out_next_config_id,
  output         io_pipe_phv_out_is_valid_processor,
  input  [7:0]   io_key_config_0_key_length,
  input  [7:0]   io_key_config_1_key_length,
  input  [191:0] io_key_in,
  input  [255:0] io_data_in,
  output         io_hit,
  output [63:0]  io_match_value
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [191:0] _RAND_278;
  reg [255:0] _RAND_279;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[matcher.scala 311:22]
  reg [7:0] phv_data_1; // @[matcher.scala 311:22]
  reg [7:0] phv_data_2; // @[matcher.scala 311:22]
  reg [7:0] phv_data_3; // @[matcher.scala 311:22]
  reg [7:0] phv_data_4; // @[matcher.scala 311:22]
  reg [7:0] phv_data_5; // @[matcher.scala 311:22]
  reg [7:0] phv_data_6; // @[matcher.scala 311:22]
  reg [7:0] phv_data_7; // @[matcher.scala 311:22]
  reg [7:0] phv_data_8; // @[matcher.scala 311:22]
  reg [7:0] phv_data_9; // @[matcher.scala 311:22]
  reg [7:0] phv_data_10; // @[matcher.scala 311:22]
  reg [7:0] phv_data_11; // @[matcher.scala 311:22]
  reg [7:0] phv_data_12; // @[matcher.scala 311:22]
  reg [7:0] phv_data_13; // @[matcher.scala 311:22]
  reg [7:0] phv_data_14; // @[matcher.scala 311:22]
  reg [7:0] phv_data_15; // @[matcher.scala 311:22]
  reg [7:0] phv_data_16; // @[matcher.scala 311:22]
  reg [7:0] phv_data_17; // @[matcher.scala 311:22]
  reg [7:0] phv_data_18; // @[matcher.scala 311:22]
  reg [7:0] phv_data_19; // @[matcher.scala 311:22]
  reg [7:0] phv_data_20; // @[matcher.scala 311:22]
  reg [7:0] phv_data_21; // @[matcher.scala 311:22]
  reg [7:0] phv_data_22; // @[matcher.scala 311:22]
  reg [7:0] phv_data_23; // @[matcher.scala 311:22]
  reg [7:0] phv_data_24; // @[matcher.scala 311:22]
  reg [7:0] phv_data_25; // @[matcher.scala 311:22]
  reg [7:0] phv_data_26; // @[matcher.scala 311:22]
  reg [7:0] phv_data_27; // @[matcher.scala 311:22]
  reg [7:0] phv_data_28; // @[matcher.scala 311:22]
  reg [7:0] phv_data_29; // @[matcher.scala 311:22]
  reg [7:0] phv_data_30; // @[matcher.scala 311:22]
  reg [7:0] phv_data_31; // @[matcher.scala 311:22]
  reg [7:0] phv_data_32; // @[matcher.scala 311:22]
  reg [7:0] phv_data_33; // @[matcher.scala 311:22]
  reg [7:0] phv_data_34; // @[matcher.scala 311:22]
  reg [7:0] phv_data_35; // @[matcher.scala 311:22]
  reg [7:0] phv_data_36; // @[matcher.scala 311:22]
  reg [7:0] phv_data_37; // @[matcher.scala 311:22]
  reg [7:0] phv_data_38; // @[matcher.scala 311:22]
  reg [7:0] phv_data_39; // @[matcher.scala 311:22]
  reg [7:0] phv_data_40; // @[matcher.scala 311:22]
  reg [7:0] phv_data_41; // @[matcher.scala 311:22]
  reg [7:0] phv_data_42; // @[matcher.scala 311:22]
  reg [7:0] phv_data_43; // @[matcher.scala 311:22]
  reg [7:0] phv_data_44; // @[matcher.scala 311:22]
  reg [7:0] phv_data_45; // @[matcher.scala 311:22]
  reg [7:0] phv_data_46; // @[matcher.scala 311:22]
  reg [7:0] phv_data_47; // @[matcher.scala 311:22]
  reg [7:0] phv_data_48; // @[matcher.scala 311:22]
  reg [7:0] phv_data_49; // @[matcher.scala 311:22]
  reg [7:0] phv_data_50; // @[matcher.scala 311:22]
  reg [7:0] phv_data_51; // @[matcher.scala 311:22]
  reg [7:0] phv_data_52; // @[matcher.scala 311:22]
  reg [7:0] phv_data_53; // @[matcher.scala 311:22]
  reg [7:0] phv_data_54; // @[matcher.scala 311:22]
  reg [7:0] phv_data_55; // @[matcher.scala 311:22]
  reg [7:0] phv_data_56; // @[matcher.scala 311:22]
  reg [7:0] phv_data_57; // @[matcher.scala 311:22]
  reg [7:0] phv_data_58; // @[matcher.scala 311:22]
  reg [7:0] phv_data_59; // @[matcher.scala 311:22]
  reg [7:0] phv_data_60; // @[matcher.scala 311:22]
  reg [7:0] phv_data_61; // @[matcher.scala 311:22]
  reg [7:0] phv_data_62; // @[matcher.scala 311:22]
  reg [7:0] phv_data_63; // @[matcher.scala 311:22]
  reg [7:0] phv_data_64; // @[matcher.scala 311:22]
  reg [7:0] phv_data_65; // @[matcher.scala 311:22]
  reg [7:0] phv_data_66; // @[matcher.scala 311:22]
  reg [7:0] phv_data_67; // @[matcher.scala 311:22]
  reg [7:0] phv_data_68; // @[matcher.scala 311:22]
  reg [7:0] phv_data_69; // @[matcher.scala 311:22]
  reg [7:0] phv_data_70; // @[matcher.scala 311:22]
  reg [7:0] phv_data_71; // @[matcher.scala 311:22]
  reg [7:0] phv_data_72; // @[matcher.scala 311:22]
  reg [7:0] phv_data_73; // @[matcher.scala 311:22]
  reg [7:0] phv_data_74; // @[matcher.scala 311:22]
  reg [7:0] phv_data_75; // @[matcher.scala 311:22]
  reg [7:0] phv_data_76; // @[matcher.scala 311:22]
  reg [7:0] phv_data_77; // @[matcher.scala 311:22]
  reg [7:0] phv_data_78; // @[matcher.scala 311:22]
  reg [7:0] phv_data_79; // @[matcher.scala 311:22]
  reg [7:0] phv_data_80; // @[matcher.scala 311:22]
  reg [7:0] phv_data_81; // @[matcher.scala 311:22]
  reg [7:0] phv_data_82; // @[matcher.scala 311:22]
  reg [7:0] phv_data_83; // @[matcher.scala 311:22]
  reg [7:0] phv_data_84; // @[matcher.scala 311:22]
  reg [7:0] phv_data_85; // @[matcher.scala 311:22]
  reg [7:0] phv_data_86; // @[matcher.scala 311:22]
  reg [7:0] phv_data_87; // @[matcher.scala 311:22]
  reg [7:0] phv_data_88; // @[matcher.scala 311:22]
  reg [7:0] phv_data_89; // @[matcher.scala 311:22]
  reg [7:0] phv_data_90; // @[matcher.scala 311:22]
  reg [7:0] phv_data_91; // @[matcher.scala 311:22]
  reg [7:0] phv_data_92; // @[matcher.scala 311:22]
  reg [7:0] phv_data_93; // @[matcher.scala 311:22]
  reg [7:0] phv_data_94; // @[matcher.scala 311:22]
  reg [7:0] phv_data_95; // @[matcher.scala 311:22]
  reg [7:0] phv_data_96; // @[matcher.scala 311:22]
  reg [7:0] phv_data_97; // @[matcher.scala 311:22]
  reg [7:0] phv_data_98; // @[matcher.scala 311:22]
  reg [7:0] phv_data_99; // @[matcher.scala 311:22]
  reg [7:0] phv_data_100; // @[matcher.scala 311:22]
  reg [7:0] phv_data_101; // @[matcher.scala 311:22]
  reg [7:0] phv_data_102; // @[matcher.scala 311:22]
  reg [7:0] phv_data_103; // @[matcher.scala 311:22]
  reg [7:0] phv_data_104; // @[matcher.scala 311:22]
  reg [7:0] phv_data_105; // @[matcher.scala 311:22]
  reg [7:0] phv_data_106; // @[matcher.scala 311:22]
  reg [7:0] phv_data_107; // @[matcher.scala 311:22]
  reg [7:0] phv_data_108; // @[matcher.scala 311:22]
  reg [7:0] phv_data_109; // @[matcher.scala 311:22]
  reg [7:0] phv_data_110; // @[matcher.scala 311:22]
  reg [7:0] phv_data_111; // @[matcher.scala 311:22]
  reg [7:0] phv_data_112; // @[matcher.scala 311:22]
  reg [7:0] phv_data_113; // @[matcher.scala 311:22]
  reg [7:0] phv_data_114; // @[matcher.scala 311:22]
  reg [7:0] phv_data_115; // @[matcher.scala 311:22]
  reg [7:0] phv_data_116; // @[matcher.scala 311:22]
  reg [7:0] phv_data_117; // @[matcher.scala 311:22]
  reg [7:0] phv_data_118; // @[matcher.scala 311:22]
  reg [7:0] phv_data_119; // @[matcher.scala 311:22]
  reg [7:0] phv_data_120; // @[matcher.scala 311:22]
  reg [7:0] phv_data_121; // @[matcher.scala 311:22]
  reg [7:0] phv_data_122; // @[matcher.scala 311:22]
  reg [7:0] phv_data_123; // @[matcher.scala 311:22]
  reg [7:0] phv_data_124; // @[matcher.scala 311:22]
  reg [7:0] phv_data_125; // @[matcher.scala 311:22]
  reg [7:0] phv_data_126; // @[matcher.scala 311:22]
  reg [7:0] phv_data_127; // @[matcher.scala 311:22]
  reg [7:0] phv_data_128; // @[matcher.scala 311:22]
  reg [7:0] phv_data_129; // @[matcher.scala 311:22]
  reg [7:0] phv_data_130; // @[matcher.scala 311:22]
  reg [7:0] phv_data_131; // @[matcher.scala 311:22]
  reg [7:0] phv_data_132; // @[matcher.scala 311:22]
  reg [7:0] phv_data_133; // @[matcher.scala 311:22]
  reg [7:0] phv_data_134; // @[matcher.scala 311:22]
  reg [7:0] phv_data_135; // @[matcher.scala 311:22]
  reg [7:0] phv_data_136; // @[matcher.scala 311:22]
  reg [7:0] phv_data_137; // @[matcher.scala 311:22]
  reg [7:0] phv_data_138; // @[matcher.scala 311:22]
  reg [7:0] phv_data_139; // @[matcher.scala 311:22]
  reg [7:0] phv_data_140; // @[matcher.scala 311:22]
  reg [7:0] phv_data_141; // @[matcher.scala 311:22]
  reg [7:0] phv_data_142; // @[matcher.scala 311:22]
  reg [7:0] phv_data_143; // @[matcher.scala 311:22]
  reg [7:0] phv_data_144; // @[matcher.scala 311:22]
  reg [7:0] phv_data_145; // @[matcher.scala 311:22]
  reg [7:0] phv_data_146; // @[matcher.scala 311:22]
  reg [7:0] phv_data_147; // @[matcher.scala 311:22]
  reg [7:0] phv_data_148; // @[matcher.scala 311:22]
  reg [7:0] phv_data_149; // @[matcher.scala 311:22]
  reg [7:0] phv_data_150; // @[matcher.scala 311:22]
  reg [7:0] phv_data_151; // @[matcher.scala 311:22]
  reg [7:0] phv_data_152; // @[matcher.scala 311:22]
  reg [7:0] phv_data_153; // @[matcher.scala 311:22]
  reg [7:0] phv_data_154; // @[matcher.scala 311:22]
  reg [7:0] phv_data_155; // @[matcher.scala 311:22]
  reg [7:0] phv_data_156; // @[matcher.scala 311:22]
  reg [7:0] phv_data_157; // @[matcher.scala 311:22]
  reg [7:0] phv_data_158; // @[matcher.scala 311:22]
  reg [7:0] phv_data_159; // @[matcher.scala 311:22]
  reg [7:0] phv_data_160; // @[matcher.scala 311:22]
  reg [7:0] phv_data_161; // @[matcher.scala 311:22]
  reg [7:0] phv_data_162; // @[matcher.scala 311:22]
  reg [7:0] phv_data_163; // @[matcher.scala 311:22]
  reg [7:0] phv_data_164; // @[matcher.scala 311:22]
  reg [7:0] phv_data_165; // @[matcher.scala 311:22]
  reg [7:0] phv_data_166; // @[matcher.scala 311:22]
  reg [7:0] phv_data_167; // @[matcher.scala 311:22]
  reg [7:0] phv_data_168; // @[matcher.scala 311:22]
  reg [7:0] phv_data_169; // @[matcher.scala 311:22]
  reg [7:0] phv_data_170; // @[matcher.scala 311:22]
  reg [7:0] phv_data_171; // @[matcher.scala 311:22]
  reg [7:0] phv_data_172; // @[matcher.scala 311:22]
  reg [7:0] phv_data_173; // @[matcher.scala 311:22]
  reg [7:0] phv_data_174; // @[matcher.scala 311:22]
  reg [7:0] phv_data_175; // @[matcher.scala 311:22]
  reg [7:0] phv_data_176; // @[matcher.scala 311:22]
  reg [7:0] phv_data_177; // @[matcher.scala 311:22]
  reg [7:0] phv_data_178; // @[matcher.scala 311:22]
  reg [7:0] phv_data_179; // @[matcher.scala 311:22]
  reg [7:0] phv_data_180; // @[matcher.scala 311:22]
  reg [7:0] phv_data_181; // @[matcher.scala 311:22]
  reg [7:0] phv_data_182; // @[matcher.scala 311:22]
  reg [7:0] phv_data_183; // @[matcher.scala 311:22]
  reg [7:0] phv_data_184; // @[matcher.scala 311:22]
  reg [7:0] phv_data_185; // @[matcher.scala 311:22]
  reg [7:0] phv_data_186; // @[matcher.scala 311:22]
  reg [7:0] phv_data_187; // @[matcher.scala 311:22]
  reg [7:0] phv_data_188; // @[matcher.scala 311:22]
  reg [7:0] phv_data_189; // @[matcher.scala 311:22]
  reg [7:0] phv_data_190; // @[matcher.scala 311:22]
  reg [7:0] phv_data_191; // @[matcher.scala 311:22]
  reg [7:0] phv_data_192; // @[matcher.scala 311:22]
  reg [7:0] phv_data_193; // @[matcher.scala 311:22]
  reg [7:0] phv_data_194; // @[matcher.scala 311:22]
  reg [7:0] phv_data_195; // @[matcher.scala 311:22]
  reg [7:0] phv_data_196; // @[matcher.scala 311:22]
  reg [7:0] phv_data_197; // @[matcher.scala 311:22]
  reg [7:0] phv_data_198; // @[matcher.scala 311:22]
  reg [7:0] phv_data_199; // @[matcher.scala 311:22]
  reg [7:0] phv_data_200; // @[matcher.scala 311:22]
  reg [7:0] phv_data_201; // @[matcher.scala 311:22]
  reg [7:0] phv_data_202; // @[matcher.scala 311:22]
  reg [7:0] phv_data_203; // @[matcher.scala 311:22]
  reg [7:0] phv_data_204; // @[matcher.scala 311:22]
  reg [7:0] phv_data_205; // @[matcher.scala 311:22]
  reg [7:0] phv_data_206; // @[matcher.scala 311:22]
  reg [7:0] phv_data_207; // @[matcher.scala 311:22]
  reg [7:0] phv_data_208; // @[matcher.scala 311:22]
  reg [7:0] phv_data_209; // @[matcher.scala 311:22]
  reg [7:0] phv_data_210; // @[matcher.scala 311:22]
  reg [7:0] phv_data_211; // @[matcher.scala 311:22]
  reg [7:0] phv_data_212; // @[matcher.scala 311:22]
  reg [7:0] phv_data_213; // @[matcher.scala 311:22]
  reg [7:0] phv_data_214; // @[matcher.scala 311:22]
  reg [7:0] phv_data_215; // @[matcher.scala 311:22]
  reg [7:0] phv_data_216; // @[matcher.scala 311:22]
  reg [7:0] phv_data_217; // @[matcher.scala 311:22]
  reg [7:0] phv_data_218; // @[matcher.scala 311:22]
  reg [7:0] phv_data_219; // @[matcher.scala 311:22]
  reg [7:0] phv_data_220; // @[matcher.scala 311:22]
  reg [7:0] phv_data_221; // @[matcher.scala 311:22]
  reg [7:0] phv_data_222; // @[matcher.scala 311:22]
  reg [7:0] phv_data_223; // @[matcher.scala 311:22]
  reg [7:0] phv_data_224; // @[matcher.scala 311:22]
  reg [7:0] phv_data_225; // @[matcher.scala 311:22]
  reg [7:0] phv_data_226; // @[matcher.scala 311:22]
  reg [7:0] phv_data_227; // @[matcher.scala 311:22]
  reg [7:0] phv_data_228; // @[matcher.scala 311:22]
  reg [7:0] phv_data_229; // @[matcher.scala 311:22]
  reg [7:0] phv_data_230; // @[matcher.scala 311:22]
  reg [7:0] phv_data_231; // @[matcher.scala 311:22]
  reg [7:0] phv_data_232; // @[matcher.scala 311:22]
  reg [7:0] phv_data_233; // @[matcher.scala 311:22]
  reg [7:0] phv_data_234; // @[matcher.scala 311:22]
  reg [7:0] phv_data_235; // @[matcher.scala 311:22]
  reg [7:0] phv_data_236; // @[matcher.scala 311:22]
  reg [7:0] phv_data_237; // @[matcher.scala 311:22]
  reg [7:0] phv_data_238; // @[matcher.scala 311:22]
  reg [7:0] phv_data_239; // @[matcher.scala 311:22]
  reg [7:0] phv_data_240; // @[matcher.scala 311:22]
  reg [7:0] phv_data_241; // @[matcher.scala 311:22]
  reg [7:0] phv_data_242; // @[matcher.scala 311:22]
  reg [7:0] phv_data_243; // @[matcher.scala 311:22]
  reg [7:0] phv_data_244; // @[matcher.scala 311:22]
  reg [7:0] phv_data_245; // @[matcher.scala 311:22]
  reg [7:0] phv_data_246; // @[matcher.scala 311:22]
  reg [7:0] phv_data_247; // @[matcher.scala 311:22]
  reg [7:0] phv_data_248; // @[matcher.scala 311:22]
  reg [7:0] phv_data_249; // @[matcher.scala 311:22]
  reg [7:0] phv_data_250; // @[matcher.scala 311:22]
  reg [7:0] phv_data_251; // @[matcher.scala 311:22]
  reg [7:0] phv_data_252; // @[matcher.scala 311:22]
  reg [7:0] phv_data_253; // @[matcher.scala 311:22]
  reg [7:0] phv_data_254; // @[matcher.scala 311:22]
  reg [7:0] phv_data_255; // @[matcher.scala 311:22]
  reg [15:0] phv_header_0; // @[matcher.scala 311:22]
  reg [15:0] phv_header_1; // @[matcher.scala 311:22]
  reg [15:0] phv_header_2; // @[matcher.scala 311:22]
  reg [15:0] phv_header_3; // @[matcher.scala 311:22]
  reg [15:0] phv_header_4; // @[matcher.scala 311:22]
  reg [15:0] phv_header_5; // @[matcher.scala 311:22]
  reg [15:0] phv_header_6; // @[matcher.scala 311:22]
  reg [15:0] phv_header_7; // @[matcher.scala 311:22]
  reg [15:0] phv_header_8; // @[matcher.scala 311:22]
  reg [15:0] phv_header_9; // @[matcher.scala 311:22]
  reg [15:0] phv_header_10; // @[matcher.scala 311:22]
  reg [15:0] phv_header_11; // @[matcher.scala 311:22]
  reg [15:0] phv_header_12; // @[matcher.scala 311:22]
  reg [15:0] phv_header_13; // @[matcher.scala 311:22]
  reg [15:0] phv_header_14; // @[matcher.scala 311:22]
  reg [15:0] phv_header_15; // @[matcher.scala 311:22]
  reg [7:0] phv_parse_current_state; // @[matcher.scala 311:22]
  reg [7:0] phv_parse_current_offset; // @[matcher.scala 311:22]
  reg [15:0] phv_parse_transition_field; // @[matcher.scala 311:22]
  reg [2:0] phv_next_processor_id; // @[matcher.scala 311:22]
  reg  phv_next_config_id; // @[matcher.scala 311:22]
  reg  phv_is_valid_processor; // @[matcher.scala 311:22]
  reg [191:0] key; // @[matcher.scala 315:22]
  reg [255:0] data; // @[matcher.scala 317:23]
  wire [7:0] key_byte = key[7:0]; // @[matcher.scala 325:35]
  wire [7:0] data_byte = data[71:64]; // @[matcher.scala 326:37]
  wire [7:0] _GEN_6 = phv_next_config_id ? io_key_config_1_key_length : io_key_config_0_key_length; // @[matcher.scala 327:65 matcher.scala 327:65]
  wire  key_equal_0 = 8'h0 < _GEN_6 ? key_byte == data_byte : 1'h1; // @[matcher.scala 327:90 matcher.scala 328:34 matcher.scala 330:34]
  wire [7:0] key_byte_1 = key[15:8]; // @[matcher.scala 325:35]
  wire [7:0] data_byte_1 = data[79:72]; // @[matcher.scala 326:37]
  wire  key_equal_1 = 8'h1 < _GEN_6 ? key_byte_1 == data_byte_1 : 1'h1; // @[matcher.scala 327:90 matcher.scala 328:34 matcher.scala 330:34]
  wire [7:0] key_byte_2 = key[23:16]; // @[matcher.scala 325:35]
  wire [7:0] data_byte_2 = data[87:80]; // @[matcher.scala 326:37]
  wire  key_equal_2 = 8'h2 < _GEN_6 ? key_byte_2 == data_byte_2 : 1'h1; // @[matcher.scala 327:90 matcher.scala 328:34 matcher.scala 330:34]
  wire [7:0] key_byte_3 = key[31:24]; // @[matcher.scala 325:35]
  wire [7:0] data_byte_3 = data[95:88]; // @[matcher.scala 326:37]
  wire  key_equal_3 = 8'h3 < _GEN_6 ? key_byte_3 == data_byte_3 : 1'h1; // @[matcher.scala 327:90 matcher.scala 328:34 matcher.scala 330:34]
  wire [7:0] key_byte_4 = key[39:32]; // @[matcher.scala 325:35]
  wire [7:0] data_byte_4 = data[103:96]; // @[matcher.scala 326:37]
  wire  key_equal_4 = 8'h4 < _GEN_6 ? key_byte_4 == data_byte_4 : 1'h1; // @[matcher.scala 327:90 matcher.scala 328:34 matcher.scala 330:34]
  wire [7:0] key_byte_5 = key[47:40]; // @[matcher.scala 325:35]
  wire [7:0] data_byte_5 = data[111:104]; // @[matcher.scala 326:37]
  wire  key_equal_5 = 8'h5 < _GEN_6 ? key_byte_5 == data_byte_5 : 1'h1; // @[matcher.scala 327:90 matcher.scala 328:34 matcher.scala 330:34]
  wire [7:0] key_byte_6 = key[55:48]; // @[matcher.scala 325:35]
  wire [7:0] data_byte_6 = data[119:112]; // @[matcher.scala 326:37]
  wire  key_equal_6 = 8'h6 < _GEN_6 ? key_byte_6 == data_byte_6 : 1'h1; // @[matcher.scala 327:90 matcher.scala 328:34 matcher.scala 330:34]
  wire [7:0] key_byte_7 = key[63:56]; // @[matcher.scala 325:35]
  wire [7:0] data_byte_7 = data[127:120]; // @[matcher.scala 326:37]
  wire  key_equal_7 = 8'h7 < _GEN_6 ? key_byte_7 == data_byte_7 : 1'h1; // @[matcher.scala 327:90 matcher.scala 328:34 matcher.scala 330:34]
  wire [7:0] key_byte_8 = key[71:64]; // @[matcher.scala 325:35]
  wire [7:0] data_byte_8 = data[135:128]; // @[matcher.scala 326:37]
  wire  key_equal_8 = 8'h8 < _GEN_6 ? key_byte_8 == data_byte_8 : 1'h1; // @[matcher.scala 327:90 matcher.scala 328:34 matcher.scala 330:34]
  wire [7:0] key_byte_9 = key[79:72]; // @[matcher.scala 325:35]
  wire [7:0] data_byte_9 = data[143:136]; // @[matcher.scala 326:37]
  wire  key_equal_9 = 8'h9 < _GEN_6 ? key_byte_9 == data_byte_9 : 1'h1; // @[matcher.scala 327:90 matcher.scala 328:34 matcher.scala 330:34]
  wire [7:0] key_byte_10 = key[87:80]; // @[matcher.scala 325:35]
  wire [7:0] data_byte_10 = data[151:144]; // @[matcher.scala 326:37]
  wire  key_equal_10 = 8'ha < _GEN_6 ? key_byte_10 == data_byte_10 : 1'h1; // @[matcher.scala 327:90 matcher.scala 328:34 matcher.scala 330:34]
  wire [7:0] key_byte_11 = key[95:88]; // @[matcher.scala 325:35]
  wire [7:0] data_byte_11 = data[159:152]; // @[matcher.scala 326:37]
  wire  key_equal_11 = 8'hb < _GEN_6 ? key_byte_11 == data_byte_11 : 1'h1; // @[matcher.scala 327:90 matcher.scala 328:34 matcher.scala 330:34]
  wire [7:0] key_byte_12 = key[103:96]; // @[matcher.scala 325:35]
  wire [7:0] data_byte_12 = data[167:160]; // @[matcher.scala 326:37]
  wire  key_equal_12 = 8'hc < _GEN_6 ? key_byte_12 == data_byte_12 : 1'h1; // @[matcher.scala 327:90 matcher.scala 328:34 matcher.scala 330:34]
  wire [7:0] key_byte_13 = key[111:104]; // @[matcher.scala 325:35]
  wire [7:0] data_byte_13 = data[175:168]; // @[matcher.scala 326:37]
  wire  key_equal_13 = 8'hd < _GEN_6 ? key_byte_13 == data_byte_13 : 1'h1; // @[matcher.scala 327:90 matcher.scala 328:34 matcher.scala 330:34]
  wire [7:0] key_byte_14 = key[119:112]; // @[matcher.scala 325:35]
  wire [7:0] data_byte_14 = data[183:176]; // @[matcher.scala 326:37]
  wire  key_equal_14 = 8'he < _GEN_6 ? key_byte_14 == data_byte_14 : 1'h1; // @[matcher.scala 327:90 matcher.scala 328:34 matcher.scala 330:34]
  wire [7:0] key_byte_15 = key[127:120]; // @[matcher.scala 325:35]
  wire [7:0] data_byte_15 = data[191:184]; // @[matcher.scala 326:37]
  wire  key_equal_15 = 8'hf < _GEN_6 ? key_byte_15 == data_byte_15 : 1'h1; // @[matcher.scala 327:90 matcher.scala 328:34 matcher.scala 330:34]
  wire [7:0] key_byte_16 = key[135:128]; // @[matcher.scala 325:35]
  wire [7:0] data_byte_16 = data[199:192]; // @[matcher.scala 326:37]
  wire  key_equal_16 = 8'h10 < _GEN_6 ? key_byte_16 == data_byte_16 : 1'h1; // @[matcher.scala 327:90 matcher.scala 328:34 matcher.scala 330:34]
  wire [7:0] key_byte_17 = key[143:136]; // @[matcher.scala 325:35]
  wire [7:0] data_byte_17 = data[207:200]; // @[matcher.scala 326:37]
  wire  key_equal_17 = 8'h11 < _GEN_6 ? key_byte_17 == data_byte_17 : 1'h1; // @[matcher.scala 327:90 matcher.scala 328:34 matcher.scala 330:34]
  wire [7:0] key_byte_18 = key[151:144]; // @[matcher.scala 325:35]
  wire [7:0] data_byte_18 = data[215:208]; // @[matcher.scala 326:37]
  wire  key_equal_18 = 8'h12 < _GEN_6 ? key_byte_18 == data_byte_18 : 1'h1; // @[matcher.scala 327:90 matcher.scala 328:34 matcher.scala 330:34]
  wire [7:0] key_byte_19 = key[159:152]; // @[matcher.scala 325:35]
  wire [7:0] data_byte_19 = data[223:216]; // @[matcher.scala 326:37]
  wire  key_equal_19 = 8'h13 < _GEN_6 ? key_byte_19 == data_byte_19 : 1'h1; // @[matcher.scala 327:90 matcher.scala 328:34 matcher.scala 330:34]
  wire [7:0] key_byte_20 = key[167:160]; // @[matcher.scala 325:35]
  wire [7:0] data_byte_20 = data[231:224]; // @[matcher.scala 326:37]
  wire  key_equal_20 = 8'h14 < _GEN_6 ? key_byte_20 == data_byte_20 : 1'h1; // @[matcher.scala 327:90 matcher.scala 328:34 matcher.scala 330:34]
  wire [7:0] key_byte_21 = key[175:168]; // @[matcher.scala 325:35]
  wire [7:0] data_byte_21 = data[239:232]; // @[matcher.scala 326:37]
  wire  key_equal_21 = 8'h15 < _GEN_6 ? key_byte_21 == data_byte_21 : 1'h1; // @[matcher.scala 327:90 matcher.scala 328:34 matcher.scala 330:34]
  wire [7:0] key_byte_22 = key[183:176]; // @[matcher.scala 325:35]
  wire [7:0] data_byte_22 = data[247:240]; // @[matcher.scala 326:37]
  wire  key_equal_22 = 8'h16 < _GEN_6 ? key_byte_22 == data_byte_22 : 1'h1; // @[matcher.scala 327:90 matcher.scala 328:34 matcher.scala 330:34]
  wire [7:0] key_byte_23 = key[191:184]; // @[matcher.scala 325:35]
  wire [7:0] data_byte_23 = data[255:248]; // @[matcher.scala 326:37]
  wire  key_equal_23 = 8'h17 < _GEN_6 ? key_byte_23 == data_byte_23 : 1'h1; // @[matcher.scala 327:90 matcher.scala 328:34 matcher.scala 330:34]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_96 = phv_data_96; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_97 = phv_data_97; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_98 = phv_data_98; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_99 = phv_data_99; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_100 = phv_data_100; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_101 = phv_data_101; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_102 = phv_data_102; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_103 = phv_data_103; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_104 = phv_data_104; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_105 = phv_data_105; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_106 = phv_data_106; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_107 = phv_data_107; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_108 = phv_data_108; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_109 = phv_data_109; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_110 = phv_data_110; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_111 = phv_data_111; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_112 = phv_data_112; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_113 = phv_data_113; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_114 = phv_data_114; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_115 = phv_data_115; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_116 = phv_data_116; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_117 = phv_data_117; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_118 = phv_data_118; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_119 = phv_data_119; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_120 = phv_data_120; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_121 = phv_data_121; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_122 = phv_data_122; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_123 = phv_data_123; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_124 = phv_data_124; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_125 = phv_data_125; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_126 = phv_data_126; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_127 = phv_data_127; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_128 = phv_data_128; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_129 = phv_data_129; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_130 = phv_data_130; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_131 = phv_data_131; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_132 = phv_data_132; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_133 = phv_data_133; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_134 = phv_data_134; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_135 = phv_data_135; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_136 = phv_data_136; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_137 = phv_data_137; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_138 = phv_data_138; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_139 = phv_data_139; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_140 = phv_data_140; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_141 = phv_data_141; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_142 = phv_data_142; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_143 = phv_data_143; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_144 = phv_data_144; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_145 = phv_data_145; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_146 = phv_data_146; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_147 = phv_data_147; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_148 = phv_data_148; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_149 = phv_data_149; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_150 = phv_data_150; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_151 = phv_data_151; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_152 = phv_data_152; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_153 = phv_data_153; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_154 = phv_data_154; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_155 = phv_data_155; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_156 = phv_data_156; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_157 = phv_data_157; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_158 = phv_data_158; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_159 = phv_data_159; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_160 = phv_data_160; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_161 = phv_data_161; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_162 = phv_data_162; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_163 = phv_data_163; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_164 = phv_data_164; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_165 = phv_data_165; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_166 = phv_data_166; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_167 = phv_data_167; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_168 = phv_data_168; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_169 = phv_data_169; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_170 = phv_data_170; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_171 = phv_data_171; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_172 = phv_data_172; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_173 = phv_data_173; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_174 = phv_data_174; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_175 = phv_data_175; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_176 = phv_data_176; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_177 = phv_data_177; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_178 = phv_data_178; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_179 = phv_data_179; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_180 = phv_data_180; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_181 = phv_data_181; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_182 = phv_data_182; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_183 = phv_data_183; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_184 = phv_data_184; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_185 = phv_data_185; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_186 = phv_data_186; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_187 = phv_data_187; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_188 = phv_data_188; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_189 = phv_data_189; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_190 = phv_data_190; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_191 = phv_data_191; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_192 = phv_data_192; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_193 = phv_data_193; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_194 = phv_data_194; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_195 = phv_data_195; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_196 = phv_data_196; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_197 = phv_data_197; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_198 = phv_data_198; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_199 = phv_data_199; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_200 = phv_data_200; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_201 = phv_data_201; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_202 = phv_data_202; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_203 = phv_data_203; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_204 = phv_data_204; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_205 = phv_data_205; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_206 = phv_data_206; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_207 = phv_data_207; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_208 = phv_data_208; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_209 = phv_data_209; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_210 = phv_data_210; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_211 = phv_data_211; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_212 = phv_data_212; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_213 = phv_data_213; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_214 = phv_data_214; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_215 = phv_data_215; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_216 = phv_data_216; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_217 = phv_data_217; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_218 = phv_data_218; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_219 = phv_data_219; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_220 = phv_data_220; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_221 = phv_data_221; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_222 = phv_data_222; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_223 = phv_data_223; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_224 = phv_data_224; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_225 = phv_data_225; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_226 = phv_data_226; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_227 = phv_data_227; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_228 = phv_data_228; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_229 = phv_data_229; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_230 = phv_data_230; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_231 = phv_data_231; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_232 = phv_data_232; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_233 = phv_data_233; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_234 = phv_data_234; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_235 = phv_data_235; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_236 = phv_data_236; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_237 = phv_data_237; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_238 = phv_data_238; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_239 = phv_data_239; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_240 = phv_data_240; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_241 = phv_data_241; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_242 = phv_data_242; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_243 = phv_data_243; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_244 = phv_data_244; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_245 = phv_data_245; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_246 = phv_data_246; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_247 = phv_data_247; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_248 = phv_data_248; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_249 = phv_data_249; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_250 = phv_data_250; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_251 = phv_data_251; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_252 = phv_data_252; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_253 = phv_data_253; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_254 = phv_data_254; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_data_255 = phv_data_255; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[matcher.scala 313:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[matcher.scala 313:25]
  assign io_hit = phv_is_valid_processor & (key_equal_0 & key_equal_1 & key_equal_2 & key_equal_3 & key_equal_4 &
    key_equal_5 & key_equal_6 & key_equal_7 & key_equal_8 & key_equal_9 & key_equal_10 & key_equal_11 & key_equal_12 &
    key_equal_13 & key_equal_14 & key_equal_15 & key_equal_16 & key_equal_17 & key_equal_18 & key_equal_19 &
    key_equal_20 & key_equal_21 & key_equal_22 & key_equal_23); // @[matcher.scala 320:39 matcher.scala 334:20 matcher.scala 337:20]
  assign io_match_value = phv_is_valid_processor ? data[63:0] : 64'h0; // @[matcher.scala 320:39 matcher.scala 335:28 matcher.scala 338:28]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[matcher.scala 312:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[matcher.scala 312:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[matcher.scala 312:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[matcher.scala 312:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[matcher.scala 312:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[matcher.scala 312:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[matcher.scala 312:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[matcher.scala 312:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[matcher.scala 312:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[matcher.scala 312:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[matcher.scala 312:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[matcher.scala 312:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[matcher.scala 312:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[matcher.scala 312:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[matcher.scala 312:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[matcher.scala 312:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[matcher.scala 312:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[matcher.scala 312:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[matcher.scala 312:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[matcher.scala 312:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[matcher.scala 312:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[matcher.scala 312:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[matcher.scala 312:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[matcher.scala 312:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[matcher.scala 312:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[matcher.scala 312:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[matcher.scala 312:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[matcher.scala 312:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[matcher.scala 312:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[matcher.scala 312:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[matcher.scala 312:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[matcher.scala 312:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[matcher.scala 312:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[matcher.scala 312:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[matcher.scala 312:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[matcher.scala 312:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[matcher.scala 312:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[matcher.scala 312:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[matcher.scala 312:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[matcher.scala 312:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[matcher.scala 312:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[matcher.scala 312:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[matcher.scala 312:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[matcher.scala 312:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[matcher.scala 312:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[matcher.scala 312:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[matcher.scala 312:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[matcher.scala 312:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[matcher.scala 312:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[matcher.scala 312:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[matcher.scala 312:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[matcher.scala 312:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[matcher.scala 312:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[matcher.scala 312:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[matcher.scala 312:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[matcher.scala 312:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[matcher.scala 312:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[matcher.scala 312:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[matcher.scala 312:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[matcher.scala 312:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[matcher.scala 312:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[matcher.scala 312:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[matcher.scala 312:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[matcher.scala 312:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[matcher.scala 312:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[matcher.scala 312:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[matcher.scala 312:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[matcher.scala 312:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[matcher.scala 312:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[matcher.scala 312:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[matcher.scala 312:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[matcher.scala 312:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[matcher.scala 312:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[matcher.scala 312:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[matcher.scala 312:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[matcher.scala 312:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[matcher.scala 312:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[matcher.scala 312:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[matcher.scala 312:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[matcher.scala 312:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[matcher.scala 312:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[matcher.scala 312:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[matcher.scala 312:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[matcher.scala 312:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[matcher.scala 312:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[matcher.scala 312:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[matcher.scala 312:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[matcher.scala 312:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[matcher.scala 312:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[matcher.scala 312:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[matcher.scala 312:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[matcher.scala 312:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[matcher.scala 312:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[matcher.scala 312:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[matcher.scala 312:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[matcher.scala 312:13]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[matcher.scala 312:13]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[matcher.scala 312:13]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[matcher.scala 312:13]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[matcher.scala 312:13]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[matcher.scala 312:13]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[matcher.scala 312:13]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[matcher.scala 312:13]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[matcher.scala 312:13]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[matcher.scala 312:13]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[matcher.scala 312:13]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[matcher.scala 312:13]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[matcher.scala 312:13]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[matcher.scala 312:13]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[matcher.scala 312:13]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[matcher.scala 312:13]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[matcher.scala 312:13]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[matcher.scala 312:13]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[matcher.scala 312:13]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[matcher.scala 312:13]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[matcher.scala 312:13]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[matcher.scala 312:13]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[matcher.scala 312:13]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[matcher.scala 312:13]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[matcher.scala 312:13]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[matcher.scala 312:13]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[matcher.scala 312:13]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[matcher.scala 312:13]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[matcher.scala 312:13]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[matcher.scala 312:13]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[matcher.scala 312:13]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[matcher.scala 312:13]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[matcher.scala 312:13]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[matcher.scala 312:13]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[matcher.scala 312:13]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[matcher.scala 312:13]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[matcher.scala 312:13]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[matcher.scala 312:13]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[matcher.scala 312:13]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[matcher.scala 312:13]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[matcher.scala 312:13]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[matcher.scala 312:13]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[matcher.scala 312:13]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[matcher.scala 312:13]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[matcher.scala 312:13]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[matcher.scala 312:13]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[matcher.scala 312:13]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[matcher.scala 312:13]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[matcher.scala 312:13]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[matcher.scala 312:13]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[matcher.scala 312:13]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[matcher.scala 312:13]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[matcher.scala 312:13]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[matcher.scala 312:13]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[matcher.scala 312:13]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[matcher.scala 312:13]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[matcher.scala 312:13]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[matcher.scala 312:13]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[matcher.scala 312:13]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[matcher.scala 312:13]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[matcher.scala 312:13]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[matcher.scala 312:13]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[matcher.scala 312:13]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[matcher.scala 312:13]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[matcher.scala 312:13]
    phv_data_160 <= io_pipe_phv_in_data_160; // @[matcher.scala 312:13]
    phv_data_161 <= io_pipe_phv_in_data_161; // @[matcher.scala 312:13]
    phv_data_162 <= io_pipe_phv_in_data_162; // @[matcher.scala 312:13]
    phv_data_163 <= io_pipe_phv_in_data_163; // @[matcher.scala 312:13]
    phv_data_164 <= io_pipe_phv_in_data_164; // @[matcher.scala 312:13]
    phv_data_165 <= io_pipe_phv_in_data_165; // @[matcher.scala 312:13]
    phv_data_166 <= io_pipe_phv_in_data_166; // @[matcher.scala 312:13]
    phv_data_167 <= io_pipe_phv_in_data_167; // @[matcher.scala 312:13]
    phv_data_168 <= io_pipe_phv_in_data_168; // @[matcher.scala 312:13]
    phv_data_169 <= io_pipe_phv_in_data_169; // @[matcher.scala 312:13]
    phv_data_170 <= io_pipe_phv_in_data_170; // @[matcher.scala 312:13]
    phv_data_171 <= io_pipe_phv_in_data_171; // @[matcher.scala 312:13]
    phv_data_172 <= io_pipe_phv_in_data_172; // @[matcher.scala 312:13]
    phv_data_173 <= io_pipe_phv_in_data_173; // @[matcher.scala 312:13]
    phv_data_174 <= io_pipe_phv_in_data_174; // @[matcher.scala 312:13]
    phv_data_175 <= io_pipe_phv_in_data_175; // @[matcher.scala 312:13]
    phv_data_176 <= io_pipe_phv_in_data_176; // @[matcher.scala 312:13]
    phv_data_177 <= io_pipe_phv_in_data_177; // @[matcher.scala 312:13]
    phv_data_178 <= io_pipe_phv_in_data_178; // @[matcher.scala 312:13]
    phv_data_179 <= io_pipe_phv_in_data_179; // @[matcher.scala 312:13]
    phv_data_180 <= io_pipe_phv_in_data_180; // @[matcher.scala 312:13]
    phv_data_181 <= io_pipe_phv_in_data_181; // @[matcher.scala 312:13]
    phv_data_182 <= io_pipe_phv_in_data_182; // @[matcher.scala 312:13]
    phv_data_183 <= io_pipe_phv_in_data_183; // @[matcher.scala 312:13]
    phv_data_184 <= io_pipe_phv_in_data_184; // @[matcher.scala 312:13]
    phv_data_185 <= io_pipe_phv_in_data_185; // @[matcher.scala 312:13]
    phv_data_186 <= io_pipe_phv_in_data_186; // @[matcher.scala 312:13]
    phv_data_187 <= io_pipe_phv_in_data_187; // @[matcher.scala 312:13]
    phv_data_188 <= io_pipe_phv_in_data_188; // @[matcher.scala 312:13]
    phv_data_189 <= io_pipe_phv_in_data_189; // @[matcher.scala 312:13]
    phv_data_190 <= io_pipe_phv_in_data_190; // @[matcher.scala 312:13]
    phv_data_191 <= io_pipe_phv_in_data_191; // @[matcher.scala 312:13]
    phv_data_192 <= io_pipe_phv_in_data_192; // @[matcher.scala 312:13]
    phv_data_193 <= io_pipe_phv_in_data_193; // @[matcher.scala 312:13]
    phv_data_194 <= io_pipe_phv_in_data_194; // @[matcher.scala 312:13]
    phv_data_195 <= io_pipe_phv_in_data_195; // @[matcher.scala 312:13]
    phv_data_196 <= io_pipe_phv_in_data_196; // @[matcher.scala 312:13]
    phv_data_197 <= io_pipe_phv_in_data_197; // @[matcher.scala 312:13]
    phv_data_198 <= io_pipe_phv_in_data_198; // @[matcher.scala 312:13]
    phv_data_199 <= io_pipe_phv_in_data_199; // @[matcher.scala 312:13]
    phv_data_200 <= io_pipe_phv_in_data_200; // @[matcher.scala 312:13]
    phv_data_201 <= io_pipe_phv_in_data_201; // @[matcher.scala 312:13]
    phv_data_202 <= io_pipe_phv_in_data_202; // @[matcher.scala 312:13]
    phv_data_203 <= io_pipe_phv_in_data_203; // @[matcher.scala 312:13]
    phv_data_204 <= io_pipe_phv_in_data_204; // @[matcher.scala 312:13]
    phv_data_205 <= io_pipe_phv_in_data_205; // @[matcher.scala 312:13]
    phv_data_206 <= io_pipe_phv_in_data_206; // @[matcher.scala 312:13]
    phv_data_207 <= io_pipe_phv_in_data_207; // @[matcher.scala 312:13]
    phv_data_208 <= io_pipe_phv_in_data_208; // @[matcher.scala 312:13]
    phv_data_209 <= io_pipe_phv_in_data_209; // @[matcher.scala 312:13]
    phv_data_210 <= io_pipe_phv_in_data_210; // @[matcher.scala 312:13]
    phv_data_211 <= io_pipe_phv_in_data_211; // @[matcher.scala 312:13]
    phv_data_212 <= io_pipe_phv_in_data_212; // @[matcher.scala 312:13]
    phv_data_213 <= io_pipe_phv_in_data_213; // @[matcher.scala 312:13]
    phv_data_214 <= io_pipe_phv_in_data_214; // @[matcher.scala 312:13]
    phv_data_215 <= io_pipe_phv_in_data_215; // @[matcher.scala 312:13]
    phv_data_216 <= io_pipe_phv_in_data_216; // @[matcher.scala 312:13]
    phv_data_217 <= io_pipe_phv_in_data_217; // @[matcher.scala 312:13]
    phv_data_218 <= io_pipe_phv_in_data_218; // @[matcher.scala 312:13]
    phv_data_219 <= io_pipe_phv_in_data_219; // @[matcher.scala 312:13]
    phv_data_220 <= io_pipe_phv_in_data_220; // @[matcher.scala 312:13]
    phv_data_221 <= io_pipe_phv_in_data_221; // @[matcher.scala 312:13]
    phv_data_222 <= io_pipe_phv_in_data_222; // @[matcher.scala 312:13]
    phv_data_223 <= io_pipe_phv_in_data_223; // @[matcher.scala 312:13]
    phv_data_224 <= io_pipe_phv_in_data_224; // @[matcher.scala 312:13]
    phv_data_225 <= io_pipe_phv_in_data_225; // @[matcher.scala 312:13]
    phv_data_226 <= io_pipe_phv_in_data_226; // @[matcher.scala 312:13]
    phv_data_227 <= io_pipe_phv_in_data_227; // @[matcher.scala 312:13]
    phv_data_228 <= io_pipe_phv_in_data_228; // @[matcher.scala 312:13]
    phv_data_229 <= io_pipe_phv_in_data_229; // @[matcher.scala 312:13]
    phv_data_230 <= io_pipe_phv_in_data_230; // @[matcher.scala 312:13]
    phv_data_231 <= io_pipe_phv_in_data_231; // @[matcher.scala 312:13]
    phv_data_232 <= io_pipe_phv_in_data_232; // @[matcher.scala 312:13]
    phv_data_233 <= io_pipe_phv_in_data_233; // @[matcher.scala 312:13]
    phv_data_234 <= io_pipe_phv_in_data_234; // @[matcher.scala 312:13]
    phv_data_235 <= io_pipe_phv_in_data_235; // @[matcher.scala 312:13]
    phv_data_236 <= io_pipe_phv_in_data_236; // @[matcher.scala 312:13]
    phv_data_237 <= io_pipe_phv_in_data_237; // @[matcher.scala 312:13]
    phv_data_238 <= io_pipe_phv_in_data_238; // @[matcher.scala 312:13]
    phv_data_239 <= io_pipe_phv_in_data_239; // @[matcher.scala 312:13]
    phv_data_240 <= io_pipe_phv_in_data_240; // @[matcher.scala 312:13]
    phv_data_241 <= io_pipe_phv_in_data_241; // @[matcher.scala 312:13]
    phv_data_242 <= io_pipe_phv_in_data_242; // @[matcher.scala 312:13]
    phv_data_243 <= io_pipe_phv_in_data_243; // @[matcher.scala 312:13]
    phv_data_244 <= io_pipe_phv_in_data_244; // @[matcher.scala 312:13]
    phv_data_245 <= io_pipe_phv_in_data_245; // @[matcher.scala 312:13]
    phv_data_246 <= io_pipe_phv_in_data_246; // @[matcher.scala 312:13]
    phv_data_247 <= io_pipe_phv_in_data_247; // @[matcher.scala 312:13]
    phv_data_248 <= io_pipe_phv_in_data_248; // @[matcher.scala 312:13]
    phv_data_249 <= io_pipe_phv_in_data_249; // @[matcher.scala 312:13]
    phv_data_250 <= io_pipe_phv_in_data_250; // @[matcher.scala 312:13]
    phv_data_251 <= io_pipe_phv_in_data_251; // @[matcher.scala 312:13]
    phv_data_252 <= io_pipe_phv_in_data_252; // @[matcher.scala 312:13]
    phv_data_253 <= io_pipe_phv_in_data_253; // @[matcher.scala 312:13]
    phv_data_254 <= io_pipe_phv_in_data_254; // @[matcher.scala 312:13]
    phv_data_255 <= io_pipe_phv_in_data_255; // @[matcher.scala 312:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[matcher.scala 312:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[matcher.scala 312:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[matcher.scala 312:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[matcher.scala 312:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[matcher.scala 312:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[matcher.scala 312:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[matcher.scala 312:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[matcher.scala 312:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[matcher.scala 312:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[matcher.scala 312:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[matcher.scala 312:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[matcher.scala 312:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[matcher.scala 312:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[matcher.scala 312:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[matcher.scala 312:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[matcher.scala 312:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[matcher.scala 312:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[matcher.scala 312:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[matcher.scala 312:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[matcher.scala 312:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[matcher.scala 312:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[matcher.scala 312:13]
    key <= io_key_in; // @[matcher.scala 316:13]
    data <= io_data_in; // @[matcher.scala 318:14]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_data_160 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  phv_data_161 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  phv_data_162 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  phv_data_163 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  phv_data_164 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  phv_data_165 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  phv_data_166 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  phv_data_167 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  phv_data_168 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  phv_data_169 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  phv_data_170 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  phv_data_171 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  phv_data_172 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  phv_data_173 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  phv_data_174 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  phv_data_175 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  phv_data_176 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_data_177 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_data_178 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  phv_data_179 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  phv_data_180 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  phv_data_181 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  phv_data_182 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  phv_data_183 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  phv_data_184 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  phv_data_185 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  phv_data_186 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  phv_data_187 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  phv_data_188 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  phv_data_189 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  phv_data_190 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  phv_data_191 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  phv_data_192 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  phv_data_193 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  phv_data_194 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  phv_data_195 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  phv_data_196 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  phv_data_197 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  phv_data_198 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  phv_data_199 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  phv_data_200 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  phv_data_201 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  phv_data_202 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  phv_data_203 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  phv_data_204 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  phv_data_205 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  phv_data_206 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  phv_data_207 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  phv_data_208 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  phv_data_209 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  phv_data_210 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  phv_data_211 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  phv_data_212 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  phv_data_213 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  phv_data_214 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  phv_data_215 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  phv_data_216 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  phv_data_217 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  phv_data_218 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  phv_data_219 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  phv_data_220 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  phv_data_221 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  phv_data_222 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  phv_data_223 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  phv_data_224 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  phv_data_225 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  phv_data_226 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  phv_data_227 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  phv_data_228 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  phv_data_229 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  phv_data_230 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  phv_data_231 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  phv_data_232 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  phv_data_233 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  phv_data_234 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  phv_data_235 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  phv_data_236 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  phv_data_237 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  phv_data_238 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  phv_data_239 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  phv_data_240 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  phv_data_241 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  phv_data_242 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  phv_data_243 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  phv_data_244 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  phv_data_245 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  phv_data_246 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  phv_data_247 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  phv_data_248 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  phv_data_249 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  phv_data_250 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  phv_data_251 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  phv_data_252 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  phv_data_253 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  phv_data_254 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  phv_data_255 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  phv_header_0 = _RAND_256[15:0];
  _RAND_257 = {1{`RANDOM}};
  phv_header_1 = _RAND_257[15:0];
  _RAND_258 = {1{`RANDOM}};
  phv_header_2 = _RAND_258[15:0];
  _RAND_259 = {1{`RANDOM}};
  phv_header_3 = _RAND_259[15:0];
  _RAND_260 = {1{`RANDOM}};
  phv_header_4 = _RAND_260[15:0];
  _RAND_261 = {1{`RANDOM}};
  phv_header_5 = _RAND_261[15:0];
  _RAND_262 = {1{`RANDOM}};
  phv_header_6 = _RAND_262[15:0];
  _RAND_263 = {1{`RANDOM}};
  phv_header_7 = _RAND_263[15:0];
  _RAND_264 = {1{`RANDOM}};
  phv_header_8 = _RAND_264[15:0];
  _RAND_265 = {1{`RANDOM}};
  phv_header_9 = _RAND_265[15:0];
  _RAND_266 = {1{`RANDOM}};
  phv_header_10 = _RAND_266[15:0];
  _RAND_267 = {1{`RANDOM}};
  phv_header_11 = _RAND_267[15:0];
  _RAND_268 = {1{`RANDOM}};
  phv_header_12 = _RAND_268[15:0];
  _RAND_269 = {1{`RANDOM}};
  phv_header_13 = _RAND_269[15:0];
  _RAND_270 = {1{`RANDOM}};
  phv_header_14 = _RAND_270[15:0];
  _RAND_271 = {1{`RANDOM}};
  phv_header_15 = _RAND_271[15:0];
  _RAND_272 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_272[7:0];
  _RAND_273 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_273[7:0];
  _RAND_274 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_274[15:0];
  _RAND_275 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_275[2:0];
  _RAND_276 = {1{`RANDOM}};
  phv_next_config_id = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_277[0:0];
  _RAND_278 = {6{`RANDOM}};
  key = _RAND_278[191:0];
  _RAND_279 = {8{`RANDOM}};
  data = _RAND_279[255:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
