module PrimitiveGetSourcePISA(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [7:0]  io_pipe_phv_in_data_160,
  input  [7:0]  io_pipe_phv_in_data_161,
  input  [7:0]  io_pipe_phv_in_data_162,
  input  [7:0]  io_pipe_phv_in_data_163,
  input  [7:0]  io_pipe_phv_in_data_164,
  input  [7:0]  io_pipe_phv_in_data_165,
  input  [7:0]  io_pipe_phv_in_data_166,
  input  [7:0]  io_pipe_phv_in_data_167,
  input  [7:0]  io_pipe_phv_in_data_168,
  input  [7:0]  io_pipe_phv_in_data_169,
  input  [7:0]  io_pipe_phv_in_data_170,
  input  [7:0]  io_pipe_phv_in_data_171,
  input  [7:0]  io_pipe_phv_in_data_172,
  input  [7:0]  io_pipe_phv_in_data_173,
  input  [7:0]  io_pipe_phv_in_data_174,
  input  [7:0]  io_pipe_phv_in_data_175,
  input  [7:0]  io_pipe_phv_in_data_176,
  input  [7:0]  io_pipe_phv_in_data_177,
  input  [7:0]  io_pipe_phv_in_data_178,
  input  [7:0]  io_pipe_phv_in_data_179,
  input  [7:0]  io_pipe_phv_in_data_180,
  input  [7:0]  io_pipe_phv_in_data_181,
  input  [7:0]  io_pipe_phv_in_data_182,
  input  [7:0]  io_pipe_phv_in_data_183,
  input  [7:0]  io_pipe_phv_in_data_184,
  input  [7:0]  io_pipe_phv_in_data_185,
  input  [7:0]  io_pipe_phv_in_data_186,
  input  [7:0]  io_pipe_phv_in_data_187,
  input  [7:0]  io_pipe_phv_in_data_188,
  input  [7:0]  io_pipe_phv_in_data_189,
  input  [7:0]  io_pipe_phv_in_data_190,
  input  [7:0]  io_pipe_phv_in_data_191,
  input  [7:0]  io_pipe_phv_in_data_192,
  input  [7:0]  io_pipe_phv_in_data_193,
  input  [7:0]  io_pipe_phv_in_data_194,
  input  [7:0]  io_pipe_phv_in_data_195,
  input  [7:0]  io_pipe_phv_in_data_196,
  input  [7:0]  io_pipe_phv_in_data_197,
  input  [7:0]  io_pipe_phv_in_data_198,
  input  [7:0]  io_pipe_phv_in_data_199,
  input  [7:0]  io_pipe_phv_in_data_200,
  input  [7:0]  io_pipe_phv_in_data_201,
  input  [7:0]  io_pipe_phv_in_data_202,
  input  [7:0]  io_pipe_phv_in_data_203,
  input  [7:0]  io_pipe_phv_in_data_204,
  input  [7:0]  io_pipe_phv_in_data_205,
  input  [7:0]  io_pipe_phv_in_data_206,
  input  [7:0]  io_pipe_phv_in_data_207,
  input  [7:0]  io_pipe_phv_in_data_208,
  input  [7:0]  io_pipe_phv_in_data_209,
  input  [7:0]  io_pipe_phv_in_data_210,
  input  [7:0]  io_pipe_phv_in_data_211,
  input  [7:0]  io_pipe_phv_in_data_212,
  input  [7:0]  io_pipe_phv_in_data_213,
  input  [7:0]  io_pipe_phv_in_data_214,
  input  [7:0]  io_pipe_phv_in_data_215,
  input  [7:0]  io_pipe_phv_in_data_216,
  input  [7:0]  io_pipe_phv_in_data_217,
  input  [7:0]  io_pipe_phv_in_data_218,
  input  [7:0]  io_pipe_phv_in_data_219,
  input  [7:0]  io_pipe_phv_in_data_220,
  input  [7:0]  io_pipe_phv_in_data_221,
  input  [7:0]  io_pipe_phv_in_data_222,
  input  [7:0]  io_pipe_phv_in_data_223,
  input  [7:0]  io_pipe_phv_in_data_224,
  input  [7:0]  io_pipe_phv_in_data_225,
  input  [7:0]  io_pipe_phv_in_data_226,
  input  [7:0]  io_pipe_phv_in_data_227,
  input  [7:0]  io_pipe_phv_in_data_228,
  input  [7:0]  io_pipe_phv_in_data_229,
  input  [7:0]  io_pipe_phv_in_data_230,
  input  [7:0]  io_pipe_phv_in_data_231,
  input  [7:0]  io_pipe_phv_in_data_232,
  input  [7:0]  io_pipe_phv_in_data_233,
  input  [7:0]  io_pipe_phv_in_data_234,
  input  [7:0]  io_pipe_phv_in_data_235,
  input  [7:0]  io_pipe_phv_in_data_236,
  input  [7:0]  io_pipe_phv_in_data_237,
  input  [7:0]  io_pipe_phv_in_data_238,
  input  [7:0]  io_pipe_phv_in_data_239,
  input  [7:0]  io_pipe_phv_in_data_240,
  input  [7:0]  io_pipe_phv_in_data_241,
  input  [7:0]  io_pipe_phv_in_data_242,
  input  [7:0]  io_pipe_phv_in_data_243,
  input  [7:0]  io_pipe_phv_in_data_244,
  input  [7:0]  io_pipe_phv_in_data_245,
  input  [7:0]  io_pipe_phv_in_data_246,
  input  [7:0]  io_pipe_phv_in_data_247,
  input  [7:0]  io_pipe_phv_in_data_248,
  input  [7:0]  io_pipe_phv_in_data_249,
  input  [7:0]  io_pipe_phv_in_data_250,
  input  [7:0]  io_pipe_phv_in_data_251,
  input  [7:0]  io_pipe_phv_in_data_252,
  input  [7:0]  io_pipe_phv_in_data_253,
  input  [7:0]  io_pipe_phv_in_data_254,
  input  [7:0]  io_pipe_phv_in_data_255,
  input  [7:0]  io_pipe_phv_in_data_256,
  input  [7:0]  io_pipe_phv_in_data_257,
  input  [7:0]  io_pipe_phv_in_data_258,
  input  [7:0]  io_pipe_phv_in_data_259,
  input  [7:0]  io_pipe_phv_in_data_260,
  input  [7:0]  io_pipe_phv_in_data_261,
  input  [7:0]  io_pipe_phv_in_data_262,
  input  [7:0]  io_pipe_phv_in_data_263,
  input  [7:0]  io_pipe_phv_in_data_264,
  input  [7:0]  io_pipe_phv_in_data_265,
  input  [7:0]  io_pipe_phv_in_data_266,
  input  [7:0]  io_pipe_phv_in_data_267,
  input  [7:0]  io_pipe_phv_in_data_268,
  input  [7:0]  io_pipe_phv_in_data_269,
  input  [7:0]  io_pipe_phv_in_data_270,
  input  [7:0]  io_pipe_phv_in_data_271,
  input  [7:0]  io_pipe_phv_in_data_272,
  input  [7:0]  io_pipe_phv_in_data_273,
  input  [7:0]  io_pipe_phv_in_data_274,
  input  [7:0]  io_pipe_phv_in_data_275,
  input  [7:0]  io_pipe_phv_in_data_276,
  input  [7:0]  io_pipe_phv_in_data_277,
  input  [7:0]  io_pipe_phv_in_data_278,
  input  [7:0]  io_pipe_phv_in_data_279,
  input  [7:0]  io_pipe_phv_in_data_280,
  input  [7:0]  io_pipe_phv_in_data_281,
  input  [7:0]  io_pipe_phv_in_data_282,
  input  [7:0]  io_pipe_phv_in_data_283,
  input  [7:0]  io_pipe_phv_in_data_284,
  input  [7:0]  io_pipe_phv_in_data_285,
  input  [7:0]  io_pipe_phv_in_data_286,
  input  [7:0]  io_pipe_phv_in_data_287,
  input  [7:0]  io_pipe_phv_in_data_288,
  input  [7:0]  io_pipe_phv_in_data_289,
  input  [7:0]  io_pipe_phv_in_data_290,
  input  [7:0]  io_pipe_phv_in_data_291,
  input  [7:0]  io_pipe_phv_in_data_292,
  input  [7:0]  io_pipe_phv_in_data_293,
  input  [7:0]  io_pipe_phv_in_data_294,
  input  [7:0]  io_pipe_phv_in_data_295,
  input  [7:0]  io_pipe_phv_in_data_296,
  input  [7:0]  io_pipe_phv_in_data_297,
  input  [7:0]  io_pipe_phv_in_data_298,
  input  [7:0]  io_pipe_phv_in_data_299,
  input  [7:0]  io_pipe_phv_in_data_300,
  input  [7:0]  io_pipe_phv_in_data_301,
  input  [7:0]  io_pipe_phv_in_data_302,
  input  [7:0]  io_pipe_phv_in_data_303,
  input  [7:0]  io_pipe_phv_in_data_304,
  input  [7:0]  io_pipe_phv_in_data_305,
  input  [7:0]  io_pipe_phv_in_data_306,
  input  [7:0]  io_pipe_phv_in_data_307,
  input  [7:0]  io_pipe_phv_in_data_308,
  input  [7:0]  io_pipe_phv_in_data_309,
  input  [7:0]  io_pipe_phv_in_data_310,
  input  [7:0]  io_pipe_phv_in_data_311,
  input  [7:0]  io_pipe_phv_in_data_312,
  input  [7:0]  io_pipe_phv_in_data_313,
  input  [7:0]  io_pipe_phv_in_data_314,
  input  [7:0]  io_pipe_phv_in_data_315,
  input  [7:0]  io_pipe_phv_in_data_316,
  input  [7:0]  io_pipe_phv_in_data_317,
  input  [7:0]  io_pipe_phv_in_data_318,
  input  [7:0]  io_pipe_phv_in_data_319,
  input  [7:0]  io_pipe_phv_in_data_320,
  input  [7:0]  io_pipe_phv_in_data_321,
  input  [7:0]  io_pipe_phv_in_data_322,
  input  [7:0]  io_pipe_phv_in_data_323,
  input  [7:0]  io_pipe_phv_in_data_324,
  input  [7:0]  io_pipe_phv_in_data_325,
  input  [7:0]  io_pipe_phv_in_data_326,
  input  [7:0]  io_pipe_phv_in_data_327,
  input  [7:0]  io_pipe_phv_in_data_328,
  input  [7:0]  io_pipe_phv_in_data_329,
  input  [7:0]  io_pipe_phv_in_data_330,
  input  [7:0]  io_pipe_phv_in_data_331,
  input  [7:0]  io_pipe_phv_in_data_332,
  input  [7:0]  io_pipe_phv_in_data_333,
  input  [7:0]  io_pipe_phv_in_data_334,
  input  [7:0]  io_pipe_phv_in_data_335,
  input  [7:0]  io_pipe_phv_in_data_336,
  input  [7:0]  io_pipe_phv_in_data_337,
  input  [7:0]  io_pipe_phv_in_data_338,
  input  [7:0]  io_pipe_phv_in_data_339,
  input  [7:0]  io_pipe_phv_in_data_340,
  input  [7:0]  io_pipe_phv_in_data_341,
  input  [7:0]  io_pipe_phv_in_data_342,
  input  [7:0]  io_pipe_phv_in_data_343,
  input  [7:0]  io_pipe_phv_in_data_344,
  input  [7:0]  io_pipe_phv_in_data_345,
  input  [7:0]  io_pipe_phv_in_data_346,
  input  [7:0]  io_pipe_phv_in_data_347,
  input  [7:0]  io_pipe_phv_in_data_348,
  input  [7:0]  io_pipe_phv_in_data_349,
  input  [7:0]  io_pipe_phv_in_data_350,
  input  [7:0]  io_pipe_phv_in_data_351,
  input  [7:0]  io_pipe_phv_in_data_352,
  input  [7:0]  io_pipe_phv_in_data_353,
  input  [7:0]  io_pipe_phv_in_data_354,
  input  [7:0]  io_pipe_phv_in_data_355,
  input  [7:0]  io_pipe_phv_in_data_356,
  input  [7:0]  io_pipe_phv_in_data_357,
  input  [7:0]  io_pipe_phv_in_data_358,
  input  [7:0]  io_pipe_phv_in_data_359,
  input  [7:0]  io_pipe_phv_in_data_360,
  input  [7:0]  io_pipe_phv_in_data_361,
  input  [7:0]  io_pipe_phv_in_data_362,
  input  [7:0]  io_pipe_phv_in_data_363,
  input  [7:0]  io_pipe_phv_in_data_364,
  input  [7:0]  io_pipe_phv_in_data_365,
  input  [7:0]  io_pipe_phv_in_data_366,
  input  [7:0]  io_pipe_phv_in_data_367,
  input  [7:0]  io_pipe_phv_in_data_368,
  input  [7:0]  io_pipe_phv_in_data_369,
  input  [7:0]  io_pipe_phv_in_data_370,
  input  [7:0]  io_pipe_phv_in_data_371,
  input  [7:0]  io_pipe_phv_in_data_372,
  input  [7:0]  io_pipe_phv_in_data_373,
  input  [7:0]  io_pipe_phv_in_data_374,
  input  [7:0]  io_pipe_phv_in_data_375,
  input  [7:0]  io_pipe_phv_in_data_376,
  input  [7:0]  io_pipe_phv_in_data_377,
  input  [7:0]  io_pipe_phv_in_data_378,
  input  [7:0]  io_pipe_phv_in_data_379,
  input  [7:0]  io_pipe_phv_in_data_380,
  input  [7:0]  io_pipe_phv_in_data_381,
  input  [7:0]  io_pipe_phv_in_data_382,
  input  [7:0]  io_pipe_phv_in_data_383,
  input  [7:0]  io_pipe_phv_in_data_384,
  input  [7:0]  io_pipe_phv_in_data_385,
  input  [7:0]  io_pipe_phv_in_data_386,
  input  [7:0]  io_pipe_phv_in_data_387,
  input  [7:0]  io_pipe_phv_in_data_388,
  input  [7:0]  io_pipe_phv_in_data_389,
  input  [7:0]  io_pipe_phv_in_data_390,
  input  [7:0]  io_pipe_phv_in_data_391,
  input  [7:0]  io_pipe_phv_in_data_392,
  input  [7:0]  io_pipe_phv_in_data_393,
  input  [7:0]  io_pipe_phv_in_data_394,
  input  [7:0]  io_pipe_phv_in_data_395,
  input  [7:0]  io_pipe_phv_in_data_396,
  input  [7:0]  io_pipe_phv_in_data_397,
  input  [7:0]  io_pipe_phv_in_data_398,
  input  [7:0]  io_pipe_phv_in_data_399,
  input  [7:0]  io_pipe_phv_in_data_400,
  input  [7:0]  io_pipe_phv_in_data_401,
  input  [7:0]  io_pipe_phv_in_data_402,
  input  [7:0]  io_pipe_phv_in_data_403,
  input  [7:0]  io_pipe_phv_in_data_404,
  input  [7:0]  io_pipe_phv_in_data_405,
  input  [7:0]  io_pipe_phv_in_data_406,
  input  [7:0]  io_pipe_phv_in_data_407,
  input  [7:0]  io_pipe_phv_in_data_408,
  input  [7:0]  io_pipe_phv_in_data_409,
  input  [7:0]  io_pipe_phv_in_data_410,
  input  [7:0]  io_pipe_phv_in_data_411,
  input  [7:0]  io_pipe_phv_in_data_412,
  input  [7:0]  io_pipe_phv_in_data_413,
  input  [7:0]  io_pipe_phv_in_data_414,
  input  [7:0]  io_pipe_phv_in_data_415,
  input  [7:0]  io_pipe_phv_in_data_416,
  input  [7:0]  io_pipe_phv_in_data_417,
  input  [7:0]  io_pipe_phv_in_data_418,
  input  [7:0]  io_pipe_phv_in_data_419,
  input  [7:0]  io_pipe_phv_in_data_420,
  input  [7:0]  io_pipe_phv_in_data_421,
  input  [7:0]  io_pipe_phv_in_data_422,
  input  [7:0]  io_pipe_phv_in_data_423,
  input  [7:0]  io_pipe_phv_in_data_424,
  input  [7:0]  io_pipe_phv_in_data_425,
  input  [7:0]  io_pipe_phv_in_data_426,
  input  [7:0]  io_pipe_phv_in_data_427,
  input  [7:0]  io_pipe_phv_in_data_428,
  input  [7:0]  io_pipe_phv_in_data_429,
  input  [7:0]  io_pipe_phv_in_data_430,
  input  [7:0]  io_pipe_phv_in_data_431,
  input  [7:0]  io_pipe_phv_in_data_432,
  input  [7:0]  io_pipe_phv_in_data_433,
  input  [7:0]  io_pipe_phv_in_data_434,
  input  [7:0]  io_pipe_phv_in_data_435,
  input  [7:0]  io_pipe_phv_in_data_436,
  input  [7:0]  io_pipe_phv_in_data_437,
  input  [7:0]  io_pipe_phv_in_data_438,
  input  [7:0]  io_pipe_phv_in_data_439,
  input  [7:0]  io_pipe_phv_in_data_440,
  input  [7:0]  io_pipe_phv_in_data_441,
  input  [7:0]  io_pipe_phv_in_data_442,
  input  [7:0]  io_pipe_phv_in_data_443,
  input  [7:0]  io_pipe_phv_in_data_444,
  input  [7:0]  io_pipe_phv_in_data_445,
  input  [7:0]  io_pipe_phv_in_data_446,
  input  [7:0]  io_pipe_phv_in_data_447,
  input  [7:0]  io_pipe_phv_in_data_448,
  input  [7:0]  io_pipe_phv_in_data_449,
  input  [7:0]  io_pipe_phv_in_data_450,
  input  [7:0]  io_pipe_phv_in_data_451,
  input  [7:0]  io_pipe_phv_in_data_452,
  input  [7:0]  io_pipe_phv_in_data_453,
  input  [7:0]  io_pipe_phv_in_data_454,
  input  [7:0]  io_pipe_phv_in_data_455,
  input  [7:0]  io_pipe_phv_in_data_456,
  input  [7:0]  io_pipe_phv_in_data_457,
  input  [7:0]  io_pipe_phv_in_data_458,
  input  [7:0]  io_pipe_phv_in_data_459,
  input  [7:0]  io_pipe_phv_in_data_460,
  input  [7:0]  io_pipe_phv_in_data_461,
  input  [7:0]  io_pipe_phv_in_data_462,
  input  [7:0]  io_pipe_phv_in_data_463,
  input  [7:0]  io_pipe_phv_in_data_464,
  input  [7:0]  io_pipe_phv_in_data_465,
  input  [7:0]  io_pipe_phv_in_data_466,
  input  [7:0]  io_pipe_phv_in_data_467,
  input  [7:0]  io_pipe_phv_in_data_468,
  input  [7:0]  io_pipe_phv_in_data_469,
  input  [7:0]  io_pipe_phv_in_data_470,
  input  [7:0]  io_pipe_phv_in_data_471,
  input  [7:0]  io_pipe_phv_in_data_472,
  input  [7:0]  io_pipe_phv_in_data_473,
  input  [7:0]  io_pipe_phv_in_data_474,
  input  [7:0]  io_pipe_phv_in_data_475,
  input  [7:0]  io_pipe_phv_in_data_476,
  input  [7:0]  io_pipe_phv_in_data_477,
  input  [7:0]  io_pipe_phv_in_data_478,
  input  [7:0]  io_pipe_phv_in_data_479,
  input  [7:0]  io_pipe_phv_in_data_480,
  input  [7:0]  io_pipe_phv_in_data_481,
  input  [7:0]  io_pipe_phv_in_data_482,
  input  [7:0]  io_pipe_phv_in_data_483,
  input  [7:0]  io_pipe_phv_in_data_484,
  input  [7:0]  io_pipe_phv_in_data_485,
  input  [7:0]  io_pipe_phv_in_data_486,
  input  [7:0]  io_pipe_phv_in_data_487,
  input  [7:0]  io_pipe_phv_in_data_488,
  input  [7:0]  io_pipe_phv_in_data_489,
  input  [7:0]  io_pipe_phv_in_data_490,
  input  [7:0]  io_pipe_phv_in_data_491,
  input  [7:0]  io_pipe_phv_in_data_492,
  input  [7:0]  io_pipe_phv_in_data_493,
  input  [7:0]  io_pipe_phv_in_data_494,
  input  [7:0]  io_pipe_phv_in_data_495,
  input  [7:0]  io_pipe_phv_in_data_496,
  input  [7:0]  io_pipe_phv_in_data_497,
  input  [7:0]  io_pipe_phv_in_data_498,
  input  [7:0]  io_pipe_phv_in_data_499,
  input  [7:0]  io_pipe_phv_in_data_500,
  input  [7:0]  io_pipe_phv_in_data_501,
  input  [7:0]  io_pipe_phv_in_data_502,
  input  [7:0]  io_pipe_phv_in_data_503,
  input  [7:0]  io_pipe_phv_in_data_504,
  input  [7:0]  io_pipe_phv_in_data_505,
  input  [7:0]  io_pipe_phv_in_data_506,
  input  [7:0]  io_pipe_phv_in_data_507,
  input  [7:0]  io_pipe_phv_in_data_508,
  input  [7:0]  io_pipe_phv_in_data_509,
  input  [7:0]  io_pipe_phv_in_data_510,
  input  [7:0]  io_pipe_phv_in_data_511,
  input  [3:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [7:0]  io_pipe_phv_out_data_160,
  output [7:0]  io_pipe_phv_out_data_161,
  output [7:0]  io_pipe_phv_out_data_162,
  output [7:0]  io_pipe_phv_out_data_163,
  output [7:0]  io_pipe_phv_out_data_164,
  output [7:0]  io_pipe_phv_out_data_165,
  output [7:0]  io_pipe_phv_out_data_166,
  output [7:0]  io_pipe_phv_out_data_167,
  output [7:0]  io_pipe_phv_out_data_168,
  output [7:0]  io_pipe_phv_out_data_169,
  output [7:0]  io_pipe_phv_out_data_170,
  output [7:0]  io_pipe_phv_out_data_171,
  output [7:0]  io_pipe_phv_out_data_172,
  output [7:0]  io_pipe_phv_out_data_173,
  output [7:0]  io_pipe_phv_out_data_174,
  output [7:0]  io_pipe_phv_out_data_175,
  output [7:0]  io_pipe_phv_out_data_176,
  output [7:0]  io_pipe_phv_out_data_177,
  output [7:0]  io_pipe_phv_out_data_178,
  output [7:0]  io_pipe_phv_out_data_179,
  output [7:0]  io_pipe_phv_out_data_180,
  output [7:0]  io_pipe_phv_out_data_181,
  output [7:0]  io_pipe_phv_out_data_182,
  output [7:0]  io_pipe_phv_out_data_183,
  output [7:0]  io_pipe_phv_out_data_184,
  output [7:0]  io_pipe_phv_out_data_185,
  output [7:0]  io_pipe_phv_out_data_186,
  output [7:0]  io_pipe_phv_out_data_187,
  output [7:0]  io_pipe_phv_out_data_188,
  output [7:0]  io_pipe_phv_out_data_189,
  output [7:0]  io_pipe_phv_out_data_190,
  output [7:0]  io_pipe_phv_out_data_191,
  output [7:0]  io_pipe_phv_out_data_192,
  output [7:0]  io_pipe_phv_out_data_193,
  output [7:0]  io_pipe_phv_out_data_194,
  output [7:0]  io_pipe_phv_out_data_195,
  output [7:0]  io_pipe_phv_out_data_196,
  output [7:0]  io_pipe_phv_out_data_197,
  output [7:0]  io_pipe_phv_out_data_198,
  output [7:0]  io_pipe_phv_out_data_199,
  output [7:0]  io_pipe_phv_out_data_200,
  output [7:0]  io_pipe_phv_out_data_201,
  output [7:0]  io_pipe_phv_out_data_202,
  output [7:0]  io_pipe_phv_out_data_203,
  output [7:0]  io_pipe_phv_out_data_204,
  output [7:0]  io_pipe_phv_out_data_205,
  output [7:0]  io_pipe_phv_out_data_206,
  output [7:0]  io_pipe_phv_out_data_207,
  output [7:0]  io_pipe_phv_out_data_208,
  output [7:0]  io_pipe_phv_out_data_209,
  output [7:0]  io_pipe_phv_out_data_210,
  output [7:0]  io_pipe_phv_out_data_211,
  output [7:0]  io_pipe_phv_out_data_212,
  output [7:0]  io_pipe_phv_out_data_213,
  output [7:0]  io_pipe_phv_out_data_214,
  output [7:0]  io_pipe_phv_out_data_215,
  output [7:0]  io_pipe_phv_out_data_216,
  output [7:0]  io_pipe_phv_out_data_217,
  output [7:0]  io_pipe_phv_out_data_218,
  output [7:0]  io_pipe_phv_out_data_219,
  output [7:0]  io_pipe_phv_out_data_220,
  output [7:0]  io_pipe_phv_out_data_221,
  output [7:0]  io_pipe_phv_out_data_222,
  output [7:0]  io_pipe_phv_out_data_223,
  output [7:0]  io_pipe_phv_out_data_224,
  output [7:0]  io_pipe_phv_out_data_225,
  output [7:0]  io_pipe_phv_out_data_226,
  output [7:0]  io_pipe_phv_out_data_227,
  output [7:0]  io_pipe_phv_out_data_228,
  output [7:0]  io_pipe_phv_out_data_229,
  output [7:0]  io_pipe_phv_out_data_230,
  output [7:0]  io_pipe_phv_out_data_231,
  output [7:0]  io_pipe_phv_out_data_232,
  output [7:0]  io_pipe_phv_out_data_233,
  output [7:0]  io_pipe_phv_out_data_234,
  output [7:0]  io_pipe_phv_out_data_235,
  output [7:0]  io_pipe_phv_out_data_236,
  output [7:0]  io_pipe_phv_out_data_237,
  output [7:0]  io_pipe_phv_out_data_238,
  output [7:0]  io_pipe_phv_out_data_239,
  output [7:0]  io_pipe_phv_out_data_240,
  output [7:0]  io_pipe_phv_out_data_241,
  output [7:0]  io_pipe_phv_out_data_242,
  output [7:0]  io_pipe_phv_out_data_243,
  output [7:0]  io_pipe_phv_out_data_244,
  output [7:0]  io_pipe_phv_out_data_245,
  output [7:0]  io_pipe_phv_out_data_246,
  output [7:0]  io_pipe_phv_out_data_247,
  output [7:0]  io_pipe_phv_out_data_248,
  output [7:0]  io_pipe_phv_out_data_249,
  output [7:0]  io_pipe_phv_out_data_250,
  output [7:0]  io_pipe_phv_out_data_251,
  output [7:0]  io_pipe_phv_out_data_252,
  output [7:0]  io_pipe_phv_out_data_253,
  output [7:0]  io_pipe_phv_out_data_254,
  output [7:0]  io_pipe_phv_out_data_255,
  output [7:0]  io_pipe_phv_out_data_256,
  output [7:0]  io_pipe_phv_out_data_257,
  output [7:0]  io_pipe_phv_out_data_258,
  output [7:0]  io_pipe_phv_out_data_259,
  output [7:0]  io_pipe_phv_out_data_260,
  output [7:0]  io_pipe_phv_out_data_261,
  output [7:0]  io_pipe_phv_out_data_262,
  output [7:0]  io_pipe_phv_out_data_263,
  output [7:0]  io_pipe_phv_out_data_264,
  output [7:0]  io_pipe_phv_out_data_265,
  output [7:0]  io_pipe_phv_out_data_266,
  output [7:0]  io_pipe_phv_out_data_267,
  output [7:0]  io_pipe_phv_out_data_268,
  output [7:0]  io_pipe_phv_out_data_269,
  output [7:0]  io_pipe_phv_out_data_270,
  output [7:0]  io_pipe_phv_out_data_271,
  output [7:0]  io_pipe_phv_out_data_272,
  output [7:0]  io_pipe_phv_out_data_273,
  output [7:0]  io_pipe_phv_out_data_274,
  output [7:0]  io_pipe_phv_out_data_275,
  output [7:0]  io_pipe_phv_out_data_276,
  output [7:0]  io_pipe_phv_out_data_277,
  output [7:0]  io_pipe_phv_out_data_278,
  output [7:0]  io_pipe_phv_out_data_279,
  output [7:0]  io_pipe_phv_out_data_280,
  output [7:0]  io_pipe_phv_out_data_281,
  output [7:0]  io_pipe_phv_out_data_282,
  output [7:0]  io_pipe_phv_out_data_283,
  output [7:0]  io_pipe_phv_out_data_284,
  output [7:0]  io_pipe_phv_out_data_285,
  output [7:0]  io_pipe_phv_out_data_286,
  output [7:0]  io_pipe_phv_out_data_287,
  output [7:0]  io_pipe_phv_out_data_288,
  output [7:0]  io_pipe_phv_out_data_289,
  output [7:0]  io_pipe_phv_out_data_290,
  output [7:0]  io_pipe_phv_out_data_291,
  output [7:0]  io_pipe_phv_out_data_292,
  output [7:0]  io_pipe_phv_out_data_293,
  output [7:0]  io_pipe_phv_out_data_294,
  output [7:0]  io_pipe_phv_out_data_295,
  output [7:0]  io_pipe_phv_out_data_296,
  output [7:0]  io_pipe_phv_out_data_297,
  output [7:0]  io_pipe_phv_out_data_298,
  output [7:0]  io_pipe_phv_out_data_299,
  output [7:0]  io_pipe_phv_out_data_300,
  output [7:0]  io_pipe_phv_out_data_301,
  output [7:0]  io_pipe_phv_out_data_302,
  output [7:0]  io_pipe_phv_out_data_303,
  output [7:0]  io_pipe_phv_out_data_304,
  output [7:0]  io_pipe_phv_out_data_305,
  output [7:0]  io_pipe_phv_out_data_306,
  output [7:0]  io_pipe_phv_out_data_307,
  output [7:0]  io_pipe_phv_out_data_308,
  output [7:0]  io_pipe_phv_out_data_309,
  output [7:0]  io_pipe_phv_out_data_310,
  output [7:0]  io_pipe_phv_out_data_311,
  output [7:0]  io_pipe_phv_out_data_312,
  output [7:0]  io_pipe_phv_out_data_313,
  output [7:0]  io_pipe_phv_out_data_314,
  output [7:0]  io_pipe_phv_out_data_315,
  output [7:0]  io_pipe_phv_out_data_316,
  output [7:0]  io_pipe_phv_out_data_317,
  output [7:0]  io_pipe_phv_out_data_318,
  output [7:0]  io_pipe_phv_out_data_319,
  output [7:0]  io_pipe_phv_out_data_320,
  output [7:0]  io_pipe_phv_out_data_321,
  output [7:0]  io_pipe_phv_out_data_322,
  output [7:0]  io_pipe_phv_out_data_323,
  output [7:0]  io_pipe_phv_out_data_324,
  output [7:0]  io_pipe_phv_out_data_325,
  output [7:0]  io_pipe_phv_out_data_326,
  output [7:0]  io_pipe_phv_out_data_327,
  output [7:0]  io_pipe_phv_out_data_328,
  output [7:0]  io_pipe_phv_out_data_329,
  output [7:0]  io_pipe_phv_out_data_330,
  output [7:0]  io_pipe_phv_out_data_331,
  output [7:0]  io_pipe_phv_out_data_332,
  output [7:0]  io_pipe_phv_out_data_333,
  output [7:0]  io_pipe_phv_out_data_334,
  output [7:0]  io_pipe_phv_out_data_335,
  output [7:0]  io_pipe_phv_out_data_336,
  output [7:0]  io_pipe_phv_out_data_337,
  output [7:0]  io_pipe_phv_out_data_338,
  output [7:0]  io_pipe_phv_out_data_339,
  output [7:0]  io_pipe_phv_out_data_340,
  output [7:0]  io_pipe_phv_out_data_341,
  output [7:0]  io_pipe_phv_out_data_342,
  output [7:0]  io_pipe_phv_out_data_343,
  output [7:0]  io_pipe_phv_out_data_344,
  output [7:0]  io_pipe_phv_out_data_345,
  output [7:0]  io_pipe_phv_out_data_346,
  output [7:0]  io_pipe_phv_out_data_347,
  output [7:0]  io_pipe_phv_out_data_348,
  output [7:0]  io_pipe_phv_out_data_349,
  output [7:0]  io_pipe_phv_out_data_350,
  output [7:0]  io_pipe_phv_out_data_351,
  output [7:0]  io_pipe_phv_out_data_352,
  output [7:0]  io_pipe_phv_out_data_353,
  output [7:0]  io_pipe_phv_out_data_354,
  output [7:0]  io_pipe_phv_out_data_355,
  output [7:0]  io_pipe_phv_out_data_356,
  output [7:0]  io_pipe_phv_out_data_357,
  output [7:0]  io_pipe_phv_out_data_358,
  output [7:0]  io_pipe_phv_out_data_359,
  output [7:0]  io_pipe_phv_out_data_360,
  output [7:0]  io_pipe_phv_out_data_361,
  output [7:0]  io_pipe_phv_out_data_362,
  output [7:0]  io_pipe_phv_out_data_363,
  output [7:0]  io_pipe_phv_out_data_364,
  output [7:0]  io_pipe_phv_out_data_365,
  output [7:0]  io_pipe_phv_out_data_366,
  output [7:0]  io_pipe_phv_out_data_367,
  output [7:0]  io_pipe_phv_out_data_368,
  output [7:0]  io_pipe_phv_out_data_369,
  output [7:0]  io_pipe_phv_out_data_370,
  output [7:0]  io_pipe_phv_out_data_371,
  output [7:0]  io_pipe_phv_out_data_372,
  output [7:0]  io_pipe_phv_out_data_373,
  output [7:0]  io_pipe_phv_out_data_374,
  output [7:0]  io_pipe_phv_out_data_375,
  output [7:0]  io_pipe_phv_out_data_376,
  output [7:0]  io_pipe_phv_out_data_377,
  output [7:0]  io_pipe_phv_out_data_378,
  output [7:0]  io_pipe_phv_out_data_379,
  output [7:0]  io_pipe_phv_out_data_380,
  output [7:0]  io_pipe_phv_out_data_381,
  output [7:0]  io_pipe_phv_out_data_382,
  output [7:0]  io_pipe_phv_out_data_383,
  output [7:0]  io_pipe_phv_out_data_384,
  output [7:0]  io_pipe_phv_out_data_385,
  output [7:0]  io_pipe_phv_out_data_386,
  output [7:0]  io_pipe_phv_out_data_387,
  output [7:0]  io_pipe_phv_out_data_388,
  output [7:0]  io_pipe_phv_out_data_389,
  output [7:0]  io_pipe_phv_out_data_390,
  output [7:0]  io_pipe_phv_out_data_391,
  output [7:0]  io_pipe_phv_out_data_392,
  output [7:0]  io_pipe_phv_out_data_393,
  output [7:0]  io_pipe_phv_out_data_394,
  output [7:0]  io_pipe_phv_out_data_395,
  output [7:0]  io_pipe_phv_out_data_396,
  output [7:0]  io_pipe_phv_out_data_397,
  output [7:0]  io_pipe_phv_out_data_398,
  output [7:0]  io_pipe_phv_out_data_399,
  output [7:0]  io_pipe_phv_out_data_400,
  output [7:0]  io_pipe_phv_out_data_401,
  output [7:0]  io_pipe_phv_out_data_402,
  output [7:0]  io_pipe_phv_out_data_403,
  output [7:0]  io_pipe_phv_out_data_404,
  output [7:0]  io_pipe_phv_out_data_405,
  output [7:0]  io_pipe_phv_out_data_406,
  output [7:0]  io_pipe_phv_out_data_407,
  output [7:0]  io_pipe_phv_out_data_408,
  output [7:0]  io_pipe_phv_out_data_409,
  output [7:0]  io_pipe_phv_out_data_410,
  output [7:0]  io_pipe_phv_out_data_411,
  output [7:0]  io_pipe_phv_out_data_412,
  output [7:0]  io_pipe_phv_out_data_413,
  output [7:0]  io_pipe_phv_out_data_414,
  output [7:0]  io_pipe_phv_out_data_415,
  output [7:0]  io_pipe_phv_out_data_416,
  output [7:0]  io_pipe_phv_out_data_417,
  output [7:0]  io_pipe_phv_out_data_418,
  output [7:0]  io_pipe_phv_out_data_419,
  output [7:0]  io_pipe_phv_out_data_420,
  output [7:0]  io_pipe_phv_out_data_421,
  output [7:0]  io_pipe_phv_out_data_422,
  output [7:0]  io_pipe_phv_out_data_423,
  output [7:0]  io_pipe_phv_out_data_424,
  output [7:0]  io_pipe_phv_out_data_425,
  output [7:0]  io_pipe_phv_out_data_426,
  output [7:0]  io_pipe_phv_out_data_427,
  output [7:0]  io_pipe_phv_out_data_428,
  output [7:0]  io_pipe_phv_out_data_429,
  output [7:0]  io_pipe_phv_out_data_430,
  output [7:0]  io_pipe_phv_out_data_431,
  output [7:0]  io_pipe_phv_out_data_432,
  output [7:0]  io_pipe_phv_out_data_433,
  output [7:0]  io_pipe_phv_out_data_434,
  output [7:0]  io_pipe_phv_out_data_435,
  output [7:0]  io_pipe_phv_out_data_436,
  output [7:0]  io_pipe_phv_out_data_437,
  output [7:0]  io_pipe_phv_out_data_438,
  output [7:0]  io_pipe_phv_out_data_439,
  output [7:0]  io_pipe_phv_out_data_440,
  output [7:0]  io_pipe_phv_out_data_441,
  output [7:0]  io_pipe_phv_out_data_442,
  output [7:0]  io_pipe_phv_out_data_443,
  output [7:0]  io_pipe_phv_out_data_444,
  output [7:0]  io_pipe_phv_out_data_445,
  output [7:0]  io_pipe_phv_out_data_446,
  output [7:0]  io_pipe_phv_out_data_447,
  output [7:0]  io_pipe_phv_out_data_448,
  output [7:0]  io_pipe_phv_out_data_449,
  output [7:0]  io_pipe_phv_out_data_450,
  output [7:0]  io_pipe_phv_out_data_451,
  output [7:0]  io_pipe_phv_out_data_452,
  output [7:0]  io_pipe_phv_out_data_453,
  output [7:0]  io_pipe_phv_out_data_454,
  output [7:0]  io_pipe_phv_out_data_455,
  output [7:0]  io_pipe_phv_out_data_456,
  output [7:0]  io_pipe_phv_out_data_457,
  output [7:0]  io_pipe_phv_out_data_458,
  output [7:0]  io_pipe_phv_out_data_459,
  output [7:0]  io_pipe_phv_out_data_460,
  output [7:0]  io_pipe_phv_out_data_461,
  output [7:0]  io_pipe_phv_out_data_462,
  output [7:0]  io_pipe_phv_out_data_463,
  output [7:0]  io_pipe_phv_out_data_464,
  output [7:0]  io_pipe_phv_out_data_465,
  output [7:0]  io_pipe_phv_out_data_466,
  output [7:0]  io_pipe_phv_out_data_467,
  output [7:0]  io_pipe_phv_out_data_468,
  output [7:0]  io_pipe_phv_out_data_469,
  output [7:0]  io_pipe_phv_out_data_470,
  output [7:0]  io_pipe_phv_out_data_471,
  output [7:0]  io_pipe_phv_out_data_472,
  output [7:0]  io_pipe_phv_out_data_473,
  output [7:0]  io_pipe_phv_out_data_474,
  output [7:0]  io_pipe_phv_out_data_475,
  output [7:0]  io_pipe_phv_out_data_476,
  output [7:0]  io_pipe_phv_out_data_477,
  output [7:0]  io_pipe_phv_out_data_478,
  output [7:0]  io_pipe_phv_out_data_479,
  output [7:0]  io_pipe_phv_out_data_480,
  output [7:0]  io_pipe_phv_out_data_481,
  output [7:0]  io_pipe_phv_out_data_482,
  output [7:0]  io_pipe_phv_out_data_483,
  output [7:0]  io_pipe_phv_out_data_484,
  output [7:0]  io_pipe_phv_out_data_485,
  output [7:0]  io_pipe_phv_out_data_486,
  output [7:0]  io_pipe_phv_out_data_487,
  output [7:0]  io_pipe_phv_out_data_488,
  output [7:0]  io_pipe_phv_out_data_489,
  output [7:0]  io_pipe_phv_out_data_490,
  output [7:0]  io_pipe_phv_out_data_491,
  output [7:0]  io_pipe_phv_out_data_492,
  output [7:0]  io_pipe_phv_out_data_493,
  output [7:0]  io_pipe_phv_out_data_494,
  output [7:0]  io_pipe_phv_out_data_495,
  output [7:0]  io_pipe_phv_out_data_496,
  output [7:0]  io_pipe_phv_out_data_497,
  output [7:0]  io_pipe_phv_out_data_498,
  output [7:0]  io_pipe_phv_out_data_499,
  output [7:0]  io_pipe_phv_out_data_500,
  output [7:0]  io_pipe_phv_out_data_501,
  output [7:0]  io_pipe_phv_out_data_502,
  output [7:0]  io_pipe_phv_out_data_503,
  output [7:0]  io_pipe_phv_out_data_504,
  output [7:0]  io_pipe_phv_out_data_505,
  output [7:0]  io_pipe_phv_out_data_506,
  output [7:0]  io_pipe_phv_out_data_507,
  output [7:0]  io_pipe_phv_out_data_508,
  output [7:0]  io_pipe_phv_out_data_509,
  output [7:0]  io_pipe_phv_out_data_510,
  output [7:0]  io_pipe_phv_out_data_511,
  output [3:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  input  [7:0]  io_args_in_0,
  input  [7:0]  io_args_in_1,
  input  [7:0]  io_args_in_2,
  input  [7:0]  io_args_in_3,
  input  [7:0]  io_args_in_4,
  input  [7:0]  io_args_in_5,
  input  [7:0]  io_args_in_6,
  input  [17:0] io_vliw_in_0,
  input  [17:0] io_vliw_in_1,
  input  [17:0] io_vliw_in_2,
  input  [17:0] io_vliw_in_3,
  input  [17:0] io_vliw_in_4,
  input  [17:0] io_vliw_in_5,
  input  [17:0] io_vliw_in_6,
  input  [17:0] io_vliw_in_7,
  input  [17:0] io_vliw_in_8,
  input  [17:0] io_vliw_in_9,
  input  [17:0] io_vliw_in_10,
  input  [17:0] io_vliw_in_11,
  input  [17:0] io_vliw_in_12,
  input  [17:0] io_vliw_in_13,
  input  [17:0] io_vliw_in_14,
  input  [17:0] io_vliw_in_15,
  input  [17:0] io_vliw_in_16,
  input  [17:0] io_vliw_in_17,
  input  [17:0] io_vliw_in_18,
  input  [17:0] io_vliw_in_19,
  input  [17:0] io_vliw_in_20,
  input  [17:0] io_vliw_in_21,
  input  [17:0] io_vliw_in_22,
  input  [17:0] io_vliw_in_23,
  input  [17:0] io_vliw_in_24,
  input  [17:0] io_vliw_in_25,
  input  [17:0] io_vliw_in_26,
  input  [17:0] io_vliw_in_27,
  input  [17:0] io_vliw_in_28,
  input  [17:0] io_vliw_in_29,
  input  [17:0] io_vliw_in_30,
  input  [17:0] io_vliw_in_31,
  input  [17:0] io_vliw_in_32,
  input  [17:0] io_vliw_in_33,
  input  [17:0] io_vliw_in_34,
  input  [17:0] io_vliw_in_35,
  input  [17:0] io_vliw_in_36,
  input  [17:0] io_vliw_in_37,
  input  [17:0] io_vliw_in_38,
  input  [17:0] io_vliw_in_39,
  input  [17:0] io_vliw_in_40,
  input  [17:0] io_vliw_in_41,
  input  [17:0] io_vliw_in_42,
  input  [17:0] io_vliw_in_43,
  input  [17:0] io_vliw_in_44,
  input  [17:0] io_vliw_in_45,
  input  [17:0] io_vliw_in_46,
  input  [17:0] io_vliw_in_47,
  input  [17:0] io_vliw_in_48,
  input  [17:0] io_vliw_in_49,
  input  [17:0] io_vliw_in_50,
  input  [17:0] io_vliw_in_51,
  input  [17:0] io_vliw_in_52,
  input  [17:0] io_vliw_in_53,
  input  [17:0] io_vliw_in_54,
  input  [17:0] io_vliw_in_55,
  input  [17:0] io_vliw_in_56,
  input  [17:0] io_vliw_in_57,
  input  [17:0] io_vliw_in_58,
  input  [17:0] io_vliw_in_59,
  input  [17:0] io_vliw_in_60,
  input  [17:0] io_vliw_in_61,
  input  [17:0] io_vliw_in_62,
  input  [17:0] io_vliw_in_63,
  input  [17:0] io_vliw_in_64,
  input  [17:0] io_vliw_in_65,
  input  [17:0] io_vliw_in_66,
  input  [17:0] io_vliw_in_67,
  input  [17:0] io_vliw_in_68,
  input  [17:0] io_vliw_in_69,
  input  [14:0] io_nid_in,
  output [14:0] io_nid_out,
  output [1:0]  io_tag_out_0,
  output [1:0]  io_tag_out_1,
  output [1:0]  io_tag_out_2,
  output [1:0]  io_tag_out_3,
  output [1:0]  io_tag_out_4,
  output [1:0]  io_tag_out_5,
  output [1:0]  io_tag_out_6,
  output [1:0]  io_tag_out_7,
  output [1:0]  io_tag_out_8,
  output [1:0]  io_tag_out_9,
  output [1:0]  io_tag_out_10,
  output [1:0]  io_tag_out_11,
  output [1:0]  io_tag_out_12,
  output [1:0]  io_tag_out_13,
  output [1:0]  io_tag_out_14,
  output [1:0]  io_tag_out_15,
  output [1:0]  io_tag_out_16,
  output [1:0]  io_tag_out_17,
  output [1:0]  io_tag_out_18,
  output [1:0]  io_tag_out_19,
  output [1:0]  io_tag_out_20,
  output [1:0]  io_tag_out_21,
  output [1:0]  io_tag_out_22,
  output [1:0]  io_tag_out_23,
  output [1:0]  io_tag_out_24,
  output [1:0]  io_tag_out_25,
  output [1:0]  io_tag_out_26,
  output [1:0]  io_tag_out_27,
  output [1:0]  io_tag_out_28,
  output [1:0]  io_tag_out_29,
  output [1:0]  io_tag_out_30,
  output [1:0]  io_tag_out_31,
  output [1:0]  io_tag_out_32,
  output [1:0]  io_tag_out_33,
  output [1:0]  io_tag_out_34,
  output [1:0]  io_tag_out_35,
  output [1:0]  io_tag_out_36,
  output [1:0]  io_tag_out_37,
  output [1:0]  io_tag_out_38,
  output [1:0]  io_tag_out_39,
  output [1:0]  io_tag_out_40,
  output [1:0]  io_tag_out_41,
  output [1:0]  io_tag_out_42,
  output [1:0]  io_tag_out_43,
  output [1:0]  io_tag_out_44,
  output [1:0]  io_tag_out_45,
  output [1:0]  io_tag_out_46,
  output [1:0]  io_tag_out_47,
  output [1:0]  io_tag_out_48,
  output [1:0]  io_tag_out_49,
  output [1:0]  io_tag_out_50,
  output [1:0]  io_tag_out_51,
  output [1:0]  io_tag_out_52,
  output [1:0]  io_tag_out_53,
  output [1:0]  io_tag_out_54,
  output [1:0]  io_tag_out_55,
  output [1:0]  io_tag_out_56,
  output [1:0]  io_tag_out_57,
  output [1:0]  io_tag_out_58,
  output [1:0]  io_tag_out_59,
  output [1:0]  io_tag_out_60,
  output [1:0]  io_tag_out_61,
  output [1:0]  io_tag_out_62,
  output [1:0]  io_tag_out_63,
  output [1:0]  io_tag_out_64,
  output [1:0]  io_tag_out_65,
  output [1:0]  io_tag_out_66,
  output [1:0]  io_tag_out_67,
  output [1:0]  io_tag_out_68,
  output [1:0]  io_tag_out_69,
  output [7:0]  io_field_set_field8_0,
  output [7:0]  io_field_set_field8_1,
  output [7:0]  io_field_set_field8_2,
  output [7:0]  io_field_set_field8_3,
  output [7:0]  io_field_set_field8_4,
  output [7:0]  io_field_set_field8_5,
  output [7:0]  io_field_set_field8_6,
  output [7:0]  io_field_set_field8_7,
  output [7:0]  io_field_set_field8_8,
  output [7:0]  io_field_set_field8_9,
  output [7:0]  io_field_set_field8_10,
  output [7:0]  io_field_set_field8_11,
  output [7:0]  io_field_set_field8_12,
  output [7:0]  io_field_set_field8_13,
  output [7:0]  io_field_set_field8_14,
  output [7:0]  io_field_set_field8_15,
  output [7:0]  io_field_set_field8_16,
  output [7:0]  io_field_set_field8_17,
  output [7:0]  io_field_set_field8_18,
  output [7:0]  io_field_set_field8_19,
  output [7:0]  io_field_set_field8_20,
  output [7:0]  io_field_set_field8_21,
  output [7:0]  io_field_set_field8_22,
  output [7:0]  io_field_set_field8_23,
  output [7:0]  io_field_set_field8_24,
  output [7:0]  io_field_set_field8_25,
  output [7:0]  io_field_set_field8_26,
  output [7:0]  io_field_set_field8_27,
  output [7:0]  io_field_set_field8_28,
  output [7:0]  io_field_set_field8_29,
  output [7:0]  io_field_set_field8_30,
  output [7:0]  io_field_set_field8_31,
  output [7:0]  io_field_set_field8_32,
  output [7:0]  io_field_set_field8_33,
  output [7:0]  io_field_set_field8_34,
  output [7:0]  io_field_set_field8_35,
  output [7:0]  io_field_set_field8_36,
  output [7:0]  io_field_set_field8_37,
  output [7:0]  io_field_set_field8_38,
  output [7:0]  io_field_set_field8_39,
  output [7:0]  io_field_set_field8_40,
  output [7:0]  io_field_set_field8_41,
  output [7:0]  io_field_set_field8_42,
  output [7:0]  io_field_set_field8_43,
  output [7:0]  io_field_set_field8_44,
  output [7:0]  io_field_set_field8_45,
  output [7:0]  io_field_set_field8_46,
  output [7:0]  io_field_set_field8_47,
  output [7:0]  io_field_set_field8_48,
  output [7:0]  io_field_set_field8_49,
  output [7:0]  io_field_set_field8_50,
  output [7:0]  io_field_set_field8_51,
  output [7:0]  io_field_set_field8_52,
  output [7:0]  io_field_set_field8_53,
  output [7:0]  io_field_set_field8_54,
  output [7:0]  io_field_set_field8_55,
  output [7:0]  io_field_set_field8_56,
  output [7:0]  io_field_set_field8_57,
  output [7:0]  io_field_set_field8_58,
  output [7:0]  io_field_set_field8_59,
  output [7:0]  io_field_set_field8_60,
  output [7:0]  io_field_set_field8_61,
  output [7:0]  io_field_set_field8_62,
  output [7:0]  io_field_set_field8_63,
  output [15:0] io_field_set_field16_0,
  output [15:0] io_field_set_field16_1,
  output [15:0] io_field_set_field16_2,
  output [15:0] io_field_set_field16_3,
  output [15:0] io_field_set_field16_4,
  output [15:0] io_field_set_field16_5
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_1; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_2; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_3; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_4; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_5; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_6; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_7; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_8; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_9; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_10; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_11; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_12; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_13; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_14; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_15; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_16; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_17; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_18; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_19; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_20; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_21; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_22; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_23; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_24; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_25; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_26; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_27; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_28; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_29; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_30; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_31; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_32; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_33; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_34; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_35; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_36; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_37; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_38; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_39; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_40; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_41; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_42; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_43; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_44; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_45; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_46; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_47; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_48; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_49; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_50; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_51; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_52; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_53; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_54; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_55; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_56; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_57; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_58; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_59; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_60; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_61; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_62; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_63; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_64; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_65; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_66; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_67; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_68; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_69; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_70; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_71; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_72; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_73; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_74; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_75; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_76; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_77; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_78; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_79; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_80; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_81; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_82; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_83; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_84; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_85; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_86; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_87; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_88; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_89; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_90; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_91; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_92; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_93; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_94; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_95; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_96; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_97; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_98; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_99; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_100; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_101; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_102; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_103; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_104; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_105; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_106; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_107; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_108; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_109; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_110; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_111; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_112; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_113; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_114; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_115; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_116; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_117; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_118; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_119; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_120; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_121; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_122; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_123; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_124; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_125; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_126; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_127; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_128; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_129; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_130; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_131; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_132; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_133; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_134; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_135; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_136; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_137; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_138; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_139; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_140; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_141; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_142; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_143; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_144; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_145; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_146; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_147; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_148; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_149; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_150; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_151; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_152; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_153; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_154; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_155; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_156; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_157; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_158; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_159; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_160; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_161; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_162; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_163; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_164; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_165; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_166; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_167; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_168; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_169; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_170; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_171; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_172; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_173; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_174; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_175; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_176; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_177; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_178; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_179; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_180; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_181; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_182; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_183; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_184; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_185; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_186; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_187; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_188; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_189; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_190; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_191; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_192; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_193; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_194; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_195; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_196; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_197; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_198; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_199; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_200; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_201; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_202; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_203; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_204; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_205; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_206; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_207; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_208; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_209; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_210; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_211; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_212; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_213; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_214; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_215; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_216; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_217; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_218; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_219; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_220; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_221; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_222; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_223; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_224; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_225; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_226; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_227; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_228; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_229; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_230; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_231; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_232; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_233; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_234; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_235; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_236; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_237; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_238; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_239; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_240; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_241; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_242; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_243; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_244; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_245; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_246; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_247; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_248; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_249; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_250; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_251; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_252; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_253; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_254; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_255; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_256; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_257; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_258; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_259; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_260; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_261; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_262; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_263; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_264; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_265; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_266; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_267; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_268; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_269; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_270; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_271; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_272; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_273; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_274; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_275; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_276; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_277; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_278; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_279; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_280; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_281; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_282; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_283; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_284; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_285; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_286; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_287; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_288; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_289; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_290; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_291; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_292; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_293; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_294; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_295; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_296; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_297; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_298; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_299; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_300; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_301; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_302; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_303; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_304; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_305; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_306; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_307; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_308; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_309; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_310; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_311; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_312; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_313; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_314; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_315; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_316; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_317; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_318; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_319; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_320; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_321; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_322; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_323; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_324; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_325; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_326; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_327; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_328; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_329; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_330; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_331; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_332; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_333; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_334; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_335; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_336; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_337; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_338; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_339; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_340; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_341; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_342; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_343; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_344; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_345; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_346; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_347; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_348; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_349; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_350; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_351; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_352; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_353; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_354; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_355; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_356; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_357; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_358; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_359; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_360; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_361; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_362; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_363; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_364; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_365; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_366; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_367; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_368; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_369; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_370; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_371; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_372; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_373; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_374; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_375; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_376; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_377; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_378; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_379; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_380; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_381; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_382; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_383; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_384; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_385; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_386; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_387; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_388; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_389; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_390; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_391; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_392; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_393; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_394; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_395; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_396; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_397; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_398; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_399; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_400; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_401; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_402; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_403; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_404; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_405; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_406; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_407; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_408; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_409; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_410; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_411; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_412; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_413; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_414; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_415; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_416; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_417; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_418; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_419; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_420; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_421; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_422; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_423; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_424; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_425; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_426; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_427; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_428; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_429; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_430; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_431; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_432; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_433; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_434; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_435; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_436; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_437; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_438; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_439; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_440; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_441; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_442; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_443; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_444; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_445; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_446; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_447; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_448; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_449; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_450; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_451; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_452; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_453; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_454; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_455; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_456; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_457; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_458; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_459; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_460; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_461; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_462; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_463; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_464; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_465; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_466; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_467; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_468; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_469; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_470; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_471; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_472; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_473; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_474; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_475; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_476; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_477; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_478; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_479; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_480; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_481; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_482; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_483; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_484; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_485; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_486; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_487; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_488; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_489; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_490; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_491; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_492; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_493; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_494; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_495; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_496; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_497; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_498; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_499; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_500; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_501; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_502; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_503; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_504; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_505; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_506; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_507; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_508; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_509; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_510; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_511; // @[executor_pisa.scala 161:22]
  reg [3:0] phv_next_processor_id; // @[executor_pisa.scala 161:22]
  reg  phv_next_config_id; // @[executor_pisa.scala 161:22]
  reg [7:0] args_0; // @[executor_pisa.scala 165:23]
  reg [7:0] args_1; // @[executor_pisa.scala 165:23]
  reg [7:0] args_2; // @[executor_pisa.scala 165:23]
  reg [7:0] args_3; // @[executor_pisa.scala 165:23]
  reg [7:0] args_4; // @[executor_pisa.scala 165:23]
  reg [7:0] args_5; // @[executor_pisa.scala 165:23]
  reg [7:0] args_6; // @[executor_pisa.scala 165:23]
  reg [17:0] vliw_0; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_1; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_2; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_3; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_4; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_5; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_6; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_7; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_8; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_9; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_10; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_11; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_12; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_13; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_14; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_15; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_16; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_17; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_18; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_19; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_20; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_21; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_22; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_23; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_24; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_25; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_26; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_27; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_28; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_29; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_30; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_31; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_32; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_33; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_34; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_35; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_36; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_37; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_38; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_39; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_40; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_41; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_42; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_43; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_44; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_45; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_46; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_47; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_48; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_49; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_50; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_51; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_52; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_53; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_54; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_55; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_56; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_57; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_58; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_59; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_60; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_61; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_62; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_63; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_64; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_65; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_66; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_67; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_68; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_69; // @[executor_pisa.scala 168:23]
  reg [14:0] nid; // @[executor_pisa.scala 171:23]
  wire [3:0] opcode = vliw_0[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2 = vliw_0[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset = parameter_2[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length = parameter_2[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T = {{1'd0}, args_offset}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset = _total_offset_T[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1 = 3'h1 == total_offset ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2 = 3'h2 == total_offset ? args_2 : _GEN_1; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3 = 3'h3 == total_offset ? args_3 : _GEN_2; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4 = 3'h4 == total_offset ? args_4 : _GEN_3; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5 = 3'h5 == total_offset ? args_5 : _GEN_4; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_6 = 3'h6 == total_offset ? args_6 : _GEN_5; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_7 = total_offset < 3'h7 ? _GEN_6 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_0 = 3'h0 < args_length ? _GEN_7 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_9 = opcode == 4'ha ? field_bytes_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_10 = opcode == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_3 = opcode == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_1 = _T_3 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_11 = opcode == 4'h8 | opcode == 4'hb ? parameter_2[7:0] : _GEN_9; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_12 = opcode == 4'h8 | opcode == 4'hb ? _field_tag_T_1 : _GEN_10; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_13 = 14'h0 == parameter_2 ? phv_data_0 : _GEN_11; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_14 = 14'h1 == parameter_2 ? phv_data_1 : _GEN_13; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_15 = 14'h2 == parameter_2 ? phv_data_2 : _GEN_14; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_16 = 14'h3 == parameter_2 ? phv_data_3 : _GEN_15; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_17 = 14'h4 == parameter_2 ? phv_data_4 : _GEN_16; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_18 = 14'h5 == parameter_2 ? phv_data_5 : _GEN_17; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_19 = 14'h6 == parameter_2 ? phv_data_6 : _GEN_18; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_20 = 14'h7 == parameter_2 ? phv_data_7 : _GEN_19; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_21 = 14'h8 == parameter_2 ? phv_data_8 : _GEN_20; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_22 = 14'h9 == parameter_2 ? phv_data_9 : _GEN_21; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_23 = 14'ha == parameter_2 ? phv_data_10 : _GEN_22; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_24 = 14'hb == parameter_2 ? phv_data_11 : _GEN_23; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_25 = 14'hc == parameter_2 ? phv_data_12 : _GEN_24; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_26 = 14'hd == parameter_2 ? phv_data_13 : _GEN_25; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_27 = 14'he == parameter_2 ? phv_data_14 : _GEN_26; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_28 = 14'hf == parameter_2 ? phv_data_15 : _GEN_27; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_29 = 14'h10 == parameter_2 ? phv_data_16 : _GEN_28; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_30 = 14'h11 == parameter_2 ? phv_data_17 : _GEN_29; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_31 = 14'h12 == parameter_2 ? phv_data_18 : _GEN_30; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_32 = 14'h13 == parameter_2 ? phv_data_19 : _GEN_31; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_33 = 14'h14 == parameter_2 ? phv_data_20 : _GEN_32; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_34 = 14'h15 == parameter_2 ? phv_data_21 : _GEN_33; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_35 = 14'h16 == parameter_2 ? phv_data_22 : _GEN_34; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_36 = 14'h17 == parameter_2 ? phv_data_23 : _GEN_35; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_37 = 14'h18 == parameter_2 ? phv_data_24 : _GEN_36; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_38 = 14'h19 == parameter_2 ? phv_data_25 : _GEN_37; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_39 = 14'h1a == parameter_2 ? phv_data_26 : _GEN_38; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_40 = 14'h1b == parameter_2 ? phv_data_27 : _GEN_39; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_41 = 14'h1c == parameter_2 ? phv_data_28 : _GEN_40; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_42 = 14'h1d == parameter_2 ? phv_data_29 : _GEN_41; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_43 = 14'h1e == parameter_2 ? phv_data_30 : _GEN_42; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_44 = 14'h1f == parameter_2 ? phv_data_31 : _GEN_43; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_45 = 14'h20 == parameter_2 ? phv_data_32 : _GEN_44; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_46 = 14'h21 == parameter_2 ? phv_data_33 : _GEN_45; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_47 = 14'h22 == parameter_2 ? phv_data_34 : _GEN_46; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_48 = 14'h23 == parameter_2 ? phv_data_35 : _GEN_47; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_49 = 14'h24 == parameter_2 ? phv_data_36 : _GEN_48; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_50 = 14'h25 == parameter_2 ? phv_data_37 : _GEN_49; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_51 = 14'h26 == parameter_2 ? phv_data_38 : _GEN_50; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_52 = 14'h27 == parameter_2 ? phv_data_39 : _GEN_51; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_53 = 14'h28 == parameter_2 ? phv_data_40 : _GEN_52; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_54 = 14'h29 == parameter_2 ? phv_data_41 : _GEN_53; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_55 = 14'h2a == parameter_2 ? phv_data_42 : _GEN_54; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_56 = 14'h2b == parameter_2 ? phv_data_43 : _GEN_55; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_57 = 14'h2c == parameter_2 ? phv_data_44 : _GEN_56; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_58 = 14'h2d == parameter_2 ? phv_data_45 : _GEN_57; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_59 = 14'h2e == parameter_2 ? phv_data_46 : _GEN_58; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_60 = 14'h2f == parameter_2 ? phv_data_47 : _GEN_59; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_61 = 14'h30 == parameter_2 ? phv_data_48 : _GEN_60; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_62 = 14'h31 == parameter_2 ? phv_data_49 : _GEN_61; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_63 = 14'h32 == parameter_2 ? phv_data_50 : _GEN_62; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_64 = 14'h33 == parameter_2 ? phv_data_51 : _GEN_63; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_65 = 14'h34 == parameter_2 ? phv_data_52 : _GEN_64; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_66 = 14'h35 == parameter_2 ? phv_data_53 : _GEN_65; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_67 = 14'h36 == parameter_2 ? phv_data_54 : _GEN_66; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_68 = 14'h37 == parameter_2 ? phv_data_55 : _GEN_67; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_69 = 14'h38 == parameter_2 ? phv_data_56 : _GEN_68; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_70 = 14'h39 == parameter_2 ? phv_data_57 : _GEN_69; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_71 = 14'h3a == parameter_2 ? phv_data_58 : _GEN_70; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_72 = 14'h3b == parameter_2 ? phv_data_59 : _GEN_71; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_73 = 14'h3c == parameter_2 ? phv_data_60 : _GEN_72; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_74 = 14'h3d == parameter_2 ? phv_data_61 : _GEN_73; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_75 = 14'h3e == parameter_2 ? phv_data_62 : _GEN_74; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_76 = 14'h3f == parameter_2 ? phv_data_63 : _GEN_75; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_1 = vliw_1[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_1 = vliw_1[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_1 = parameter_2_1[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_1 = parameter_2_1[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_1 = {{1'd0}, args_offset_1}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_1 = _total_offset_T_1[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_80 = 3'h1 == total_offset_1 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_81 = 3'h2 == total_offset_1 ? args_2 : _GEN_80; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_82 = 3'h3 == total_offset_1 ? args_3 : _GEN_81; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_83 = 3'h4 == total_offset_1 ? args_4 : _GEN_82; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_84 = 3'h5 == total_offset_1 ? args_5 : _GEN_83; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_85 = 3'h6 == total_offset_1 ? args_6 : _GEN_84; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_86 = total_offset_1 < 3'h7 ? _GEN_85 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_1_0 = 3'h0 < args_length_1 ? _GEN_86 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_88 = opcode_1 == 4'ha ? field_bytes_1_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_89 = opcode_1 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_74 = opcode_1 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_3 = _T_74 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_90 = opcode_1 == 4'h8 | opcode_1 == 4'hb ? parameter_2_1[7:0] : _GEN_88; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_91 = opcode_1 == 4'h8 | opcode_1 == 4'hb ? _field_tag_T_3 : _GEN_89; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_92 = 14'h0 == parameter_2_1 ? phv_data_0 : _GEN_90; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_93 = 14'h1 == parameter_2_1 ? phv_data_1 : _GEN_92; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_94 = 14'h2 == parameter_2_1 ? phv_data_2 : _GEN_93; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_95 = 14'h3 == parameter_2_1 ? phv_data_3 : _GEN_94; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_96 = 14'h4 == parameter_2_1 ? phv_data_4 : _GEN_95; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_97 = 14'h5 == parameter_2_1 ? phv_data_5 : _GEN_96; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_98 = 14'h6 == parameter_2_1 ? phv_data_6 : _GEN_97; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_99 = 14'h7 == parameter_2_1 ? phv_data_7 : _GEN_98; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_100 = 14'h8 == parameter_2_1 ? phv_data_8 : _GEN_99; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_101 = 14'h9 == parameter_2_1 ? phv_data_9 : _GEN_100; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_102 = 14'ha == parameter_2_1 ? phv_data_10 : _GEN_101; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_103 = 14'hb == parameter_2_1 ? phv_data_11 : _GEN_102; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_104 = 14'hc == parameter_2_1 ? phv_data_12 : _GEN_103; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_105 = 14'hd == parameter_2_1 ? phv_data_13 : _GEN_104; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_106 = 14'he == parameter_2_1 ? phv_data_14 : _GEN_105; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_107 = 14'hf == parameter_2_1 ? phv_data_15 : _GEN_106; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_108 = 14'h10 == parameter_2_1 ? phv_data_16 : _GEN_107; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_109 = 14'h11 == parameter_2_1 ? phv_data_17 : _GEN_108; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_110 = 14'h12 == parameter_2_1 ? phv_data_18 : _GEN_109; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_111 = 14'h13 == parameter_2_1 ? phv_data_19 : _GEN_110; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_112 = 14'h14 == parameter_2_1 ? phv_data_20 : _GEN_111; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_113 = 14'h15 == parameter_2_1 ? phv_data_21 : _GEN_112; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_114 = 14'h16 == parameter_2_1 ? phv_data_22 : _GEN_113; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_115 = 14'h17 == parameter_2_1 ? phv_data_23 : _GEN_114; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_116 = 14'h18 == parameter_2_1 ? phv_data_24 : _GEN_115; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_117 = 14'h19 == parameter_2_1 ? phv_data_25 : _GEN_116; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_118 = 14'h1a == parameter_2_1 ? phv_data_26 : _GEN_117; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_119 = 14'h1b == parameter_2_1 ? phv_data_27 : _GEN_118; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_120 = 14'h1c == parameter_2_1 ? phv_data_28 : _GEN_119; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_121 = 14'h1d == parameter_2_1 ? phv_data_29 : _GEN_120; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_122 = 14'h1e == parameter_2_1 ? phv_data_30 : _GEN_121; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_123 = 14'h1f == parameter_2_1 ? phv_data_31 : _GEN_122; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_124 = 14'h20 == parameter_2_1 ? phv_data_32 : _GEN_123; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_125 = 14'h21 == parameter_2_1 ? phv_data_33 : _GEN_124; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_126 = 14'h22 == parameter_2_1 ? phv_data_34 : _GEN_125; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_127 = 14'h23 == parameter_2_1 ? phv_data_35 : _GEN_126; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_128 = 14'h24 == parameter_2_1 ? phv_data_36 : _GEN_127; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_129 = 14'h25 == parameter_2_1 ? phv_data_37 : _GEN_128; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_130 = 14'h26 == parameter_2_1 ? phv_data_38 : _GEN_129; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_131 = 14'h27 == parameter_2_1 ? phv_data_39 : _GEN_130; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_132 = 14'h28 == parameter_2_1 ? phv_data_40 : _GEN_131; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_133 = 14'h29 == parameter_2_1 ? phv_data_41 : _GEN_132; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_134 = 14'h2a == parameter_2_1 ? phv_data_42 : _GEN_133; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_135 = 14'h2b == parameter_2_1 ? phv_data_43 : _GEN_134; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_136 = 14'h2c == parameter_2_1 ? phv_data_44 : _GEN_135; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_137 = 14'h2d == parameter_2_1 ? phv_data_45 : _GEN_136; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_138 = 14'h2e == parameter_2_1 ? phv_data_46 : _GEN_137; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_139 = 14'h2f == parameter_2_1 ? phv_data_47 : _GEN_138; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_140 = 14'h30 == parameter_2_1 ? phv_data_48 : _GEN_139; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_141 = 14'h31 == parameter_2_1 ? phv_data_49 : _GEN_140; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_142 = 14'h32 == parameter_2_1 ? phv_data_50 : _GEN_141; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_143 = 14'h33 == parameter_2_1 ? phv_data_51 : _GEN_142; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_144 = 14'h34 == parameter_2_1 ? phv_data_52 : _GEN_143; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_145 = 14'h35 == parameter_2_1 ? phv_data_53 : _GEN_144; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_146 = 14'h36 == parameter_2_1 ? phv_data_54 : _GEN_145; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_147 = 14'h37 == parameter_2_1 ? phv_data_55 : _GEN_146; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_148 = 14'h38 == parameter_2_1 ? phv_data_56 : _GEN_147; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_149 = 14'h39 == parameter_2_1 ? phv_data_57 : _GEN_148; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_150 = 14'h3a == parameter_2_1 ? phv_data_58 : _GEN_149; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_151 = 14'h3b == parameter_2_1 ? phv_data_59 : _GEN_150; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_152 = 14'h3c == parameter_2_1 ? phv_data_60 : _GEN_151; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_153 = 14'h3d == parameter_2_1 ? phv_data_61 : _GEN_152; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_154 = 14'h3e == parameter_2_1 ? phv_data_62 : _GEN_153; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_155 = 14'h3f == parameter_2_1 ? phv_data_63 : _GEN_154; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_2 = vliw_2[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_2 = vliw_2[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_2 = parameter_2_2[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_2 = parameter_2_2[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_2 = {{1'd0}, args_offset_2}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_2 = _total_offset_T_2[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_159 = 3'h1 == total_offset_2 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_160 = 3'h2 == total_offset_2 ? args_2 : _GEN_159; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_161 = 3'h3 == total_offset_2 ? args_3 : _GEN_160; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_162 = 3'h4 == total_offset_2 ? args_4 : _GEN_161; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_163 = 3'h5 == total_offset_2 ? args_5 : _GEN_162; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_164 = 3'h6 == total_offset_2 ? args_6 : _GEN_163; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_165 = total_offset_2 < 3'h7 ? _GEN_164 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_2_0 = 3'h0 < args_length_2 ? _GEN_165 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_167 = opcode_2 == 4'ha ? field_bytes_2_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_168 = opcode_2 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_145 = opcode_2 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_5 = _T_145 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_169 = opcode_2 == 4'h8 | opcode_2 == 4'hb ? parameter_2_2[7:0] : _GEN_167; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_170 = opcode_2 == 4'h8 | opcode_2 == 4'hb ? _field_tag_T_5 : _GEN_168; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_171 = 14'h0 == parameter_2_2 ? phv_data_0 : _GEN_169; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_172 = 14'h1 == parameter_2_2 ? phv_data_1 : _GEN_171; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_173 = 14'h2 == parameter_2_2 ? phv_data_2 : _GEN_172; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_174 = 14'h3 == parameter_2_2 ? phv_data_3 : _GEN_173; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_175 = 14'h4 == parameter_2_2 ? phv_data_4 : _GEN_174; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_176 = 14'h5 == parameter_2_2 ? phv_data_5 : _GEN_175; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_177 = 14'h6 == parameter_2_2 ? phv_data_6 : _GEN_176; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_178 = 14'h7 == parameter_2_2 ? phv_data_7 : _GEN_177; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_179 = 14'h8 == parameter_2_2 ? phv_data_8 : _GEN_178; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_180 = 14'h9 == parameter_2_2 ? phv_data_9 : _GEN_179; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_181 = 14'ha == parameter_2_2 ? phv_data_10 : _GEN_180; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_182 = 14'hb == parameter_2_2 ? phv_data_11 : _GEN_181; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_183 = 14'hc == parameter_2_2 ? phv_data_12 : _GEN_182; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_184 = 14'hd == parameter_2_2 ? phv_data_13 : _GEN_183; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_185 = 14'he == parameter_2_2 ? phv_data_14 : _GEN_184; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_186 = 14'hf == parameter_2_2 ? phv_data_15 : _GEN_185; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_187 = 14'h10 == parameter_2_2 ? phv_data_16 : _GEN_186; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_188 = 14'h11 == parameter_2_2 ? phv_data_17 : _GEN_187; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_189 = 14'h12 == parameter_2_2 ? phv_data_18 : _GEN_188; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_190 = 14'h13 == parameter_2_2 ? phv_data_19 : _GEN_189; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_191 = 14'h14 == parameter_2_2 ? phv_data_20 : _GEN_190; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_192 = 14'h15 == parameter_2_2 ? phv_data_21 : _GEN_191; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_193 = 14'h16 == parameter_2_2 ? phv_data_22 : _GEN_192; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_194 = 14'h17 == parameter_2_2 ? phv_data_23 : _GEN_193; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_195 = 14'h18 == parameter_2_2 ? phv_data_24 : _GEN_194; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_196 = 14'h19 == parameter_2_2 ? phv_data_25 : _GEN_195; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_197 = 14'h1a == parameter_2_2 ? phv_data_26 : _GEN_196; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_198 = 14'h1b == parameter_2_2 ? phv_data_27 : _GEN_197; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_199 = 14'h1c == parameter_2_2 ? phv_data_28 : _GEN_198; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_200 = 14'h1d == parameter_2_2 ? phv_data_29 : _GEN_199; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_201 = 14'h1e == parameter_2_2 ? phv_data_30 : _GEN_200; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_202 = 14'h1f == parameter_2_2 ? phv_data_31 : _GEN_201; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_203 = 14'h20 == parameter_2_2 ? phv_data_32 : _GEN_202; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_204 = 14'h21 == parameter_2_2 ? phv_data_33 : _GEN_203; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_205 = 14'h22 == parameter_2_2 ? phv_data_34 : _GEN_204; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_206 = 14'h23 == parameter_2_2 ? phv_data_35 : _GEN_205; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_207 = 14'h24 == parameter_2_2 ? phv_data_36 : _GEN_206; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_208 = 14'h25 == parameter_2_2 ? phv_data_37 : _GEN_207; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_209 = 14'h26 == parameter_2_2 ? phv_data_38 : _GEN_208; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_210 = 14'h27 == parameter_2_2 ? phv_data_39 : _GEN_209; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_211 = 14'h28 == parameter_2_2 ? phv_data_40 : _GEN_210; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_212 = 14'h29 == parameter_2_2 ? phv_data_41 : _GEN_211; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_213 = 14'h2a == parameter_2_2 ? phv_data_42 : _GEN_212; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_214 = 14'h2b == parameter_2_2 ? phv_data_43 : _GEN_213; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_215 = 14'h2c == parameter_2_2 ? phv_data_44 : _GEN_214; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_216 = 14'h2d == parameter_2_2 ? phv_data_45 : _GEN_215; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_217 = 14'h2e == parameter_2_2 ? phv_data_46 : _GEN_216; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_218 = 14'h2f == parameter_2_2 ? phv_data_47 : _GEN_217; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_219 = 14'h30 == parameter_2_2 ? phv_data_48 : _GEN_218; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_220 = 14'h31 == parameter_2_2 ? phv_data_49 : _GEN_219; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_221 = 14'h32 == parameter_2_2 ? phv_data_50 : _GEN_220; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_222 = 14'h33 == parameter_2_2 ? phv_data_51 : _GEN_221; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_223 = 14'h34 == parameter_2_2 ? phv_data_52 : _GEN_222; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_224 = 14'h35 == parameter_2_2 ? phv_data_53 : _GEN_223; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_225 = 14'h36 == parameter_2_2 ? phv_data_54 : _GEN_224; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_226 = 14'h37 == parameter_2_2 ? phv_data_55 : _GEN_225; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_227 = 14'h38 == parameter_2_2 ? phv_data_56 : _GEN_226; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_228 = 14'h39 == parameter_2_2 ? phv_data_57 : _GEN_227; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_229 = 14'h3a == parameter_2_2 ? phv_data_58 : _GEN_228; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_230 = 14'h3b == parameter_2_2 ? phv_data_59 : _GEN_229; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_231 = 14'h3c == parameter_2_2 ? phv_data_60 : _GEN_230; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_232 = 14'h3d == parameter_2_2 ? phv_data_61 : _GEN_231; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_233 = 14'h3e == parameter_2_2 ? phv_data_62 : _GEN_232; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_234 = 14'h3f == parameter_2_2 ? phv_data_63 : _GEN_233; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_3 = vliw_3[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_3 = vliw_3[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_3 = parameter_2_3[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_3 = parameter_2_3[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_3 = {{1'd0}, args_offset_3}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_3 = _total_offset_T_3[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_238 = 3'h1 == total_offset_3 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_239 = 3'h2 == total_offset_3 ? args_2 : _GEN_238; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_240 = 3'h3 == total_offset_3 ? args_3 : _GEN_239; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_241 = 3'h4 == total_offset_3 ? args_4 : _GEN_240; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_242 = 3'h5 == total_offset_3 ? args_5 : _GEN_241; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_243 = 3'h6 == total_offset_3 ? args_6 : _GEN_242; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_244 = total_offset_3 < 3'h7 ? _GEN_243 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_3_0 = 3'h0 < args_length_3 ? _GEN_244 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_246 = opcode_3 == 4'ha ? field_bytes_3_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_247 = opcode_3 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_216 = opcode_3 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_7 = _T_216 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_248 = opcode_3 == 4'h8 | opcode_3 == 4'hb ? parameter_2_3[7:0] : _GEN_246; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_249 = opcode_3 == 4'h8 | opcode_3 == 4'hb ? _field_tag_T_7 : _GEN_247; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_250 = 14'h0 == parameter_2_3 ? phv_data_0 : _GEN_248; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_251 = 14'h1 == parameter_2_3 ? phv_data_1 : _GEN_250; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_252 = 14'h2 == parameter_2_3 ? phv_data_2 : _GEN_251; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_253 = 14'h3 == parameter_2_3 ? phv_data_3 : _GEN_252; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_254 = 14'h4 == parameter_2_3 ? phv_data_4 : _GEN_253; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_255 = 14'h5 == parameter_2_3 ? phv_data_5 : _GEN_254; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_256 = 14'h6 == parameter_2_3 ? phv_data_6 : _GEN_255; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_257 = 14'h7 == parameter_2_3 ? phv_data_7 : _GEN_256; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_258 = 14'h8 == parameter_2_3 ? phv_data_8 : _GEN_257; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_259 = 14'h9 == parameter_2_3 ? phv_data_9 : _GEN_258; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_260 = 14'ha == parameter_2_3 ? phv_data_10 : _GEN_259; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_261 = 14'hb == parameter_2_3 ? phv_data_11 : _GEN_260; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_262 = 14'hc == parameter_2_3 ? phv_data_12 : _GEN_261; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_263 = 14'hd == parameter_2_3 ? phv_data_13 : _GEN_262; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_264 = 14'he == parameter_2_3 ? phv_data_14 : _GEN_263; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_265 = 14'hf == parameter_2_3 ? phv_data_15 : _GEN_264; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_266 = 14'h10 == parameter_2_3 ? phv_data_16 : _GEN_265; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_267 = 14'h11 == parameter_2_3 ? phv_data_17 : _GEN_266; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_268 = 14'h12 == parameter_2_3 ? phv_data_18 : _GEN_267; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_269 = 14'h13 == parameter_2_3 ? phv_data_19 : _GEN_268; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_270 = 14'h14 == parameter_2_3 ? phv_data_20 : _GEN_269; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_271 = 14'h15 == parameter_2_3 ? phv_data_21 : _GEN_270; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_272 = 14'h16 == parameter_2_3 ? phv_data_22 : _GEN_271; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_273 = 14'h17 == parameter_2_3 ? phv_data_23 : _GEN_272; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_274 = 14'h18 == parameter_2_3 ? phv_data_24 : _GEN_273; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_275 = 14'h19 == parameter_2_3 ? phv_data_25 : _GEN_274; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_276 = 14'h1a == parameter_2_3 ? phv_data_26 : _GEN_275; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_277 = 14'h1b == parameter_2_3 ? phv_data_27 : _GEN_276; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_278 = 14'h1c == parameter_2_3 ? phv_data_28 : _GEN_277; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_279 = 14'h1d == parameter_2_3 ? phv_data_29 : _GEN_278; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_280 = 14'h1e == parameter_2_3 ? phv_data_30 : _GEN_279; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_281 = 14'h1f == parameter_2_3 ? phv_data_31 : _GEN_280; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_282 = 14'h20 == parameter_2_3 ? phv_data_32 : _GEN_281; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_283 = 14'h21 == parameter_2_3 ? phv_data_33 : _GEN_282; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_284 = 14'h22 == parameter_2_3 ? phv_data_34 : _GEN_283; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_285 = 14'h23 == parameter_2_3 ? phv_data_35 : _GEN_284; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_286 = 14'h24 == parameter_2_3 ? phv_data_36 : _GEN_285; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_287 = 14'h25 == parameter_2_3 ? phv_data_37 : _GEN_286; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_288 = 14'h26 == parameter_2_3 ? phv_data_38 : _GEN_287; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_289 = 14'h27 == parameter_2_3 ? phv_data_39 : _GEN_288; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_290 = 14'h28 == parameter_2_3 ? phv_data_40 : _GEN_289; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_291 = 14'h29 == parameter_2_3 ? phv_data_41 : _GEN_290; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_292 = 14'h2a == parameter_2_3 ? phv_data_42 : _GEN_291; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_293 = 14'h2b == parameter_2_3 ? phv_data_43 : _GEN_292; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_294 = 14'h2c == parameter_2_3 ? phv_data_44 : _GEN_293; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_295 = 14'h2d == parameter_2_3 ? phv_data_45 : _GEN_294; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_296 = 14'h2e == parameter_2_3 ? phv_data_46 : _GEN_295; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_297 = 14'h2f == parameter_2_3 ? phv_data_47 : _GEN_296; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_298 = 14'h30 == parameter_2_3 ? phv_data_48 : _GEN_297; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_299 = 14'h31 == parameter_2_3 ? phv_data_49 : _GEN_298; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_300 = 14'h32 == parameter_2_3 ? phv_data_50 : _GEN_299; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_301 = 14'h33 == parameter_2_3 ? phv_data_51 : _GEN_300; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_302 = 14'h34 == parameter_2_3 ? phv_data_52 : _GEN_301; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_303 = 14'h35 == parameter_2_3 ? phv_data_53 : _GEN_302; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_304 = 14'h36 == parameter_2_3 ? phv_data_54 : _GEN_303; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_305 = 14'h37 == parameter_2_3 ? phv_data_55 : _GEN_304; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_306 = 14'h38 == parameter_2_3 ? phv_data_56 : _GEN_305; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_307 = 14'h39 == parameter_2_3 ? phv_data_57 : _GEN_306; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_308 = 14'h3a == parameter_2_3 ? phv_data_58 : _GEN_307; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_309 = 14'h3b == parameter_2_3 ? phv_data_59 : _GEN_308; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_310 = 14'h3c == parameter_2_3 ? phv_data_60 : _GEN_309; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_311 = 14'h3d == parameter_2_3 ? phv_data_61 : _GEN_310; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_312 = 14'h3e == parameter_2_3 ? phv_data_62 : _GEN_311; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_313 = 14'h3f == parameter_2_3 ? phv_data_63 : _GEN_312; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_4 = vliw_4[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_4 = vliw_4[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_4 = parameter_2_4[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_4 = parameter_2_4[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_4 = {{1'd0}, args_offset_4}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_4 = _total_offset_T_4[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_317 = 3'h1 == total_offset_4 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_318 = 3'h2 == total_offset_4 ? args_2 : _GEN_317; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_319 = 3'h3 == total_offset_4 ? args_3 : _GEN_318; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_320 = 3'h4 == total_offset_4 ? args_4 : _GEN_319; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_321 = 3'h5 == total_offset_4 ? args_5 : _GEN_320; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_322 = 3'h6 == total_offset_4 ? args_6 : _GEN_321; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_323 = total_offset_4 < 3'h7 ? _GEN_322 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_4_0 = 3'h0 < args_length_4 ? _GEN_323 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_325 = opcode_4 == 4'ha ? field_bytes_4_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_326 = opcode_4 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_287 = opcode_4 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_9 = _T_287 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_327 = opcode_4 == 4'h8 | opcode_4 == 4'hb ? parameter_2_4[7:0] : _GEN_325; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_328 = opcode_4 == 4'h8 | opcode_4 == 4'hb ? _field_tag_T_9 : _GEN_326; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_329 = 14'h0 == parameter_2_4 ? phv_data_0 : _GEN_327; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_330 = 14'h1 == parameter_2_4 ? phv_data_1 : _GEN_329; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_331 = 14'h2 == parameter_2_4 ? phv_data_2 : _GEN_330; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_332 = 14'h3 == parameter_2_4 ? phv_data_3 : _GEN_331; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_333 = 14'h4 == parameter_2_4 ? phv_data_4 : _GEN_332; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_334 = 14'h5 == parameter_2_4 ? phv_data_5 : _GEN_333; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_335 = 14'h6 == parameter_2_4 ? phv_data_6 : _GEN_334; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_336 = 14'h7 == parameter_2_4 ? phv_data_7 : _GEN_335; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_337 = 14'h8 == parameter_2_4 ? phv_data_8 : _GEN_336; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_338 = 14'h9 == parameter_2_4 ? phv_data_9 : _GEN_337; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_339 = 14'ha == parameter_2_4 ? phv_data_10 : _GEN_338; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_340 = 14'hb == parameter_2_4 ? phv_data_11 : _GEN_339; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_341 = 14'hc == parameter_2_4 ? phv_data_12 : _GEN_340; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_342 = 14'hd == parameter_2_4 ? phv_data_13 : _GEN_341; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_343 = 14'he == parameter_2_4 ? phv_data_14 : _GEN_342; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_344 = 14'hf == parameter_2_4 ? phv_data_15 : _GEN_343; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_345 = 14'h10 == parameter_2_4 ? phv_data_16 : _GEN_344; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_346 = 14'h11 == parameter_2_4 ? phv_data_17 : _GEN_345; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_347 = 14'h12 == parameter_2_4 ? phv_data_18 : _GEN_346; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_348 = 14'h13 == parameter_2_4 ? phv_data_19 : _GEN_347; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_349 = 14'h14 == parameter_2_4 ? phv_data_20 : _GEN_348; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_350 = 14'h15 == parameter_2_4 ? phv_data_21 : _GEN_349; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_351 = 14'h16 == parameter_2_4 ? phv_data_22 : _GEN_350; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_352 = 14'h17 == parameter_2_4 ? phv_data_23 : _GEN_351; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_353 = 14'h18 == parameter_2_4 ? phv_data_24 : _GEN_352; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_354 = 14'h19 == parameter_2_4 ? phv_data_25 : _GEN_353; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_355 = 14'h1a == parameter_2_4 ? phv_data_26 : _GEN_354; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_356 = 14'h1b == parameter_2_4 ? phv_data_27 : _GEN_355; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_357 = 14'h1c == parameter_2_4 ? phv_data_28 : _GEN_356; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_358 = 14'h1d == parameter_2_4 ? phv_data_29 : _GEN_357; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_359 = 14'h1e == parameter_2_4 ? phv_data_30 : _GEN_358; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_360 = 14'h1f == parameter_2_4 ? phv_data_31 : _GEN_359; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_361 = 14'h20 == parameter_2_4 ? phv_data_32 : _GEN_360; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_362 = 14'h21 == parameter_2_4 ? phv_data_33 : _GEN_361; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_363 = 14'h22 == parameter_2_4 ? phv_data_34 : _GEN_362; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_364 = 14'h23 == parameter_2_4 ? phv_data_35 : _GEN_363; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_365 = 14'h24 == parameter_2_4 ? phv_data_36 : _GEN_364; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_366 = 14'h25 == parameter_2_4 ? phv_data_37 : _GEN_365; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_367 = 14'h26 == parameter_2_4 ? phv_data_38 : _GEN_366; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_368 = 14'h27 == parameter_2_4 ? phv_data_39 : _GEN_367; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_369 = 14'h28 == parameter_2_4 ? phv_data_40 : _GEN_368; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_370 = 14'h29 == parameter_2_4 ? phv_data_41 : _GEN_369; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_371 = 14'h2a == parameter_2_4 ? phv_data_42 : _GEN_370; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_372 = 14'h2b == parameter_2_4 ? phv_data_43 : _GEN_371; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_373 = 14'h2c == parameter_2_4 ? phv_data_44 : _GEN_372; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_374 = 14'h2d == parameter_2_4 ? phv_data_45 : _GEN_373; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_375 = 14'h2e == parameter_2_4 ? phv_data_46 : _GEN_374; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_376 = 14'h2f == parameter_2_4 ? phv_data_47 : _GEN_375; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_377 = 14'h30 == parameter_2_4 ? phv_data_48 : _GEN_376; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_378 = 14'h31 == parameter_2_4 ? phv_data_49 : _GEN_377; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_379 = 14'h32 == parameter_2_4 ? phv_data_50 : _GEN_378; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_380 = 14'h33 == parameter_2_4 ? phv_data_51 : _GEN_379; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_381 = 14'h34 == parameter_2_4 ? phv_data_52 : _GEN_380; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_382 = 14'h35 == parameter_2_4 ? phv_data_53 : _GEN_381; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_383 = 14'h36 == parameter_2_4 ? phv_data_54 : _GEN_382; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_384 = 14'h37 == parameter_2_4 ? phv_data_55 : _GEN_383; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_385 = 14'h38 == parameter_2_4 ? phv_data_56 : _GEN_384; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_386 = 14'h39 == parameter_2_4 ? phv_data_57 : _GEN_385; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_387 = 14'h3a == parameter_2_4 ? phv_data_58 : _GEN_386; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_388 = 14'h3b == parameter_2_4 ? phv_data_59 : _GEN_387; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_389 = 14'h3c == parameter_2_4 ? phv_data_60 : _GEN_388; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_390 = 14'h3d == parameter_2_4 ? phv_data_61 : _GEN_389; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_391 = 14'h3e == parameter_2_4 ? phv_data_62 : _GEN_390; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_392 = 14'h3f == parameter_2_4 ? phv_data_63 : _GEN_391; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_5 = vliw_5[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_5 = vliw_5[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_5 = parameter_2_5[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_5 = parameter_2_5[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_5 = {{1'd0}, args_offset_5}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_5 = _total_offset_T_5[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_396 = 3'h1 == total_offset_5 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_397 = 3'h2 == total_offset_5 ? args_2 : _GEN_396; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_398 = 3'h3 == total_offset_5 ? args_3 : _GEN_397; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_399 = 3'h4 == total_offset_5 ? args_4 : _GEN_398; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_400 = 3'h5 == total_offset_5 ? args_5 : _GEN_399; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_401 = 3'h6 == total_offset_5 ? args_6 : _GEN_400; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_402 = total_offset_5 < 3'h7 ? _GEN_401 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_5_0 = 3'h0 < args_length_5 ? _GEN_402 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_404 = opcode_5 == 4'ha ? field_bytes_5_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_405 = opcode_5 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_358 = opcode_5 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_11 = _T_358 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_406 = opcode_5 == 4'h8 | opcode_5 == 4'hb ? parameter_2_5[7:0] : _GEN_404; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_407 = opcode_5 == 4'h8 | opcode_5 == 4'hb ? _field_tag_T_11 : _GEN_405; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_408 = 14'h0 == parameter_2_5 ? phv_data_0 : _GEN_406; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_409 = 14'h1 == parameter_2_5 ? phv_data_1 : _GEN_408; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_410 = 14'h2 == parameter_2_5 ? phv_data_2 : _GEN_409; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_411 = 14'h3 == parameter_2_5 ? phv_data_3 : _GEN_410; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_412 = 14'h4 == parameter_2_5 ? phv_data_4 : _GEN_411; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_413 = 14'h5 == parameter_2_5 ? phv_data_5 : _GEN_412; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_414 = 14'h6 == parameter_2_5 ? phv_data_6 : _GEN_413; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_415 = 14'h7 == parameter_2_5 ? phv_data_7 : _GEN_414; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_416 = 14'h8 == parameter_2_5 ? phv_data_8 : _GEN_415; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_417 = 14'h9 == parameter_2_5 ? phv_data_9 : _GEN_416; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_418 = 14'ha == parameter_2_5 ? phv_data_10 : _GEN_417; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_419 = 14'hb == parameter_2_5 ? phv_data_11 : _GEN_418; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_420 = 14'hc == parameter_2_5 ? phv_data_12 : _GEN_419; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_421 = 14'hd == parameter_2_5 ? phv_data_13 : _GEN_420; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_422 = 14'he == parameter_2_5 ? phv_data_14 : _GEN_421; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_423 = 14'hf == parameter_2_5 ? phv_data_15 : _GEN_422; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_424 = 14'h10 == parameter_2_5 ? phv_data_16 : _GEN_423; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_425 = 14'h11 == parameter_2_5 ? phv_data_17 : _GEN_424; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_426 = 14'h12 == parameter_2_5 ? phv_data_18 : _GEN_425; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_427 = 14'h13 == parameter_2_5 ? phv_data_19 : _GEN_426; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_428 = 14'h14 == parameter_2_5 ? phv_data_20 : _GEN_427; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_429 = 14'h15 == parameter_2_5 ? phv_data_21 : _GEN_428; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_430 = 14'h16 == parameter_2_5 ? phv_data_22 : _GEN_429; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_431 = 14'h17 == parameter_2_5 ? phv_data_23 : _GEN_430; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_432 = 14'h18 == parameter_2_5 ? phv_data_24 : _GEN_431; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_433 = 14'h19 == parameter_2_5 ? phv_data_25 : _GEN_432; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_434 = 14'h1a == parameter_2_5 ? phv_data_26 : _GEN_433; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_435 = 14'h1b == parameter_2_5 ? phv_data_27 : _GEN_434; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_436 = 14'h1c == parameter_2_5 ? phv_data_28 : _GEN_435; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_437 = 14'h1d == parameter_2_5 ? phv_data_29 : _GEN_436; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_438 = 14'h1e == parameter_2_5 ? phv_data_30 : _GEN_437; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_439 = 14'h1f == parameter_2_5 ? phv_data_31 : _GEN_438; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_440 = 14'h20 == parameter_2_5 ? phv_data_32 : _GEN_439; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_441 = 14'h21 == parameter_2_5 ? phv_data_33 : _GEN_440; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_442 = 14'h22 == parameter_2_5 ? phv_data_34 : _GEN_441; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_443 = 14'h23 == parameter_2_5 ? phv_data_35 : _GEN_442; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_444 = 14'h24 == parameter_2_5 ? phv_data_36 : _GEN_443; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_445 = 14'h25 == parameter_2_5 ? phv_data_37 : _GEN_444; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_446 = 14'h26 == parameter_2_5 ? phv_data_38 : _GEN_445; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_447 = 14'h27 == parameter_2_5 ? phv_data_39 : _GEN_446; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_448 = 14'h28 == parameter_2_5 ? phv_data_40 : _GEN_447; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_449 = 14'h29 == parameter_2_5 ? phv_data_41 : _GEN_448; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_450 = 14'h2a == parameter_2_5 ? phv_data_42 : _GEN_449; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_451 = 14'h2b == parameter_2_5 ? phv_data_43 : _GEN_450; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_452 = 14'h2c == parameter_2_5 ? phv_data_44 : _GEN_451; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_453 = 14'h2d == parameter_2_5 ? phv_data_45 : _GEN_452; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_454 = 14'h2e == parameter_2_5 ? phv_data_46 : _GEN_453; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_455 = 14'h2f == parameter_2_5 ? phv_data_47 : _GEN_454; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_456 = 14'h30 == parameter_2_5 ? phv_data_48 : _GEN_455; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_457 = 14'h31 == parameter_2_5 ? phv_data_49 : _GEN_456; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_458 = 14'h32 == parameter_2_5 ? phv_data_50 : _GEN_457; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_459 = 14'h33 == parameter_2_5 ? phv_data_51 : _GEN_458; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_460 = 14'h34 == parameter_2_5 ? phv_data_52 : _GEN_459; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_461 = 14'h35 == parameter_2_5 ? phv_data_53 : _GEN_460; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_462 = 14'h36 == parameter_2_5 ? phv_data_54 : _GEN_461; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_463 = 14'h37 == parameter_2_5 ? phv_data_55 : _GEN_462; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_464 = 14'h38 == parameter_2_5 ? phv_data_56 : _GEN_463; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_465 = 14'h39 == parameter_2_5 ? phv_data_57 : _GEN_464; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_466 = 14'h3a == parameter_2_5 ? phv_data_58 : _GEN_465; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_467 = 14'h3b == parameter_2_5 ? phv_data_59 : _GEN_466; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_468 = 14'h3c == parameter_2_5 ? phv_data_60 : _GEN_467; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_469 = 14'h3d == parameter_2_5 ? phv_data_61 : _GEN_468; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_470 = 14'h3e == parameter_2_5 ? phv_data_62 : _GEN_469; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_471 = 14'h3f == parameter_2_5 ? phv_data_63 : _GEN_470; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_6 = vliw_6[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_6 = vliw_6[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_6 = parameter_2_6[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_6 = parameter_2_6[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_6 = {{1'd0}, args_offset_6}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_6 = _total_offset_T_6[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_475 = 3'h1 == total_offset_6 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_476 = 3'h2 == total_offset_6 ? args_2 : _GEN_475; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_477 = 3'h3 == total_offset_6 ? args_3 : _GEN_476; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_478 = 3'h4 == total_offset_6 ? args_4 : _GEN_477; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_479 = 3'h5 == total_offset_6 ? args_5 : _GEN_478; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_480 = 3'h6 == total_offset_6 ? args_6 : _GEN_479; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_481 = total_offset_6 < 3'h7 ? _GEN_480 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_6_0 = 3'h0 < args_length_6 ? _GEN_481 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_483 = opcode_6 == 4'ha ? field_bytes_6_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_484 = opcode_6 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_429 = opcode_6 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_13 = _T_429 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_485 = opcode_6 == 4'h8 | opcode_6 == 4'hb ? parameter_2_6[7:0] : _GEN_483; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_486 = opcode_6 == 4'h8 | opcode_6 == 4'hb ? _field_tag_T_13 : _GEN_484; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_487 = 14'h0 == parameter_2_6 ? phv_data_0 : _GEN_485; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_488 = 14'h1 == parameter_2_6 ? phv_data_1 : _GEN_487; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_489 = 14'h2 == parameter_2_6 ? phv_data_2 : _GEN_488; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_490 = 14'h3 == parameter_2_6 ? phv_data_3 : _GEN_489; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_491 = 14'h4 == parameter_2_6 ? phv_data_4 : _GEN_490; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_492 = 14'h5 == parameter_2_6 ? phv_data_5 : _GEN_491; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_493 = 14'h6 == parameter_2_6 ? phv_data_6 : _GEN_492; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_494 = 14'h7 == parameter_2_6 ? phv_data_7 : _GEN_493; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_495 = 14'h8 == parameter_2_6 ? phv_data_8 : _GEN_494; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_496 = 14'h9 == parameter_2_6 ? phv_data_9 : _GEN_495; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_497 = 14'ha == parameter_2_6 ? phv_data_10 : _GEN_496; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_498 = 14'hb == parameter_2_6 ? phv_data_11 : _GEN_497; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_499 = 14'hc == parameter_2_6 ? phv_data_12 : _GEN_498; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_500 = 14'hd == parameter_2_6 ? phv_data_13 : _GEN_499; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_501 = 14'he == parameter_2_6 ? phv_data_14 : _GEN_500; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_502 = 14'hf == parameter_2_6 ? phv_data_15 : _GEN_501; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_503 = 14'h10 == parameter_2_6 ? phv_data_16 : _GEN_502; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_504 = 14'h11 == parameter_2_6 ? phv_data_17 : _GEN_503; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_505 = 14'h12 == parameter_2_6 ? phv_data_18 : _GEN_504; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_506 = 14'h13 == parameter_2_6 ? phv_data_19 : _GEN_505; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_507 = 14'h14 == parameter_2_6 ? phv_data_20 : _GEN_506; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_508 = 14'h15 == parameter_2_6 ? phv_data_21 : _GEN_507; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_509 = 14'h16 == parameter_2_6 ? phv_data_22 : _GEN_508; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_510 = 14'h17 == parameter_2_6 ? phv_data_23 : _GEN_509; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_511 = 14'h18 == parameter_2_6 ? phv_data_24 : _GEN_510; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_512 = 14'h19 == parameter_2_6 ? phv_data_25 : _GEN_511; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_513 = 14'h1a == parameter_2_6 ? phv_data_26 : _GEN_512; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_514 = 14'h1b == parameter_2_6 ? phv_data_27 : _GEN_513; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_515 = 14'h1c == parameter_2_6 ? phv_data_28 : _GEN_514; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_516 = 14'h1d == parameter_2_6 ? phv_data_29 : _GEN_515; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_517 = 14'h1e == parameter_2_6 ? phv_data_30 : _GEN_516; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_518 = 14'h1f == parameter_2_6 ? phv_data_31 : _GEN_517; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_519 = 14'h20 == parameter_2_6 ? phv_data_32 : _GEN_518; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_520 = 14'h21 == parameter_2_6 ? phv_data_33 : _GEN_519; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_521 = 14'h22 == parameter_2_6 ? phv_data_34 : _GEN_520; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_522 = 14'h23 == parameter_2_6 ? phv_data_35 : _GEN_521; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_523 = 14'h24 == parameter_2_6 ? phv_data_36 : _GEN_522; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_524 = 14'h25 == parameter_2_6 ? phv_data_37 : _GEN_523; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_525 = 14'h26 == parameter_2_6 ? phv_data_38 : _GEN_524; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_526 = 14'h27 == parameter_2_6 ? phv_data_39 : _GEN_525; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_527 = 14'h28 == parameter_2_6 ? phv_data_40 : _GEN_526; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_528 = 14'h29 == parameter_2_6 ? phv_data_41 : _GEN_527; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_529 = 14'h2a == parameter_2_6 ? phv_data_42 : _GEN_528; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_530 = 14'h2b == parameter_2_6 ? phv_data_43 : _GEN_529; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_531 = 14'h2c == parameter_2_6 ? phv_data_44 : _GEN_530; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_532 = 14'h2d == parameter_2_6 ? phv_data_45 : _GEN_531; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_533 = 14'h2e == parameter_2_6 ? phv_data_46 : _GEN_532; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_534 = 14'h2f == parameter_2_6 ? phv_data_47 : _GEN_533; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_535 = 14'h30 == parameter_2_6 ? phv_data_48 : _GEN_534; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_536 = 14'h31 == parameter_2_6 ? phv_data_49 : _GEN_535; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_537 = 14'h32 == parameter_2_6 ? phv_data_50 : _GEN_536; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_538 = 14'h33 == parameter_2_6 ? phv_data_51 : _GEN_537; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_539 = 14'h34 == parameter_2_6 ? phv_data_52 : _GEN_538; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_540 = 14'h35 == parameter_2_6 ? phv_data_53 : _GEN_539; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_541 = 14'h36 == parameter_2_6 ? phv_data_54 : _GEN_540; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_542 = 14'h37 == parameter_2_6 ? phv_data_55 : _GEN_541; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_543 = 14'h38 == parameter_2_6 ? phv_data_56 : _GEN_542; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_544 = 14'h39 == parameter_2_6 ? phv_data_57 : _GEN_543; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_545 = 14'h3a == parameter_2_6 ? phv_data_58 : _GEN_544; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_546 = 14'h3b == parameter_2_6 ? phv_data_59 : _GEN_545; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_547 = 14'h3c == parameter_2_6 ? phv_data_60 : _GEN_546; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_548 = 14'h3d == parameter_2_6 ? phv_data_61 : _GEN_547; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_549 = 14'h3e == parameter_2_6 ? phv_data_62 : _GEN_548; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_550 = 14'h3f == parameter_2_6 ? phv_data_63 : _GEN_549; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_7 = vliw_7[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_7 = vliw_7[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_7 = parameter_2_7[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_7 = parameter_2_7[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_7 = {{1'd0}, args_offset_7}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_7 = _total_offset_T_7[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_554 = 3'h1 == total_offset_7 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_555 = 3'h2 == total_offset_7 ? args_2 : _GEN_554; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_556 = 3'h3 == total_offset_7 ? args_3 : _GEN_555; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_557 = 3'h4 == total_offset_7 ? args_4 : _GEN_556; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_558 = 3'h5 == total_offset_7 ? args_5 : _GEN_557; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_559 = 3'h6 == total_offset_7 ? args_6 : _GEN_558; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_560 = total_offset_7 < 3'h7 ? _GEN_559 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_7_0 = 3'h0 < args_length_7 ? _GEN_560 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_562 = opcode_7 == 4'ha ? field_bytes_7_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_563 = opcode_7 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_500 = opcode_7 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_15 = _T_500 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_564 = opcode_7 == 4'h8 | opcode_7 == 4'hb ? parameter_2_7[7:0] : _GEN_562; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_565 = opcode_7 == 4'h8 | opcode_7 == 4'hb ? _field_tag_T_15 : _GEN_563; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_566 = 14'h0 == parameter_2_7 ? phv_data_0 : _GEN_564; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_567 = 14'h1 == parameter_2_7 ? phv_data_1 : _GEN_566; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_568 = 14'h2 == parameter_2_7 ? phv_data_2 : _GEN_567; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_569 = 14'h3 == parameter_2_7 ? phv_data_3 : _GEN_568; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_570 = 14'h4 == parameter_2_7 ? phv_data_4 : _GEN_569; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_571 = 14'h5 == parameter_2_7 ? phv_data_5 : _GEN_570; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_572 = 14'h6 == parameter_2_7 ? phv_data_6 : _GEN_571; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_573 = 14'h7 == parameter_2_7 ? phv_data_7 : _GEN_572; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_574 = 14'h8 == parameter_2_7 ? phv_data_8 : _GEN_573; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_575 = 14'h9 == parameter_2_7 ? phv_data_9 : _GEN_574; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_576 = 14'ha == parameter_2_7 ? phv_data_10 : _GEN_575; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_577 = 14'hb == parameter_2_7 ? phv_data_11 : _GEN_576; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_578 = 14'hc == parameter_2_7 ? phv_data_12 : _GEN_577; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_579 = 14'hd == parameter_2_7 ? phv_data_13 : _GEN_578; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_580 = 14'he == parameter_2_7 ? phv_data_14 : _GEN_579; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_581 = 14'hf == parameter_2_7 ? phv_data_15 : _GEN_580; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_582 = 14'h10 == parameter_2_7 ? phv_data_16 : _GEN_581; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_583 = 14'h11 == parameter_2_7 ? phv_data_17 : _GEN_582; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_584 = 14'h12 == parameter_2_7 ? phv_data_18 : _GEN_583; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_585 = 14'h13 == parameter_2_7 ? phv_data_19 : _GEN_584; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_586 = 14'h14 == parameter_2_7 ? phv_data_20 : _GEN_585; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_587 = 14'h15 == parameter_2_7 ? phv_data_21 : _GEN_586; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_588 = 14'h16 == parameter_2_7 ? phv_data_22 : _GEN_587; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_589 = 14'h17 == parameter_2_7 ? phv_data_23 : _GEN_588; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_590 = 14'h18 == parameter_2_7 ? phv_data_24 : _GEN_589; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_591 = 14'h19 == parameter_2_7 ? phv_data_25 : _GEN_590; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_592 = 14'h1a == parameter_2_7 ? phv_data_26 : _GEN_591; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_593 = 14'h1b == parameter_2_7 ? phv_data_27 : _GEN_592; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_594 = 14'h1c == parameter_2_7 ? phv_data_28 : _GEN_593; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_595 = 14'h1d == parameter_2_7 ? phv_data_29 : _GEN_594; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_596 = 14'h1e == parameter_2_7 ? phv_data_30 : _GEN_595; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_597 = 14'h1f == parameter_2_7 ? phv_data_31 : _GEN_596; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_598 = 14'h20 == parameter_2_7 ? phv_data_32 : _GEN_597; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_599 = 14'h21 == parameter_2_7 ? phv_data_33 : _GEN_598; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_600 = 14'h22 == parameter_2_7 ? phv_data_34 : _GEN_599; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_601 = 14'h23 == parameter_2_7 ? phv_data_35 : _GEN_600; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_602 = 14'h24 == parameter_2_7 ? phv_data_36 : _GEN_601; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_603 = 14'h25 == parameter_2_7 ? phv_data_37 : _GEN_602; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_604 = 14'h26 == parameter_2_7 ? phv_data_38 : _GEN_603; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_605 = 14'h27 == parameter_2_7 ? phv_data_39 : _GEN_604; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_606 = 14'h28 == parameter_2_7 ? phv_data_40 : _GEN_605; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_607 = 14'h29 == parameter_2_7 ? phv_data_41 : _GEN_606; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_608 = 14'h2a == parameter_2_7 ? phv_data_42 : _GEN_607; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_609 = 14'h2b == parameter_2_7 ? phv_data_43 : _GEN_608; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_610 = 14'h2c == parameter_2_7 ? phv_data_44 : _GEN_609; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_611 = 14'h2d == parameter_2_7 ? phv_data_45 : _GEN_610; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_612 = 14'h2e == parameter_2_7 ? phv_data_46 : _GEN_611; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_613 = 14'h2f == parameter_2_7 ? phv_data_47 : _GEN_612; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_614 = 14'h30 == parameter_2_7 ? phv_data_48 : _GEN_613; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_615 = 14'h31 == parameter_2_7 ? phv_data_49 : _GEN_614; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_616 = 14'h32 == parameter_2_7 ? phv_data_50 : _GEN_615; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_617 = 14'h33 == parameter_2_7 ? phv_data_51 : _GEN_616; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_618 = 14'h34 == parameter_2_7 ? phv_data_52 : _GEN_617; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_619 = 14'h35 == parameter_2_7 ? phv_data_53 : _GEN_618; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_620 = 14'h36 == parameter_2_7 ? phv_data_54 : _GEN_619; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_621 = 14'h37 == parameter_2_7 ? phv_data_55 : _GEN_620; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_622 = 14'h38 == parameter_2_7 ? phv_data_56 : _GEN_621; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_623 = 14'h39 == parameter_2_7 ? phv_data_57 : _GEN_622; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_624 = 14'h3a == parameter_2_7 ? phv_data_58 : _GEN_623; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_625 = 14'h3b == parameter_2_7 ? phv_data_59 : _GEN_624; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_626 = 14'h3c == parameter_2_7 ? phv_data_60 : _GEN_625; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_627 = 14'h3d == parameter_2_7 ? phv_data_61 : _GEN_626; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_628 = 14'h3e == parameter_2_7 ? phv_data_62 : _GEN_627; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_629 = 14'h3f == parameter_2_7 ? phv_data_63 : _GEN_628; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_8 = vliw_8[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_8 = vliw_8[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_8 = parameter_2_8[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_8 = parameter_2_8[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_8 = {{1'd0}, args_offset_8}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_8 = _total_offset_T_8[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_633 = 3'h1 == total_offset_8 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_634 = 3'h2 == total_offset_8 ? args_2 : _GEN_633; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_635 = 3'h3 == total_offset_8 ? args_3 : _GEN_634; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_636 = 3'h4 == total_offset_8 ? args_4 : _GEN_635; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_637 = 3'h5 == total_offset_8 ? args_5 : _GEN_636; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_638 = 3'h6 == total_offset_8 ? args_6 : _GEN_637; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_639 = total_offset_8 < 3'h7 ? _GEN_638 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_8_0 = 3'h0 < args_length_8 ? _GEN_639 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_641 = opcode_8 == 4'ha ? field_bytes_8_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_642 = opcode_8 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_571 = opcode_8 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_17 = _T_571 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_643 = opcode_8 == 4'h8 | opcode_8 == 4'hb ? parameter_2_8[7:0] : _GEN_641; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_644 = opcode_8 == 4'h8 | opcode_8 == 4'hb ? _field_tag_T_17 : _GEN_642; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_645 = 14'h0 == parameter_2_8 ? phv_data_0 : _GEN_643; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_646 = 14'h1 == parameter_2_8 ? phv_data_1 : _GEN_645; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_647 = 14'h2 == parameter_2_8 ? phv_data_2 : _GEN_646; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_648 = 14'h3 == parameter_2_8 ? phv_data_3 : _GEN_647; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_649 = 14'h4 == parameter_2_8 ? phv_data_4 : _GEN_648; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_650 = 14'h5 == parameter_2_8 ? phv_data_5 : _GEN_649; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_651 = 14'h6 == parameter_2_8 ? phv_data_6 : _GEN_650; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_652 = 14'h7 == parameter_2_8 ? phv_data_7 : _GEN_651; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_653 = 14'h8 == parameter_2_8 ? phv_data_8 : _GEN_652; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_654 = 14'h9 == parameter_2_8 ? phv_data_9 : _GEN_653; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_655 = 14'ha == parameter_2_8 ? phv_data_10 : _GEN_654; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_656 = 14'hb == parameter_2_8 ? phv_data_11 : _GEN_655; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_657 = 14'hc == parameter_2_8 ? phv_data_12 : _GEN_656; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_658 = 14'hd == parameter_2_8 ? phv_data_13 : _GEN_657; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_659 = 14'he == parameter_2_8 ? phv_data_14 : _GEN_658; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_660 = 14'hf == parameter_2_8 ? phv_data_15 : _GEN_659; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_661 = 14'h10 == parameter_2_8 ? phv_data_16 : _GEN_660; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_662 = 14'h11 == parameter_2_8 ? phv_data_17 : _GEN_661; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_663 = 14'h12 == parameter_2_8 ? phv_data_18 : _GEN_662; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_664 = 14'h13 == parameter_2_8 ? phv_data_19 : _GEN_663; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_665 = 14'h14 == parameter_2_8 ? phv_data_20 : _GEN_664; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_666 = 14'h15 == parameter_2_8 ? phv_data_21 : _GEN_665; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_667 = 14'h16 == parameter_2_8 ? phv_data_22 : _GEN_666; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_668 = 14'h17 == parameter_2_8 ? phv_data_23 : _GEN_667; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_669 = 14'h18 == parameter_2_8 ? phv_data_24 : _GEN_668; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_670 = 14'h19 == parameter_2_8 ? phv_data_25 : _GEN_669; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_671 = 14'h1a == parameter_2_8 ? phv_data_26 : _GEN_670; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_672 = 14'h1b == parameter_2_8 ? phv_data_27 : _GEN_671; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_673 = 14'h1c == parameter_2_8 ? phv_data_28 : _GEN_672; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_674 = 14'h1d == parameter_2_8 ? phv_data_29 : _GEN_673; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_675 = 14'h1e == parameter_2_8 ? phv_data_30 : _GEN_674; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_676 = 14'h1f == parameter_2_8 ? phv_data_31 : _GEN_675; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_677 = 14'h20 == parameter_2_8 ? phv_data_32 : _GEN_676; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_678 = 14'h21 == parameter_2_8 ? phv_data_33 : _GEN_677; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_679 = 14'h22 == parameter_2_8 ? phv_data_34 : _GEN_678; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_680 = 14'h23 == parameter_2_8 ? phv_data_35 : _GEN_679; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_681 = 14'h24 == parameter_2_8 ? phv_data_36 : _GEN_680; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_682 = 14'h25 == parameter_2_8 ? phv_data_37 : _GEN_681; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_683 = 14'h26 == parameter_2_8 ? phv_data_38 : _GEN_682; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_684 = 14'h27 == parameter_2_8 ? phv_data_39 : _GEN_683; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_685 = 14'h28 == parameter_2_8 ? phv_data_40 : _GEN_684; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_686 = 14'h29 == parameter_2_8 ? phv_data_41 : _GEN_685; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_687 = 14'h2a == parameter_2_8 ? phv_data_42 : _GEN_686; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_688 = 14'h2b == parameter_2_8 ? phv_data_43 : _GEN_687; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_689 = 14'h2c == parameter_2_8 ? phv_data_44 : _GEN_688; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_690 = 14'h2d == parameter_2_8 ? phv_data_45 : _GEN_689; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_691 = 14'h2e == parameter_2_8 ? phv_data_46 : _GEN_690; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_692 = 14'h2f == parameter_2_8 ? phv_data_47 : _GEN_691; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_693 = 14'h30 == parameter_2_8 ? phv_data_48 : _GEN_692; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_694 = 14'h31 == parameter_2_8 ? phv_data_49 : _GEN_693; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_695 = 14'h32 == parameter_2_8 ? phv_data_50 : _GEN_694; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_696 = 14'h33 == parameter_2_8 ? phv_data_51 : _GEN_695; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_697 = 14'h34 == parameter_2_8 ? phv_data_52 : _GEN_696; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_698 = 14'h35 == parameter_2_8 ? phv_data_53 : _GEN_697; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_699 = 14'h36 == parameter_2_8 ? phv_data_54 : _GEN_698; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_700 = 14'h37 == parameter_2_8 ? phv_data_55 : _GEN_699; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_701 = 14'h38 == parameter_2_8 ? phv_data_56 : _GEN_700; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_702 = 14'h39 == parameter_2_8 ? phv_data_57 : _GEN_701; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_703 = 14'h3a == parameter_2_8 ? phv_data_58 : _GEN_702; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_704 = 14'h3b == parameter_2_8 ? phv_data_59 : _GEN_703; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_705 = 14'h3c == parameter_2_8 ? phv_data_60 : _GEN_704; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_706 = 14'h3d == parameter_2_8 ? phv_data_61 : _GEN_705; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_707 = 14'h3e == parameter_2_8 ? phv_data_62 : _GEN_706; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_708 = 14'h3f == parameter_2_8 ? phv_data_63 : _GEN_707; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_9 = vliw_9[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_9 = vliw_9[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_9 = parameter_2_9[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_9 = parameter_2_9[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_9 = {{1'd0}, args_offset_9}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_9 = _total_offset_T_9[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_712 = 3'h1 == total_offset_9 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_713 = 3'h2 == total_offset_9 ? args_2 : _GEN_712; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_714 = 3'h3 == total_offset_9 ? args_3 : _GEN_713; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_715 = 3'h4 == total_offset_9 ? args_4 : _GEN_714; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_716 = 3'h5 == total_offset_9 ? args_5 : _GEN_715; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_717 = 3'h6 == total_offset_9 ? args_6 : _GEN_716; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_718 = total_offset_9 < 3'h7 ? _GEN_717 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_9_0 = 3'h0 < args_length_9 ? _GEN_718 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_720 = opcode_9 == 4'ha ? field_bytes_9_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_721 = opcode_9 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_642 = opcode_9 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_19 = _T_642 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_722 = opcode_9 == 4'h8 | opcode_9 == 4'hb ? parameter_2_9[7:0] : _GEN_720; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_723 = opcode_9 == 4'h8 | opcode_9 == 4'hb ? _field_tag_T_19 : _GEN_721; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_724 = 14'h0 == parameter_2_9 ? phv_data_0 : _GEN_722; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_725 = 14'h1 == parameter_2_9 ? phv_data_1 : _GEN_724; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_726 = 14'h2 == parameter_2_9 ? phv_data_2 : _GEN_725; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_727 = 14'h3 == parameter_2_9 ? phv_data_3 : _GEN_726; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_728 = 14'h4 == parameter_2_9 ? phv_data_4 : _GEN_727; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_729 = 14'h5 == parameter_2_9 ? phv_data_5 : _GEN_728; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_730 = 14'h6 == parameter_2_9 ? phv_data_6 : _GEN_729; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_731 = 14'h7 == parameter_2_9 ? phv_data_7 : _GEN_730; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_732 = 14'h8 == parameter_2_9 ? phv_data_8 : _GEN_731; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_733 = 14'h9 == parameter_2_9 ? phv_data_9 : _GEN_732; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_734 = 14'ha == parameter_2_9 ? phv_data_10 : _GEN_733; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_735 = 14'hb == parameter_2_9 ? phv_data_11 : _GEN_734; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_736 = 14'hc == parameter_2_9 ? phv_data_12 : _GEN_735; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_737 = 14'hd == parameter_2_9 ? phv_data_13 : _GEN_736; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_738 = 14'he == parameter_2_9 ? phv_data_14 : _GEN_737; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_739 = 14'hf == parameter_2_9 ? phv_data_15 : _GEN_738; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_740 = 14'h10 == parameter_2_9 ? phv_data_16 : _GEN_739; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_741 = 14'h11 == parameter_2_9 ? phv_data_17 : _GEN_740; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_742 = 14'h12 == parameter_2_9 ? phv_data_18 : _GEN_741; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_743 = 14'h13 == parameter_2_9 ? phv_data_19 : _GEN_742; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_744 = 14'h14 == parameter_2_9 ? phv_data_20 : _GEN_743; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_745 = 14'h15 == parameter_2_9 ? phv_data_21 : _GEN_744; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_746 = 14'h16 == parameter_2_9 ? phv_data_22 : _GEN_745; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_747 = 14'h17 == parameter_2_9 ? phv_data_23 : _GEN_746; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_748 = 14'h18 == parameter_2_9 ? phv_data_24 : _GEN_747; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_749 = 14'h19 == parameter_2_9 ? phv_data_25 : _GEN_748; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_750 = 14'h1a == parameter_2_9 ? phv_data_26 : _GEN_749; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_751 = 14'h1b == parameter_2_9 ? phv_data_27 : _GEN_750; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_752 = 14'h1c == parameter_2_9 ? phv_data_28 : _GEN_751; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_753 = 14'h1d == parameter_2_9 ? phv_data_29 : _GEN_752; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_754 = 14'h1e == parameter_2_9 ? phv_data_30 : _GEN_753; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_755 = 14'h1f == parameter_2_9 ? phv_data_31 : _GEN_754; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_756 = 14'h20 == parameter_2_9 ? phv_data_32 : _GEN_755; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_757 = 14'h21 == parameter_2_9 ? phv_data_33 : _GEN_756; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_758 = 14'h22 == parameter_2_9 ? phv_data_34 : _GEN_757; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_759 = 14'h23 == parameter_2_9 ? phv_data_35 : _GEN_758; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_760 = 14'h24 == parameter_2_9 ? phv_data_36 : _GEN_759; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_761 = 14'h25 == parameter_2_9 ? phv_data_37 : _GEN_760; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_762 = 14'h26 == parameter_2_9 ? phv_data_38 : _GEN_761; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_763 = 14'h27 == parameter_2_9 ? phv_data_39 : _GEN_762; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_764 = 14'h28 == parameter_2_9 ? phv_data_40 : _GEN_763; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_765 = 14'h29 == parameter_2_9 ? phv_data_41 : _GEN_764; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_766 = 14'h2a == parameter_2_9 ? phv_data_42 : _GEN_765; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_767 = 14'h2b == parameter_2_9 ? phv_data_43 : _GEN_766; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_768 = 14'h2c == parameter_2_9 ? phv_data_44 : _GEN_767; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_769 = 14'h2d == parameter_2_9 ? phv_data_45 : _GEN_768; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_770 = 14'h2e == parameter_2_9 ? phv_data_46 : _GEN_769; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_771 = 14'h2f == parameter_2_9 ? phv_data_47 : _GEN_770; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_772 = 14'h30 == parameter_2_9 ? phv_data_48 : _GEN_771; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_773 = 14'h31 == parameter_2_9 ? phv_data_49 : _GEN_772; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_774 = 14'h32 == parameter_2_9 ? phv_data_50 : _GEN_773; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_775 = 14'h33 == parameter_2_9 ? phv_data_51 : _GEN_774; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_776 = 14'h34 == parameter_2_9 ? phv_data_52 : _GEN_775; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_777 = 14'h35 == parameter_2_9 ? phv_data_53 : _GEN_776; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_778 = 14'h36 == parameter_2_9 ? phv_data_54 : _GEN_777; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_779 = 14'h37 == parameter_2_9 ? phv_data_55 : _GEN_778; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_780 = 14'h38 == parameter_2_9 ? phv_data_56 : _GEN_779; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_781 = 14'h39 == parameter_2_9 ? phv_data_57 : _GEN_780; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_782 = 14'h3a == parameter_2_9 ? phv_data_58 : _GEN_781; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_783 = 14'h3b == parameter_2_9 ? phv_data_59 : _GEN_782; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_784 = 14'h3c == parameter_2_9 ? phv_data_60 : _GEN_783; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_785 = 14'h3d == parameter_2_9 ? phv_data_61 : _GEN_784; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_786 = 14'h3e == parameter_2_9 ? phv_data_62 : _GEN_785; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_787 = 14'h3f == parameter_2_9 ? phv_data_63 : _GEN_786; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_10 = vliw_10[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_10 = vliw_10[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_10 = parameter_2_10[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_10 = parameter_2_10[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_10 = {{1'd0}, args_offset_10}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_10 = _total_offset_T_10[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_791 = 3'h1 == total_offset_10 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_792 = 3'h2 == total_offset_10 ? args_2 : _GEN_791; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_793 = 3'h3 == total_offset_10 ? args_3 : _GEN_792; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_794 = 3'h4 == total_offset_10 ? args_4 : _GEN_793; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_795 = 3'h5 == total_offset_10 ? args_5 : _GEN_794; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_796 = 3'h6 == total_offset_10 ? args_6 : _GEN_795; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_797 = total_offset_10 < 3'h7 ? _GEN_796 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_10_0 = 3'h0 < args_length_10 ? _GEN_797 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_799 = opcode_10 == 4'ha ? field_bytes_10_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_800 = opcode_10 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_713 = opcode_10 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_21 = _T_713 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_801 = opcode_10 == 4'h8 | opcode_10 == 4'hb ? parameter_2_10[7:0] : _GEN_799; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_802 = opcode_10 == 4'h8 | opcode_10 == 4'hb ? _field_tag_T_21 : _GEN_800; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_803 = 14'h0 == parameter_2_10 ? phv_data_0 : _GEN_801; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_804 = 14'h1 == parameter_2_10 ? phv_data_1 : _GEN_803; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_805 = 14'h2 == parameter_2_10 ? phv_data_2 : _GEN_804; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_806 = 14'h3 == parameter_2_10 ? phv_data_3 : _GEN_805; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_807 = 14'h4 == parameter_2_10 ? phv_data_4 : _GEN_806; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_808 = 14'h5 == parameter_2_10 ? phv_data_5 : _GEN_807; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_809 = 14'h6 == parameter_2_10 ? phv_data_6 : _GEN_808; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_810 = 14'h7 == parameter_2_10 ? phv_data_7 : _GEN_809; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_811 = 14'h8 == parameter_2_10 ? phv_data_8 : _GEN_810; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_812 = 14'h9 == parameter_2_10 ? phv_data_9 : _GEN_811; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_813 = 14'ha == parameter_2_10 ? phv_data_10 : _GEN_812; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_814 = 14'hb == parameter_2_10 ? phv_data_11 : _GEN_813; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_815 = 14'hc == parameter_2_10 ? phv_data_12 : _GEN_814; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_816 = 14'hd == parameter_2_10 ? phv_data_13 : _GEN_815; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_817 = 14'he == parameter_2_10 ? phv_data_14 : _GEN_816; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_818 = 14'hf == parameter_2_10 ? phv_data_15 : _GEN_817; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_819 = 14'h10 == parameter_2_10 ? phv_data_16 : _GEN_818; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_820 = 14'h11 == parameter_2_10 ? phv_data_17 : _GEN_819; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_821 = 14'h12 == parameter_2_10 ? phv_data_18 : _GEN_820; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_822 = 14'h13 == parameter_2_10 ? phv_data_19 : _GEN_821; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_823 = 14'h14 == parameter_2_10 ? phv_data_20 : _GEN_822; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_824 = 14'h15 == parameter_2_10 ? phv_data_21 : _GEN_823; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_825 = 14'h16 == parameter_2_10 ? phv_data_22 : _GEN_824; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_826 = 14'h17 == parameter_2_10 ? phv_data_23 : _GEN_825; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_827 = 14'h18 == parameter_2_10 ? phv_data_24 : _GEN_826; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_828 = 14'h19 == parameter_2_10 ? phv_data_25 : _GEN_827; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_829 = 14'h1a == parameter_2_10 ? phv_data_26 : _GEN_828; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_830 = 14'h1b == parameter_2_10 ? phv_data_27 : _GEN_829; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_831 = 14'h1c == parameter_2_10 ? phv_data_28 : _GEN_830; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_832 = 14'h1d == parameter_2_10 ? phv_data_29 : _GEN_831; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_833 = 14'h1e == parameter_2_10 ? phv_data_30 : _GEN_832; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_834 = 14'h1f == parameter_2_10 ? phv_data_31 : _GEN_833; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_835 = 14'h20 == parameter_2_10 ? phv_data_32 : _GEN_834; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_836 = 14'h21 == parameter_2_10 ? phv_data_33 : _GEN_835; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_837 = 14'h22 == parameter_2_10 ? phv_data_34 : _GEN_836; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_838 = 14'h23 == parameter_2_10 ? phv_data_35 : _GEN_837; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_839 = 14'h24 == parameter_2_10 ? phv_data_36 : _GEN_838; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_840 = 14'h25 == parameter_2_10 ? phv_data_37 : _GEN_839; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_841 = 14'h26 == parameter_2_10 ? phv_data_38 : _GEN_840; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_842 = 14'h27 == parameter_2_10 ? phv_data_39 : _GEN_841; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_843 = 14'h28 == parameter_2_10 ? phv_data_40 : _GEN_842; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_844 = 14'h29 == parameter_2_10 ? phv_data_41 : _GEN_843; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_845 = 14'h2a == parameter_2_10 ? phv_data_42 : _GEN_844; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_846 = 14'h2b == parameter_2_10 ? phv_data_43 : _GEN_845; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_847 = 14'h2c == parameter_2_10 ? phv_data_44 : _GEN_846; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_848 = 14'h2d == parameter_2_10 ? phv_data_45 : _GEN_847; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_849 = 14'h2e == parameter_2_10 ? phv_data_46 : _GEN_848; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_850 = 14'h2f == parameter_2_10 ? phv_data_47 : _GEN_849; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_851 = 14'h30 == parameter_2_10 ? phv_data_48 : _GEN_850; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_852 = 14'h31 == parameter_2_10 ? phv_data_49 : _GEN_851; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_853 = 14'h32 == parameter_2_10 ? phv_data_50 : _GEN_852; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_854 = 14'h33 == parameter_2_10 ? phv_data_51 : _GEN_853; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_855 = 14'h34 == parameter_2_10 ? phv_data_52 : _GEN_854; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_856 = 14'h35 == parameter_2_10 ? phv_data_53 : _GEN_855; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_857 = 14'h36 == parameter_2_10 ? phv_data_54 : _GEN_856; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_858 = 14'h37 == parameter_2_10 ? phv_data_55 : _GEN_857; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_859 = 14'h38 == parameter_2_10 ? phv_data_56 : _GEN_858; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_860 = 14'h39 == parameter_2_10 ? phv_data_57 : _GEN_859; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_861 = 14'h3a == parameter_2_10 ? phv_data_58 : _GEN_860; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_862 = 14'h3b == parameter_2_10 ? phv_data_59 : _GEN_861; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_863 = 14'h3c == parameter_2_10 ? phv_data_60 : _GEN_862; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_864 = 14'h3d == parameter_2_10 ? phv_data_61 : _GEN_863; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_865 = 14'h3e == parameter_2_10 ? phv_data_62 : _GEN_864; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_866 = 14'h3f == parameter_2_10 ? phv_data_63 : _GEN_865; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_11 = vliw_11[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_11 = vliw_11[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_11 = parameter_2_11[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_11 = parameter_2_11[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_11 = {{1'd0}, args_offset_11}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_11 = _total_offset_T_11[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_870 = 3'h1 == total_offset_11 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_871 = 3'h2 == total_offset_11 ? args_2 : _GEN_870; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_872 = 3'h3 == total_offset_11 ? args_3 : _GEN_871; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_873 = 3'h4 == total_offset_11 ? args_4 : _GEN_872; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_874 = 3'h5 == total_offset_11 ? args_5 : _GEN_873; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_875 = 3'h6 == total_offset_11 ? args_6 : _GEN_874; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_876 = total_offset_11 < 3'h7 ? _GEN_875 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_11_0 = 3'h0 < args_length_11 ? _GEN_876 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_878 = opcode_11 == 4'ha ? field_bytes_11_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_879 = opcode_11 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_784 = opcode_11 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_23 = _T_784 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_880 = opcode_11 == 4'h8 | opcode_11 == 4'hb ? parameter_2_11[7:0] : _GEN_878; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_881 = opcode_11 == 4'h8 | opcode_11 == 4'hb ? _field_tag_T_23 : _GEN_879; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_882 = 14'h0 == parameter_2_11 ? phv_data_0 : _GEN_880; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_883 = 14'h1 == parameter_2_11 ? phv_data_1 : _GEN_882; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_884 = 14'h2 == parameter_2_11 ? phv_data_2 : _GEN_883; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_885 = 14'h3 == parameter_2_11 ? phv_data_3 : _GEN_884; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_886 = 14'h4 == parameter_2_11 ? phv_data_4 : _GEN_885; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_887 = 14'h5 == parameter_2_11 ? phv_data_5 : _GEN_886; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_888 = 14'h6 == parameter_2_11 ? phv_data_6 : _GEN_887; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_889 = 14'h7 == parameter_2_11 ? phv_data_7 : _GEN_888; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_890 = 14'h8 == parameter_2_11 ? phv_data_8 : _GEN_889; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_891 = 14'h9 == parameter_2_11 ? phv_data_9 : _GEN_890; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_892 = 14'ha == parameter_2_11 ? phv_data_10 : _GEN_891; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_893 = 14'hb == parameter_2_11 ? phv_data_11 : _GEN_892; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_894 = 14'hc == parameter_2_11 ? phv_data_12 : _GEN_893; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_895 = 14'hd == parameter_2_11 ? phv_data_13 : _GEN_894; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_896 = 14'he == parameter_2_11 ? phv_data_14 : _GEN_895; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_897 = 14'hf == parameter_2_11 ? phv_data_15 : _GEN_896; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_898 = 14'h10 == parameter_2_11 ? phv_data_16 : _GEN_897; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_899 = 14'h11 == parameter_2_11 ? phv_data_17 : _GEN_898; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_900 = 14'h12 == parameter_2_11 ? phv_data_18 : _GEN_899; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_901 = 14'h13 == parameter_2_11 ? phv_data_19 : _GEN_900; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_902 = 14'h14 == parameter_2_11 ? phv_data_20 : _GEN_901; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_903 = 14'h15 == parameter_2_11 ? phv_data_21 : _GEN_902; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_904 = 14'h16 == parameter_2_11 ? phv_data_22 : _GEN_903; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_905 = 14'h17 == parameter_2_11 ? phv_data_23 : _GEN_904; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_906 = 14'h18 == parameter_2_11 ? phv_data_24 : _GEN_905; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_907 = 14'h19 == parameter_2_11 ? phv_data_25 : _GEN_906; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_908 = 14'h1a == parameter_2_11 ? phv_data_26 : _GEN_907; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_909 = 14'h1b == parameter_2_11 ? phv_data_27 : _GEN_908; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_910 = 14'h1c == parameter_2_11 ? phv_data_28 : _GEN_909; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_911 = 14'h1d == parameter_2_11 ? phv_data_29 : _GEN_910; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_912 = 14'h1e == parameter_2_11 ? phv_data_30 : _GEN_911; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_913 = 14'h1f == parameter_2_11 ? phv_data_31 : _GEN_912; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_914 = 14'h20 == parameter_2_11 ? phv_data_32 : _GEN_913; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_915 = 14'h21 == parameter_2_11 ? phv_data_33 : _GEN_914; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_916 = 14'h22 == parameter_2_11 ? phv_data_34 : _GEN_915; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_917 = 14'h23 == parameter_2_11 ? phv_data_35 : _GEN_916; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_918 = 14'h24 == parameter_2_11 ? phv_data_36 : _GEN_917; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_919 = 14'h25 == parameter_2_11 ? phv_data_37 : _GEN_918; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_920 = 14'h26 == parameter_2_11 ? phv_data_38 : _GEN_919; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_921 = 14'h27 == parameter_2_11 ? phv_data_39 : _GEN_920; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_922 = 14'h28 == parameter_2_11 ? phv_data_40 : _GEN_921; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_923 = 14'h29 == parameter_2_11 ? phv_data_41 : _GEN_922; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_924 = 14'h2a == parameter_2_11 ? phv_data_42 : _GEN_923; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_925 = 14'h2b == parameter_2_11 ? phv_data_43 : _GEN_924; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_926 = 14'h2c == parameter_2_11 ? phv_data_44 : _GEN_925; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_927 = 14'h2d == parameter_2_11 ? phv_data_45 : _GEN_926; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_928 = 14'h2e == parameter_2_11 ? phv_data_46 : _GEN_927; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_929 = 14'h2f == parameter_2_11 ? phv_data_47 : _GEN_928; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_930 = 14'h30 == parameter_2_11 ? phv_data_48 : _GEN_929; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_931 = 14'h31 == parameter_2_11 ? phv_data_49 : _GEN_930; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_932 = 14'h32 == parameter_2_11 ? phv_data_50 : _GEN_931; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_933 = 14'h33 == parameter_2_11 ? phv_data_51 : _GEN_932; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_934 = 14'h34 == parameter_2_11 ? phv_data_52 : _GEN_933; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_935 = 14'h35 == parameter_2_11 ? phv_data_53 : _GEN_934; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_936 = 14'h36 == parameter_2_11 ? phv_data_54 : _GEN_935; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_937 = 14'h37 == parameter_2_11 ? phv_data_55 : _GEN_936; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_938 = 14'h38 == parameter_2_11 ? phv_data_56 : _GEN_937; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_939 = 14'h39 == parameter_2_11 ? phv_data_57 : _GEN_938; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_940 = 14'h3a == parameter_2_11 ? phv_data_58 : _GEN_939; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_941 = 14'h3b == parameter_2_11 ? phv_data_59 : _GEN_940; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_942 = 14'h3c == parameter_2_11 ? phv_data_60 : _GEN_941; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_943 = 14'h3d == parameter_2_11 ? phv_data_61 : _GEN_942; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_944 = 14'h3e == parameter_2_11 ? phv_data_62 : _GEN_943; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_945 = 14'h3f == parameter_2_11 ? phv_data_63 : _GEN_944; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_12 = vliw_12[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_12 = vliw_12[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_12 = parameter_2_12[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_12 = parameter_2_12[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_12 = {{1'd0}, args_offset_12}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_12 = _total_offset_T_12[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_949 = 3'h1 == total_offset_12 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_950 = 3'h2 == total_offset_12 ? args_2 : _GEN_949; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_951 = 3'h3 == total_offset_12 ? args_3 : _GEN_950; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_952 = 3'h4 == total_offset_12 ? args_4 : _GEN_951; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_953 = 3'h5 == total_offset_12 ? args_5 : _GEN_952; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_954 = 3'h6 == total_offset_12 ? args_6 : _GEN_953; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_955 = total_offset_12 < 3'h7 ? _GEN_954 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_12_0 = 3'h0 < args_length_12 ? _GEN_955 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_957 = opcode_12 == 4'ha ? field_bytes_12_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_958 = opcode_12 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_855 = opcode_12 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_25 = _T_855 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_959 = opcode_12 == 4'h8 | opcode_12 == 4'hb ? parameter_2_12[7:0] : _GEN_957; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_960 = opcode_12 == 4'h8 | opcode_12 == 4'hb ? _field_tag_T_25 : _GEN_958; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_961 = 14'h0 == parameter_2_12 ? phv_data_0 : _GEN_959; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_962 = 14'h1 == parameter_2_12 ? phv_data_1 : _GEN_961; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_963 = 14'h2 == parameter_2_12 ? phv_data_2 : _GEN_962; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_964 = 14'h3 == parameter_2_12 ? phv_data_3 : _GEN_963; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_965 = 14'h4 == parameter_2_12 ? phv_data_4 : _GEN_964; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_966 = 14'h5 == parameter_2_12 ? phv_data_5 : _GEN_965; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_967 = 14'h6 == parameter_2_12 ? phv_data_6 : _GEN_966; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_968 = 14'h7 == parameter_2_12 ? phv_data_7 : _GEN_967; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_969 = 14'h8 == parameter_2_12 ? phv_data_8 : _GEN_968; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_970 = 14'h9 == parameter_2_12 ? phv_data_9 : _GEN_969; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_971 = 14'ha == parameter_2_12 ? phv_data_10 : _GEN_970; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_972 = 14'hb == parameter_2_12 ? phv_data_11 : _GEN_971; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_973 = 14'hc == parameter_2_12 ? phv_data_12 : _GEN_972; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_974 = 14'hd == parameter_2_12 ? phv_data_13 : _GEN_973; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_975 = 14'he == parameter_2_12 ? phv_data_14 : _GEN_974; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_976 = 14'hf == parameter_2_12 ? phv_data_15 : _GEN_975; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_977 = 14'h10 == parameter_2_12 ? phv_data_16 : _GEN_976; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_978 = 14'h11 == parameter_2_12 ? phv_data_17 : _GEN_977; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_979 = 14'h12 == parameter_2_12 ? phv_data_18 : _GEN_978; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_980 = 14'h13 == parameter_2_12 ? phv_data_19 : _GEN_979; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_981 = 14'h14 == parameter_2_12 ? phv_data_20 : _GEN_980; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_982 = 14'h15 == parameter_2_12 ? phv_data_21 : _GEN_981; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_983 = 14'h16 == parameter_2_12 ? phv_data_22 : _GEN_982; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_984 = 14'h17 == parameter_2_12 ? phv_data_23 : _GEN_983; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_985 = 14'h18 == parameter_2_12 ? phv_data_24 : _GEN_984; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_986 = 14'h19 == parameter_2_12 ? phv_data_25 : _GEN_985; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_987 = 14'h1a == parameter_2_12 ? phv_data_26 : _GEN_986; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_988 = 14'h1b == parameter_2_12 ? phv_data_27 : _GEN_987; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_989 = 14'h1c == parameter_2_12 ? phv_data_28 : _GEN_988; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_990 = 14'h1d == parameter_2_12 ? phv_data_29 : _GEN_989; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_991 = 14'h1e == parameter_2_12 ? phv_data_30 : _GEN_990; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_992 = 14'h1f == parameter_2_12 ? phv_data_31 : _GEN_991; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_993 = 14'h20 == parameter_2_12 ? phv_data_32 : _GEN_992; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_994 = 14'h21 == parameter_2_12 ? phv_data_33 : _GEN_993; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_995 = 14'h22 == parameter_2_12 ? phv_data_34 : _GEN_994; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_996 = 14'h23 == parameter_2_12 ? phv_data_35 : _GEN_995; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_997 = 14'h24 == parameter_2_12 ? phv_data_36 : _GEN_996; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_998 = 14'h25 == parameter_2_12 ? phv_data_37 : _GEN_997; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_999 = 14'h26 == parameter_2_12 ? phv_data_38 : _GEN_998; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1000 = 14'h27 == parameter_2_12 ? phv_data_39 : _GEN_999; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1001 = 14'h28 == parameter_2_12 ? phv_data_40 : _GEN_1000; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1002 = 14'h29 == parameter_2_12 ? phv_data_41 : _GEN_1001; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1003 = 14'h2a == parameter_2_12 ? phv_data_42 : _GEN_1002; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1004 = 14'h2b == parameter_2_12 ? phv_data_43 : _GEN_1003; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1005 = 14'h2c == parameter_2_12 ? phv_data_44 : _GEN_1004; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1006 = 14'h2d == parameter_2_12 ? phv_data_45 : _GEN_1005; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1007 = 14'h2e == parameter_2_12 ? phv_data_46 : _GEN_1006; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1008 = 14'h2f == parameter_2_12 ? phv_data_47 : _GEN_1007; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1009 = 14'h30 == parameter_2_12 ? phv_data_48 : _GEN_1008; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1010 = 14'h31 == parameter_2_12 ? phv_data_49 : _GEN_1009; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1011 = 14'h32 == parameter_2_12 ? phv_data_50 : _GEN_1010; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1012 = 14'h33 == parameter_2_12 ? phv_data_51 : _GEN_1011; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1013 = 14'h34 == parameter_2_12 ? phv_data_52 : _GEN_1012; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1014 = 14'h35 == parameter_2_12 ? phv_data_53 : _GEN_1013; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1015 = 14'h36 == parameter_2_12 ? phv_data_54 : _GEN_1014; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1016 = 14'h37 == parameter_2_12 ? phv_data_55 : _GEN_1015; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1017 = 14'h38 == parameter_2_12 ? phv_data_56 : _GEN_1016; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1018 = 14'h39 == parameter_2_12 ? phv_data_57 : _GEN_1017; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1019 = 14'h3a == parameter_2_12 ? phv_data_58 : _GEN_1018; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1020 = 14'h3b == parameter_2_12 ? phv_data_59 : _GEN_1019; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1021 = 14'h3c == parameter_2_12 ? phv_data_60 : _GEN_1020; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1022 = 14'h3d == parameter_2_12 ? phv_data_61 : _GEN_1021; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1023 = 14'h3e == parameter_2_12 ? phv_data_62 : _GEN_1022; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1024 = 14'h3f == parameter_2_12 ? phv_data_63 : _GEN_1023; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_13 = vliw_13[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_13 = vliw_13[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_13 = parameter_2_13[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_13 = parameter_2_13[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_13 = {{1'd0}, args_offset_13}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_13 = _total_offset_T_13[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1028 = 3'h1 == total_offset_13 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1029 = 3'h2 == total_offset_13 ? args_2 : _GEN_1028; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1030 = 3'h3 == total_offset_13 ? args_3 : _GEN_1029; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1031 = 3'h4 == total_offset_13 ? args_4 : _GEN_1030; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1032 = 3'h5 == total_offset_13 ? args_5 : _GEN_1031; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1033 = 3'h6 == total_offset_13 ? args_6 : _GEN_1032; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1034 = total_offset_13 < 3'h7 ? _GEN_1033 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_13_0 = 3'h0 < args_length_13 ? _GEN_1034 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_1036 = opcode_13 == 4'ha ? field_bytes_13_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1037 = opcode_13 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_926 = opcode_13 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_27 = _T_926 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_1038 = opcode_13 == 4'h8 | opcode_13 == 4'hb ? parameter_2_13[7:0] : _GEN_1036; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_1039 = opcode_13 == 4'h8 | opcode_13 == 4'hb ? _field_tag_T_27 : _GEN_1037; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_1040 = 14'h0 == parameter_2_13 ? phv_data_0 : _GEN_1038; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1041 = 14'h1 == parameter_2_13 ? phv_data_1 : _GEN_1040; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1042 = 14'h2 == parameter_2_13 ? phv_data_2 : _GEN_1041; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1043 = 14'h3 == parameter_2_13 ? phv_data_3 : _GEN_1042; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1044 = 14'h4 == parameter_2_13 ? phv_data_4 : _GEN_1043; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1045 = 14'h5 == parameter_2_13 ? phv_data_5 : _GEN_1044; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1046 = 14'h6 == parameter_2_13 ? phv_data_6 : _GEN_1045; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1047 = 14'h7 == parameter_2_13 ? phv_data_7 : _GEN_1046; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1048 = 14'h8 == parameter_2_13 ? phv_data_8 : _GEN_1047; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1049 = 14'h9 == parameter_2_13 ? phv_data_9 : _GEN_1048; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1050 = 14'ha == parameter_2_13 ? phv_data_10 : _GEN_1049; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1051 = 14'hb == parameter_2_13 ? phv_data_11 : _GEN_1050; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1052 = 14'hc == parameter_2_13 ? phv_data_12 : _GEN_1051; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1053 = 14'hd == parameter_2_13 ? phv_data_13 : _GEN_1052; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1054 = 14'he == parameter_2_13 ? phv_data_14 : _GEN_1053; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1055 = 14'hf == parameter_2_13 ? phv_data_15 : _GEN_1054; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1056 = 14'h10 == parameter_2_13 ? phv_data_16 : _GEN_1055; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1057 = 14'h11 == parameter_2_13 ? phv_data_17 : _GEN_1056; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1058 = 14'h12 == parameter_2_13 ? phv_data_18 : _GEN_1057; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1059 = 14'h13 == parameter_2_13 ? phv_data_19 : _GEN_1058; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1060 = 14'h14 == parameter_2_13 ? phv_data_20 : _GEN_1059; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1061 = 14'h15 == parameter_2_13 ? phv_data_21 : _GEN_1060; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1062 = 14'h16 == parameter_2_13 ? phv_data_22 : _GEN_1061; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1063 = 14'h17 == parameter_2_13 ? phv_data_23 : _GEN_1062; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1064 = 14'h18 == parameter_2_13 ? phv_data_24 : _GEN_1063; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1065 = 14'h19 == parameter_2_13 ? phv_data_25 : _GEN_1064; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1066 = 14'h1a == parameter_2_13 ? phv_data_26 : _GEN_1065; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1067 = 14'h1b == parameter_2_13 ? phv_data_27 : _GEN_1066; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1068 = 14'h1c == parameter_2_13 ? phv_data_28 : _GEN_1067; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1069 = 14'h1d == parameter_2_13 ? phv_data_29 : _GEN_1068; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1070 = 14'h1e == parameter_2_13 ? phv_data_30 : _GEN_1069; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1071 = 14'h1f == parameter_2_13 ? phv_data_31 : _GEN_1070; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1072 = 14'h20 == parameter_2_13 ? phv_data_32 : _GEN_1071; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1073 = 14'h21 == parameter_2_13 ? phv_data_33 : _GEN_1072; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1074 = 14'h22 == parameter_2_13 ? phv_data_34 : _GEN_1073; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1075 = 14'h23 == parameter_2_13 ? phv_data_35 : _GEN_1074; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1076 = 14'h24 == parameter_2_13 ? phv_data_36 : _GEN_1075; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1077 = 14'h25 == parameter_2_13 ? phv_data_37 : _GEN_1076; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1078 = 14'h26 == parameter_2_13 ? phv_data_38 : _GEN_1077; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1079 = 14'h27 == parameter_2_13 ? phv_data_39 : _GEN_1078; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1080 = 14'h28 == parameter_2_13 ? phv_data_40 : _GEN_1079; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1081 = 14'h29 == parameter_2_13 ? phv_data_41 : _GEN_1080; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1082 = 14'h2a == parameter_2_13 ? phv_data_42 : _GEN_1081; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1083 = 14'h2b == parameter_2_13 ? phv_data_43 : _GEN_1082; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1084 = 14'h2c == parameter_2_13 ? phv_data_44 : _GEN_1083; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1085 = 14'h2d == parameter_2_13 ? phv_data_45 : _GEN_1084; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1086 = 14'h2e == parameter_2_13 ? phv_data_46 : _GEN_1085; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1087 = 14'h2f == parameter_2_13 ? phv_data_47 : _GEN_1086; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1088 = 14'h30 == parameter_2_13 ? phv_data_48 : _GEN_1087; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1089 = 14'h31 == parameter_2_13 ? phv_data_49 : _GEN_1088; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1090 = 14'h32 == parameter_2_13 ? phv_data_50 : _GEN_1089; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1091 = 14'h33 == parameter_2_13 ? phv_data_51 : _GEN_1090; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1092 = 14'h34 == parameter_2_13 ? phv_data_52 : _GEN_1091; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1093 = 14'h35 == parameter_2_13 ? phv_data_53 : _GEN_1092; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1094 = 14'h36 == parameter_2_13 ? phv_data_54 : _GEN_1093; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1095 = 14'h37 == parameter_2_13 ? phv_data_55 : _GEN_1094; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1096 = 14'h38 == parameter_2_13 ? phv_data_56 : _GEN_1095; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1097 = 14'h39 == parameter_2_13 ? phv_data_57 : _GEN_1096; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1098 = 14'h3a == parameter_2_13 ? phv_data_58 : _GEN_1097; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1099 = 14'h3b == parameter_2_13 ? phv_data_59 : _GEN_1098; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1100 = 14'h3c == parameter_2_13 ? phv_data_60 : _GEN_1099; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1101 = 14'h3d == parameter_2_13 ? phv_data_61 : _GEN_1100; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1102 = 14'h3e == parameter_2_13 ? phv_data_62 : _GEN_1101; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1103 = 14'h3f == parameter_2_13 ? phv_data_63 : _GEN_1102; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_14 = vliw_14[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_14 = vliw_14[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_14 = parameter_2_14[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_14 = parameter_2_14[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_14 = {{1'd0}, args_offset_14}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_14 = _total_offset_T_14[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1107 = 3'h1 == total_offset_14 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1108 = 3'h2 == total_offset_14 ? args_2 : _GEN_1107; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1109 = 3'h3 == total_offset_14 ? args_3 : _GEN_1108; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1110 = 3'h4 == total_offset_14 ? args_4 : _GEN_1109; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1111 = 3'h5 == total_offset_14 ? args_5 : _GEN_1110; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1112 = 3'h6 == total_offset_14 ? args_6 : _GEN_1111; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1113 = total_offset_14 < 3'h7 ? _GEN_1112 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_14_0 = 3'h0 < args_length_14 ? _GEN_1113 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_1115 = opcode_14 == 4'ha ? field_bytes_14_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1116 = opcode_14 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_997 = opcode_14 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_29 = _T_997 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_1117 = opcode_14 == 4'h8 | opcode_14 == 4'hb ? parameter_2_14[7:0] : _GEN_1115; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_1118 = opcode_14 == 4'h8 | opcode_14 == 4'hb ? _field_tag_T_29 : _GEN_1116; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_1119 = 14'h0 == parameter_2_14 ? phv_data_0 : _GEN_1117; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1120 = 14'h1 == parameter_2_14 ? phv_data_1 : _GEN_1119; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1121 = 14'h2 == parameter_2_14 ? phv_data_2 : _GEN_1120; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1122 = 14'h3 == parameter_2_14 ? phv_data_3 : _GEN_1121; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1123 = 14'h4 == parameter_2_14 ? phv_data_4 : _GEN_1122; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1124 = 14'h5 == parameter_2_14 ? phv_data_5 : _GEN_1123; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1125 = 14'h6 == parameter_2_14 ? phv_data_6 : _GEN_1124; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1126 = 14'h7 == parameter_2_14 ? phv_data_7 : _GEN_1125; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1127 = 14'h8 == parameter_2_14 ? phv_data_8 : _GEN_1126; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1128 = 14'h9 == parameter_2_14 ? phv_data_9 : _GEN_1127; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1129 = 14'ha == parameter_2_14 ? phv_data_10 : _GEN_1128; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1130 = 14'hb == parameter_2_14 ? phv_data_11 : _GEN_1129; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1131 = 14'hc == parameter_2_14 ? phv_data_12 : _GEN_1130; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1132 = 14'hd == parameter_2_14 ? phv_data_13 : _GEN_1131; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1133 = 14'he == parameter_2_14 ? phv_data_14 : _GEN_1132; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1134 = 14'hf == parameter_2_14 ? phv_data_15 : _GEN_1133; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1135 = 14'h10 == parameter_2_14 ? phv_data_16 : _GEN_1134; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1136 = 14'h11 == parameter_2_14 ? phv_data_17 : _GEN_1135; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1137 = 14'h12 == parameter_2_14 ? phv_data_18 : _GEN_1136; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1138 = 14'h13 == parameter_2_14 ? phv_data_19 : _GEN_1137; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1139 = 14'h14 == parameter_2_14 ? phv_data_20 : _GEN_1138; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1140 = 14'h15 == parameter_2_14 ? phv_data_21 : _GEN_1139; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1141 = 14'h16 == parameter_2_14 ? phv_data_22 : _GEN_1140; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1142 = 14'h17 == parameter_2_14 ? phv_data_23 : _GEN_1141; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1143 = 14'h18 == parameter_2_14 ? phv_data_24 : _GEN_1142; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1144 = 14'h19 == parameter_2_14 ? phv_data_25 : _GEN_1143; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1145 = 14'h1a == parameter_2_14 ? phv_data_26 : _GEN_1144; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1146 = 14'h1b == parameter_2_14 ? phv_data_27 : _GEN_1145; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1147 = 14'h1c == parameter_2_14 ? phv_data_28 : _GEN_1146; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1148 = 14'h1d == parameter_2_14 ? phv_data_29 : _GEN_1147; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1149 = 14'h1e == parameter_2_14 ? phv_data_30 : _GEN_1148; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1150 = 14'h1f == parameter_2_14 ? phv_data_31 : _GEN_1149; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1151 = 14'h20 == parameter_2_14 ? phv_data_32 : _GEN_1150; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1152 = 14'h21 == parameter_2_14 ? phv_data_33 : _GEN_1151; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1153 = 14'h22 == parameter_2_14 ? phv_data_34 : _GEN_1152; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1154 = 14'h23 == parameter_2_14 ? phv_data_35 : _GEN_1153; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1155 = 14'h24 == parameter_2_14 ? phv_data_36 : _GEN_1154; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1156 = 14'h25 == parameter_2_14 ? phv_data_37 : _GEN_1155; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1157 = 14'h26 == parameter_2_14 ? phv_data_38 : _GEN_1156; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1158 = 14'h27 == parameter_2_14 ? phv_data_39 : _GEN_1157; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1159 = 14'h28 == parameter_2_14 ? phv_data_40 : _GEN_1158; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1160 = 14'h29 == parameter_2_14 ? phv_data_41 : _GEN_1159; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1161 = 14'h2a == parameter_2_14 ? phv_data_42 : _GEN_1160; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1162 = 14'h2b == parameter_2_14 ? phv_data_43 : _GEN_1161; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1163 = 14'h2c == parameter_2_14 ? phv_data_44 : _GEN_1162; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1164 = 14'h2d == parameter_2_14 ? phv_data_45 : _GEN_1163; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1165 = 14'h2e == parameter_2_14 ? phv_data_46 : _GEN_1164; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1166 = 14'h2f == parameter_2_14 ? phv_data_47 : _GEN_1165; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1167 = 14'h30 == parameter_2_14 ? phv_data_48 : _GEN_1166; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1168 = 14'h31 == parameter_2_14 ? phv_data_49 : _GEN_1167; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1169 = 14'h32 == parameter_2_14 ? phv_data_50 : _GEN_1168; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1170 = 14'h33 == parameter_2_14 ? phv_data_51 : _GEN_1169; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1171 = 14'h34 == parameter_2_14 ? phv_data_52 : _GEN_1170; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1172 = 14'h35 == parameter_2_14 ? phv_data_53 : _GEN_1171; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1173 = 14'h36 == parameter_2_14 ? phv_data_54 : _GEN_1172; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1174 = 14'h37 == parameter_2_14 ? phv_data_55 : _GEN_1173; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1175 = 14'h38 == parameter_2_14 ? phv_data_56 : _GEN_1174; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1176 = 14'h39 == parameter_2_14 ? phv_data_57 : _GEN_1175; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1177 = 14'h3a == parameter_2_14 ? phv_data_58 : _GEN_1176; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1178 = 14'h3b == parameter_2_14 ? phv_data_59 : _GEN_1177; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1179 = 14'h3c == parameter_2_14 ? phv_data_60 : _GEN_1178; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1180 = 14'h3d == parameter_2_14 ? phv_data_61 : _GEN_1179; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1181 = 14'h3e == parameter_2_14 ? phv_data_62 : _GEN_1180; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1182 = 14'h3f == parameter_2_14 ? phv_data_63 : _GEN_1181; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_15 = vliw_15[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_15 = vliw_15[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_15 = parameter_2_15[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_15 = parameter_2_15[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_15 = {{1'd0}, args_offset_15}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_15 = _total_offset_T_15[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1186 = 3'h1 == total_offset_15 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1187 = 3'h2 == total_offset_15 ? args_2 : _GEN_1186; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1188 = 3'h3 == total_offset_15 ? args_3 : _GEN_1187; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1189 = 3'h4 == total_offset_15 ? args_4 : _GEN_1188; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1190 = 3'h5 == total_offset_15 ? args_5 : _GEN_1189; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1191 = 3'h6 == total_offset_15 ? args_6 : _GEN_1190; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1192 = total_offset_15 < 3'h7 ? _GEN_1191 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_15_0 = 3'h0 < args_length_15 ? _GEN_1192 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_1194 = opcode_15 == 4'ha ? field_bytes_15_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1195 = opcode_15 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1068 = opcode_15 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_31 = _T_1068 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_1196 = opcode_15 == 4'h8 | opcode_15 == 4'hb ? parameter_2_15[7:0] : _GEN_1194; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_1197 = opcode_15 == 4'h8 | opcode_15 == 4'hb ? _field_tag_T_31 : _GEN_1195; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_1198 = 14'h0 == parameter_2_15 ? phv_data_0 : _GEN_1196; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1199 = 14'h1 == parameter_2_15 ? phv_data_1 : _GEN_1198; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1200 = 14'h2 == parameter_2_15 ? phv_data_2 : _GEN_1199; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1201 = 14'h3 == parameter_2_15 ? phv_data_3 : _GEN_1200; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1202 = 14'h4 == parameter_2_15 ? phv_data_4 : _GEN_1201; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1203 = 14'h5 == parameter_2_15 ? phv_data_5 : _GEN_1202; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1204 = 14'h6 == parameter_2_15 ? phv_data_6 : _GEN_1203; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1205 = 14'h7 == parameter_2_15 ? phv_data_7 : _GEN_1204; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1206 = 14'h8 == parameter_2_15 ? phv_data_8 : _GEN_1205; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1207 = 14'h9 == parameter_2_15 ? phv_data_9 : _GEN_1206; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1208 = 14'ha == parameter_2_15 ? phv_data_10 : _GEN_1207; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1209 = 14'hb == parameter_2_15 ? phv_data_11 : _GEN_1208; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1210 = 14'hc == parameter_2_15 ? phv_data_12 : _GEN_1209; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1211 = 14'hd == parameter_2_15 ? phv_data_13 : _GEN_1210; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1212 = 14'he == parameter_2_15 ? phv_data_14 : _GEN_1211; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1213 = 14'hf == parameter_2_15 ? phv_data_15 : _GEN_1212; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1214 = 14'h10 == parameter_2_15 ? phv_data_16 : _GEN_1213; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1215 = 14'h11 == parameter_2_15 ? phv_data_17 : _GEN_1214; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1216 = 14'h12 == parameter_2_15 ? phv_data_18 : _GEN_1215; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1217 = 14'h13 == parameter_2_15 ? phv_data_19 : _GEN_1216; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1218 = 14'h14 == parameter_2_15 ? phv_data_20 : _GEN_1217; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1219 = 14'h15 == parameter_2_15 ? phv_data_21 : _GEN_1218; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1220 = 14'h16 == parameter_2_15 ? phv_data_22 : _GEN_1219; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1221 = 14'h17 == parameter_2_15 ? phv_data_23 : _GEN_1220; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1222 = 14'h18 == parameter_2_15 ? phv_data_24 : _GEN_1221; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1223 = 14'h19 == parameter_2_15 ? phv_data_25 : _GEN_1222; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1224 = 14'h1a == parameter_2_15 ? phv_data_26 : _GEN_1223; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1225 = 14'h1b == parameter_2_15 ? phv_data_27 : _GEN_1224; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1226 = 14'h1c == parameter_2_15 ? phv_data_28 : _GEN_1225; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1227 = 14'h1d == parameter_2_15 ? phv_data_29 : _GEN_1226; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1228 = 14'h1e == parameter_2_15 ? phv_data_30 : _GEN_1227; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1229 = 14'h1f == parameter_2_15 ? phv_data_31 : _GEN_1228; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1230 = 14'h20 == parameter_2_15 ? phv_data_32 : _GEN_1229; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1231 = 14'h21 == parameter_2_15 ? phv_data_33 : _GEN_1230; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1232 = 14'h22 == parameter_2_15 ? phv_data_34 : _GEN_1231; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1233 = 14'h23 == parameter_2_15 ? phv_data_35 : _GEN_1232; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1234 = 14'h24 == parameter_2_15 ? phv_data_36 : _GEN_1233; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1235 = 14'h25 == parameter_2_15 ? phv_data_37 : _GEN_1234; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1236 = 14'h26 == parameter_2_15 ? phv_data_38 : _GEN_1235; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1237 = 14'h27 == parameter_2_15 ? phv_data_39 : _GEN_1236; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1238 = 14'h28 == parameter_2_15 ? phv_data_40 : _GEN_1237; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1239 = 14'h29 == parameter_2_15 ? phv_data_41 : _GEN_1238; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1240 = 14'h2a == parameter_2_15 ? phv_data_42 : _GEN_1239; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1241 = 14'h2b == parameter_2_15 ? phv_data_43 : _GEN_1240; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1242 = 14'h2c == parameter_2_15 ? phv_data_44 : _GEN_1241; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1243 = 14'h2d == parameter_2_15 ? phv_data_45 : _GEN_1242; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1244 = 14'h2e == parameter_2_15 ? phv_data_46 : _GEN_1243; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1245 = 14'h2f == parameter_2_15 ? phv_data_47 : _GEN_1244; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1246 = 14'h30 == parameter_2_15 ? phv_data_48 : _GEN_1245; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1247 = 14'h31 == parameter_2_15 ? phv_data_49 : _GEN_1246; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1248 = 14'h32 == parameter_2_15 ? phv_data_50 : _GEN_1247; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1249 = 14'h33 == parameter_2_15 ? phv_data_51 : _GEN_1248; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1250 = 14'h34 == parameter_2_15 ? phv_data_52 : _GEN_1249; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1251 = 14'h35 == parameter_2_15 ? phv_data_53 : _GEN_1250; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1252 = 14'h36 == parameter_2_15 ? phv_data_54 : _GEN_1251; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1253 = 14'h37 == parameter_2_15 ? phv_data_55 : _GEN_1252; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1254 = 14'h38 == parameter_2_15 ? phv_data_56 : _GEN_1253; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1255 = 14'h39 == parameter_2_15 ? phv_data_57 : _GEN_1254; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1256 = 14'h3a == parameter_2_15 ? phv_data_58 : _GEN_1255; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1257 = 14'h3b == parameter_2_15 ? phv_data_59 : _GEN_1256; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1258 = 14'h3c == parameter_2_15 ? phv_data_60 : _GEN_1257; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1259 = 14'h3d == parameter_2_15 ? phv_data_61 : _GEN_1258; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1260 = 14'h3e == parameter_2_15 ? phv_data_62 : _GEN_1259; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1261 = 14'h3f == parameter_2_15 ? phv_data_63 : _GEN_1260; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_16 = vliw_16[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_16 = vliw_16[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_16 = parameter_2_16[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_16 = parameter_2_16[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_16 = {{1'd0}, args_offset_16}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_16 = _total_offset_T_16[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1265 = 3'h1 == total_offset_16 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1266 = 3'h2 == total_offset_16 ? args_2 : _GEN_1265; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1267 = 3'h3 == total_offset_16 ? args_3 : _GEN_1266; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1268 = 3'h4 == total_offset_16 ? args_4 : _GEN_1267; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1269 = 3'h5 == total_offset_16 ? args_5 : _GEN_1268; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1270 = 3'h6 == total_offset_16 ? args_6 : _GEN_1269; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1271 = total_offset_16 < 3'h7 ? _GEN_1270 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_16_0 = 3'h0 < args_length_16 ? _GEN_1271 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_1273 = opcode_16 == 4'ha ? field_bytes_16_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1274 = opcode_16 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1139 = opcode_16 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_33 = _T_1139 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_1275 = opcode_16 == 4'h8 | opcode_16 == 4'hb ? parameter_2_16[7:0] : _GEN_1273; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_1276 = opcode_16 == 4'h8 | opcode_16 == 4'hb ? _field_tag_T_33 : _GEN_1274; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_1277 = 14'h0 == parameter_2_16 ? phv_data_0 : _GEN_1275; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1278 = 14'h1 == parameter_2_16 ? phv_data_1 : _GEN_1277; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1279 = 14'h2 == parameter_2_16 ? phv_data_2 : _GEN_1278; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1280 = 14'h3 == parameter_2_16 ? phv_data_3 : _GEN_1279; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1281 = 14'h4 == parameter_2_16 ? phv_data_4 : _GEN_1280; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1282 = 14'h5 == parameter_2_16 ? phv_data_5 : _GEN_1281; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1283 = 14'h6 == parameter_2_16 ? phv_data_6 : _GEN_1282; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1284 = 14'h7 == parameter_2_16 ? phv_data_7 : _GEN_1283; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1285 = 14'h8 == parameter_2_16 ? phv_data_8 : _GEN_1284; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1286 = 14'h9 == parameter_2_16 ? phv_data_9 : _GEN_1285; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1287 = 14'ha == parameter_2_16 ? phv_data_10 : _GEN_1286; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1288 = 14'hb == parameter_2_16 ? phv_data_11 : _GEN_1287; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1289 = 14'hc == parameter_2_16 ? phv_data_12 : _GEN_1288; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1290 = 14'hd == parameter_2_16 ? phv_data_13 : _GEN_1289; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1291 = 14'he == parameter_2_16 ? phv_data_14 : _GEN_1290; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1292 = 14'hf == parameter_2_16 ? phv_data_15 : _GEN_1291; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1293 = 14'h10 == parameter_2_16 ? phv_data_16 : _GEN_1292; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1294 = 14'h11 == parameter_2_16 ? phv_data_17 : _GEN_1293; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1295 = 14'h12 == parameter_2_16 ? phv_data_18 : _GEN_1294; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1296 = 14'h13 == parameter_2_16 ? phv_data_19 : _GEN_1295; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1297 = 14'h14 == parameter_2_16 ? phv_data_20 : _GEN_1296; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1298 = 14'h15 == parameter_2_16 ? phv_data_21 : _GEN_1297; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1299 = 14'h16 == parameter_2_16 ? phv_data_22 : _GEN_1298; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1300 = 14'h17 == parameter_2_16 ? phv_data_23 : _GEN_1299; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1301 = 14'h18 == parameter_2_16 ? phv_data_24 : _GEN_1300; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1302 = 14'h19 == parameter_2_16 ? phv_data_25 : _GEN_1301; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1303 = 14'h1a == parameter_2_16 ? phv_data_26 : _GEN_1302; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1304 = 14'h1b == parameter_2_16 ? phv_data_27 : _GEN_1303; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1305 = 14'h1c == parameter_2_16 ? phv_data_28 : _GEN_1304; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1306 = 14'h1d == parameter_2_16 ? phv_data_29 : _GEN_1305; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1307 = 14'h1e == parameter_2_16 ? phv_data_30 : _GEN_1306; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1308 = 14'h1f == parameter_2_16 ? phv_data_31 : _GEN_1307; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1309 = 14'h20 == parameter_2_16 ? phv_data_32 : _GEN_1308; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1310 = 14'h21 == parameter_2_16 ? phv_data_33 : _GEN_1309; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1311 = 14'h22 == parameter_2_16 ? phv_data_34 : _GEN_1310; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1312 = 14'h23 == parameter_2_16 ? phv_data_35 : _GEN_1311; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1313 = 14'h24 == parameter_2_16 ? phv_data_36 : _GEN_1312; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1314 = 14'h25 == parameter_2_16 ? phv_data_37 : _GEN_1313; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1315 = 14'h26 == parameter_2_16 ? phv_data_38 : _GEN_1314; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1316 = 14'h27 == parameter_2_16 ? phv_data_39 : _GEN_1315; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1317 = 14'h28 == parameter_2_16 ? phv_data_40 : _GEN_1316; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1318 = 14'h29 == parameter_2_16 ? phv_data_41 : _GEN_1317; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1319 = 14'h2a == parameter_2_16 ? phv_data_42 : _GEN_1318; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1320 = 14'h2b == parameter_2_16 ? phv_data_43 : _GEN_1319; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1321 = 14'h2c == parameter_2_16 ? phv_data_44 : _GEN_1320; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1322 = 14'h2d == parameter_2_16 ? phv_data_45 : _GEN_1321; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1323 = 14'h2e == parameter_2_16 ? phv_data_46 : _GEN_1322; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1324 = 14'h2f == parameter_2_16 ? phv_data_47 : _GEN_1323; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1325 = 14'h30 == parameter_2_16 ? phv_data_48 : _GEN_1324; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1326 = 14'h31 == parameter_2_16 ? phv_data_49 : _GEN_1325; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1327 = 14'h32 == parameter_2_16 ? phv_data_50 : _GEN_1326; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1328 = 14'h33 == parameter_2_16 ? phv_data_51 : _GEN_1327; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1329 = 14'h34 == parameter_2_16 ? phv_data_52 : _GEN_1328; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1330 = 14'h35 == parameter_2_16 ? phv_data_53 : _GEN_1329; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1331 = 14'h36 == parameter_2_16 ? phv_data_54 : _GEN_1330; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1332 = 14'h37 == parameter_2_16 ? phv_data_55 : _GEN_1331; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1333 = 14'h38 == parameter_2_16 ? phv_data_56 : _GEN_1332; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1334 = 14'h39 == parameter_2_16 ? phv_data_57 : _GEN_1333; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1335 = 14'h3a == parameter_2_16 ? phv_data_58 : _GEN_1334; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1336 = 14'h3b == parameter_2_16 ? phv_data_59 : _GEN_1335; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1337 = 14'h3c == parameter_2_16 ? phv_data_60 : _GEN_1336; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1338 = 14'h3d == parameter_2_16 ? phv_data_61 : _GEN_1337; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1339 = 14'h3e == parameter_2_16 ? phv_data_62 : _GEN_1338; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1340 = 14'h3f == parameter_2_16 ? phv_data_63 : _GEN_1339; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_17 = vliw_17[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_17 = vliw_17[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_17 = parameter_2_17[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_17 = parameter_2_17[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_17 = {{1'd0}, args_offset_17}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_17 = _total_offset_T_17[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1344 = 3'h1 == total_offset_17 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1345 = 3'h2 == total_offset_17 ? args_2 : _GEN_1344; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1346 = 3'h3 == total_offset_17 ? args_3 : _GEN_1345; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1347 = 3'h4 == total_offset_17 ? args_4 : _GEN_1346; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1348 = 3'h5 == total_offset_17 ? args_5 : _GEN_1347; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1349 = 3'h6 == total_offset_17 ? args_6 : _GEN_1348; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1350 = total_offset_17 < 3'h7 ? _GEN_1349 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_17_0 = 3'h0 < args_length_17 ? _GEN_1350 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_1352 = opcode_17 == 4'ha ? field_bytes_17_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1353 = opcode_17 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1210 = opcode_17 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_35 = _T_1210 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_1354 = opcode_17 == 4'h8 | opcode_17 == 4'hb ? parameter_2_17[7:0] : _GEN_1352; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_1355 = opcode_17 == 4'h8 | opcode_17 == 4'hb ? _field_tag_T_35 : _GEN_1353; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_1356 = 14'h0 == parameter_2_17 ? phv_data_0 : _GEN_1354; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1357 = 14'h1 == parameter_2_17 ? phv_data_1 : _GEN_1356; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1358 = 14'h2 == parameter_2_17 ? phv_data_2 : _GEN_1357; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1359 = 14'h3 == parameter_2_17 ? phv_data_3 : _GEN_1358; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1360 = 14'h4 == parameter_2_17 ? phv_data_4 : _GEN_1359; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1361 = 14'h5 == parameter_2_17 ? phv_data_5 : _GEN_1360; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1362 = 14'h6 == parameter_2_17 ? phv_data_6 : _GEN_1361; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1363 = 14'h7 == parameter_2_17 ? phv_data_7 : _GEN_1362; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1364 = 14'h8 == parameter_2_17 ? phv_data_8 : _GEN_1363; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1365 = 14'h9 == parameter_2_17 ? phv_data_9 : _GEN_1364; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1366 = 14'ha == parameter_2_17 ? phv_data_10 : _GEN_1365; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1367 = 14'hb == parameter_2_17 ? phv_data_11 : _GEN_1366; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1368 = 14'hc == parameter_2_17 ? phv_data_12 : _GEN_1367; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1369 = 14'hd == parameter_2_17 ? phv_data_13 : _GEN_1368; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1370 = 14'he == parameter_2_17 ? phv_data_14 : _GEN_1369; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1371 = 14'hf == parameter_2_17 ? phv_data_15 : _GEN_1370; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1372 = 14'h10 == parameter_2_17 ? phv_data_16 : _GEN_1371; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1373 = 14'h11 == parameter_2_17 ? phv_data_17 : _GEN_1372; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1374 = 14'h12 == parameter_2_17 ? phv_data_18 : _GEN_1373; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1375 = 14'h13 == parameter_2_17 ? phv_data_19 : _GEN_1374; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1376 = 14'h14 == parameter_2_17 ? phv_data_20 : _GEN_1375; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1377 = 14'h15 == parameter_2_17 ? phv_data_21 : _GEN_1376; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1378 = 14'h16 == parameter_2_17 ? phv_data_22 : _GEN_1377; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1379 = 14'h17 == parameter_2_17 ? phv_data_23 : _GEN_1378; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1380 = 14'h18 == parameter_2_17 ? phv_data_24 : _GEN_1379; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1381 = 14'h19 == parameter_2_17 ? phv_data_25 : _GEN_1380; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1382 = 14'h1a == parameter_2_17 ? phv_data_26 : _GEN_1381; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1383 = 14'h1b == parameter_2_17 ? phv_data_27 : _GEN_1382; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1384 = 14'h1c == parameter_2_17 ? phv_data_28 : _GEN_1383; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1385 = 14'h1d == parameter_2_17 ? phv_data_29 : _GEN_1384; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1386 = 14'h1e == parameter_2_17 ? phv_data_30 : _GEN_1385; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1387 = 14'h1f == parameter_2_17 ? phv_data_31 : _GEN_1386; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1388 = 14'h20 == parameter_2_17 ? phv_data_32 : _GEN_1387; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1389 = 14'h21 == parameter_2_17 ? phv_data_33 : _GEN_1388; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1390 = 14'h22 == parameter_2_17 ? phv_data_34 : _GEN_1389; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1391 = 14'h23 == parameter_2_17 ? phv_data_35 : _GEN_1390; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1392 = 14'h24 == parameter_2_17 ? phv_data_36 : _GEN_1391; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1393 = 14'h25 == parameter_2_17 ? phv_data_37 : _GEN_1392; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1394 = 14'h26 == parameter_2_17 ? phv_data_38 : _GEN_1393; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1395 = 14'h27 == parameter_2_17 ? phv_data_39 : _GEN_1394; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1396 = 14'h28 == parameter_2_17 ? phv_data_40 : _GEN_1395; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1397 = 14'h29 == parameter_2_17 ? phv_data_41 : _GEN_1396; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1398 = 14'h2a == parameter_2_17 ? phv_data_42 : _GEN_1397; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1399 = 14'h2b == parameter_2_17 ? phv_data_43 : _GEN_1398; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1400 = 14'h2c == parameter_2_17 ? phv_data_44 : _GEN_1399; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1401 = 14'h2d == parameter_2_17 ? phv_data_45 : _GEN_1400; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1402 = 14'h2e == parameter_2_17 ? phv_data_46 : _GEN_1401; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1403 = 14'h2f == parameter_2_17 ? phv_data_47 : _GEN_1402; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1404 = 14'h30 == parameter_2_17 ? phv_data_48 : _GEN_1403; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1405 = 14'h31 == parameter_2_17 ? phv_data_49 : _GEN_1404; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1406 = 14'h32 == parameter_2_17 ? phv_data_50 : _GEN_1405; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1407 = 14'h33 == parameter_2_17 ? phv_data_51 : _GEN_1406; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1408 = 14'h34 == parameter_2_17 ? phv_data_52 : _GEN_1407; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1409 = 14'h35 == parameter_2_17 ? phv_data_53 : _GEN_1408; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1410 = 14'h36 == parameter_2_17 ? phv_data_54 : _GEN_1409; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1411 = 14'h37 == parameter_2_17 ? phv_data_55 : _GEN_1410; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1412 = 14'h38 == parameter_2_17 ? phv_data_56 : _GEN_1411; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1413 = 14'h39 == parameter_2_17 ? phv_data_57 : _GEN_1412; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1414 = 14'h3a == parameter_2_17 ? phv_data_58 : _GEN_1413; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1415 = 14'h3b == parameter_2_17 ? phv_data_59 : _GEN_1414; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1416 = 14'h3c == parameter_2_17 ? phv_data_60 : _GEN_1415; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1417 = 14'h3d == parameter_2_17 ? phv_data_61 : _GEN_1416; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1418 = 14'h3e == parameter_2_17 ? phv_data_62 : _GEN_1417; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1419 = 14'h3f == parameter_2_17 ? phv_data_63 : _GEN_1418; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_18 = vliw_18[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_18 = vliw_18[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_18 = parameter_2_18[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_18 = parameter_2_18[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_18 = {{1'd0}, args_offset_18}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_18 = _total_offset_T_18[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1423 = 3'h1 == total_offset_18 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1424 = 3'h2 == total_offset_18 ? args_2 : _GEN_1423; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1425 = 3'h3 == total_offset_18 ? args_3 : _GEN_1424; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1426 = 3'h4 == total_offset_18 ? args_4 : _GEN_1425; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1427 = 3'h5 == total_offset_18 ? args_5 : _GEN_1426; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1428 = 3'h6 == total_offset_18 ? args_6 : _GEN_1427; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1429 = total_offset_18 < 3'h7 ? _GEN_1428 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_18_0 = 3'h0 < args_length_18 ? _GEN_1429 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_1431 = opcode_18 == 4'ha ? field_bytes_18_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1432 = opcode_18 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1281 = opcode_18 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_37 = _T_1281 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_1433 = opcode_18 == 4'h8 | opcode_18 == 4'hb ? parameter_2_18[7:0] : _GEN_1431; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_1434 = opcode_18 == 4'h8 | opcode_18 == 4'hb ? _field_tag_T_37 : _GEN_1432; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_1435 = 14'h0 == parameter_2_18 ? phv_data_0 : _GEN_1433; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1436 = 14'h1 == parameter_2_18 ? phv_data_1 : _GEN_1435; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1437 = 14'h2 == parameter_2_18 ? phv_data_2 : _GEN_1436; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1438 = 14'h3 == parameter_2_18 ? phv_data_3 : _GEN_1437; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1439 = 14'h4 == parameter_2_18 ? phv_data_4 : _GEN_1438; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1440 = 14'h5 == parameter_2_18 ? phv_data_5 : _GEN_1439; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1441 = 14'h6 == parameter_2_18 ? phv_data_6 : _GEN_1440; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1442 = 14'h7 == parameter_2_18 ? phv_data_7 : _GEN_1441; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1443 = 14'h8 == parameter_2_18 ? phv_data_8 : _GEN_1442; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1444 = 14'h9 == parameter_2_18 ? phv_data_9 : _GEN_1443; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1445 = 14'ha == parameter_2_18 ? phv_data_10 : _GEN_1444; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1446 = 14'hb == parameter_2_18 ? phv_data_11 : _GEN_1445; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1447 = 14'hc == parameter_2_18 ? phv_data_12 : _GEN_1446; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1448 = 14'hd == parameter_2_18 ? phv_data_13 : _GEN_1447; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1449 = 14'he == parameter_2_18 ? phv_data_14 : _GEN_1448; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1450 = 14'hf == parameter_2_18 ? phv_data_15 : _GEN_1449; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1451 = 14'h10 == parameter_2_18 ? phv_data_16 : _GEN_1450; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1452 = 14'h11 == parameter_2_18 ? phv_data_17 : _GEN_1451; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1453 = 14'h12 == parameter_2_18 ? phv_data_18 : _GEN_1452; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1454 = 14'h13 == parameter_2_18 ? phv_data_19 : _GEN_1453; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1455 = 14'h14 == parameter_2_18 ? phv_data_20 : _GEN_1454; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1456 = 14'h15 == parameter_2_18 ? phv_data_21 : _GEN_1455; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1457 = 14'h16 == parameter_2_18 ? phv_data_22 : _GEN_1456; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1458 = 14'h17 == parameter_2_18 ? phv_data_23 : _GEN_1457; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1459 = 14'h18 == parameter_2_18 ? phv_data_24 : _GEN_1458; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1460 = 14'h19 == parameter_2_18 ? phv_data_25 : _GEN_1459; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1461 = 14'h1a == parameter_2_18 ? phv_data_26 : _GEN_1460; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1462 = 14'h1b == parameter_2_18 ? phv_data_27 : _GEN_1461; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1463 = 14'h1c == parameter_2_18 ? phv_data_28 : _GEN_1462; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1464 = 14'h1d == parameter_2_18 ? phv_data_29 : _GEN_1463; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1465 = 14'h1e == parameter_2_18 ? phv_data_30 : _GEN_1464; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1466 = 14'h1f == parameter_2_18 ? phv_data_31 : _GEN_1465; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1467 = 14'h20 == parameter_2_18 ? phv_data_32 : _GEN_1466; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1468 = 14'h21 == parameter_2_18 ? phv_data_33 : _GEN_1467; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1469 = 14'h22 == parameter_2_18 ? phv_data_34 : _GEN_1468; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1470 = 14'h23 == parameter_2_18 ? phv_data_35 : _GEN_1469; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1471 = 14'h24 == parameter_2_18 ? phv_data_36 : _GEN_1470; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1472 = 14'h25 == parameter_2_18 ? phv_data_37 : _GEN_1471; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1473 = 14'h26 == parameter_2_18 ? phv_data_38 : _GEN_1472; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1474 = 14'h27 == parameter_2_18 ? phv_data_39 : _GEN_1473; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1475 = 14'h28 == parameter_2_18 ? phv_data_40 : _GEN_1474; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1476 = 14'h29 == parameter_2_18 ? phv_data_41 : _GEN_1475; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1477 = 14'h2a == parameter_2_18 ? phv_data_42 : _GEN_1476; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1478 = 14'h2b == parameter_2_18 ? phv_data_43 : _GEN_1477; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1479 = 14'h2c == parameter_2_18 ? phv_data_44 : _GEN_1478; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1480 = 14'h2d == parameter_2_18 ? phv_data_45 : _GEN_1479; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1481 = 14'h2e == parameter_2_18 ? phv_data_46 : _GEN_1480; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1482 = 14'h2f == parameter_2_18 ? phv_data_47 : _GEN_1481; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1483 = 14'h30 == parameter_2_18 ? phv_data_48 : _GEN_1482; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1484 = 14'h31 == parameter_2_18 ? phv_data_49 : _GEN_1483; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1485 = 14'h32 == parameter_2_18 ? phv_data_50 : _GEN_1484; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1486 = 14'h33 == parameter_2_18 ? phv_data_51 : _GEN_1485; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1487 = 14'h34 == parameter_2_18 ? phv_data_52 : _GEN_1486; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1488 = 14'h35 == parameter_2_18 ? phv_data_53 : _GEN_1487; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1489 = 14'h36 == parameter_2_18 ? phv_data_54 : _GEN_1488; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1490 = 14'h37 == parameter_2_18 ? phv_data_55 : _GEN_1489; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1491 = 14'h38 == parameter_2_18 ? phv_data_56 : _GEN_1490; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1492 = 14'h39 == parameter_2_18 ? phv_data_57 : _GEN_1491; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1493 = 14'h3a == parameter_2_18 ? phv_data_58 : _GEN_1492; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1494 = 14'h3b == parameter_2_18 ? phv_data_59 : _GEN_1493; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1495 = 14'h3c == parameter_2_18 ? phv_data_60 : _GEN_1494; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1496 = 14'h3d == parameter_2_18 ? phv_data_61 : _GEN_1495; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1497 = 14'h3e == parameter_2_18 ? phv_data_62 : _GEN_1496; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1498 = 14'h3f == parameter_2_18 ? phv_data_63 : _GEN_1497; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_19 = vliw_19[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_19 = vliw_19[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_19 = parameter_2_19[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_19 = parameter_2_19[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_19 = {{1'd0}, args_offset_19}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_19 = _total_offset_T_19[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1502 = 3'h1 == total_offset_19 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1503 = 3'h2 == total_offset_19 ? args_2 : _GEN_1502; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1504 = 3'h3 == total_offset_19 ? args_3 : _GEN_1503; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1505 = 3'h4 == total_offset_19 ? args_4 : _GEN_1504; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1506 = 3'h5 == total_offset_19 ? args_5 : _GEN_1505; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1507 = 3'h6 == total_offset_19 ? args_6 : _GEN_1506; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1508 = total_offset_19 < 3'h7 ? _GEN_1507 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_19_0 = 3'h0 < args_length_19 ? _GEN_1508 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_1510 = opcode_19 == 4'ha ? field_bytes_19_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1511 = opcode_19 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1352 = opcode_19 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_39 = _T_1352 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_1512 = opcode_19 == 4'h8 | opcode_19 == 4'hb ? parameter_2_19[7:0] : _GEN_1510; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_1513 = opcode_19 == 4'h8 | opcode_19 == 4'hb ? _field_tag_T_39 : _GEN_1511; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_1514 = 14'h0 == parameter_2_19 ? phv_data_0 : _GEN_1512; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1515 = 14'h1 == parameter_2_19 ? phv_data_1 : _GEN_1514; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1516 = 14'h2 == parameter_2_19 ? phv_data_2 : _GEN_1515; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1517 = 14'h3 == parameter_2_19 ? phv_data_3 : _GEN_1516; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1518 = 14'h4 == parameter_2_19 ? phv_data_4 : _GEN_1517; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1519 = 14'h5 == parameter_2_19 ? phv_data_5 : _GEN_1518; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1520 = 14'h6 == parameter_2_19 ? phv_data_6 : _GEN_1519; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1521 = 14'h7 == parameter_2_19 ? phv_data_7 : _GEN_1520; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1522 = 14'h8 == parameter_2_19 ? phv_data_8 : _GEN_1521; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1523 = 14'h9 == parameter_2_19 ? phv_data_9 : _GEN_1522; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1524 = 14'ha == parameter_2_19 ? phv_data_10 : _GEN_1523; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1525 = 14'hb == parameter_2_19 ? phv_data_11 : _GEN_1524; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1526 = 14'hc == parameter_2_19 ? phv_data_12 : _GEN_1525; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1527 = 14'hd == parameter_2_19 ? phv_data_13 : _GEN_1526; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1528 = 14'he == parameter_2_19 ? phv_data_14 : _GEN_1527; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1529 = 14'hf == parameter_2_19 ? phv_data_15 : _GEN_1528; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1530 = 14'h10 == parameter_2_19 ? phv_data_16 : _GEN_1529; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1531 = 14'h11 == parameter_2_19 ? phv_data_17 : _GEN_1530; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1532 = 14'h12 == parameter_2_19 ? phv_data_18 : _GEN_1531; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1533 = 14'h13 == parameter_2_19 ? phv_data_19 : _GEN_1532; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1534 = 14'h14 == parameter_2_19 ? phv_data_20 : _GEN_1533; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1535 = 14'h15 == parameter_2_19 ? phv_data_21 : _GEN_1534; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1536 = 14'h16 == parameter_2_19 ? phv_data_22 : _GEN_1535; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1537 = 14'h17 == parameter_2_19 ? phv_data_23 : _GEN_1536; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1538 = 14'h18 == parameter_2_19 ? phv_data_24 : _GEN_1537; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1539 = 14'h19 == parameter_2_19 ? phv_data_25 : _GEN_1538; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1540 = 14'h1a == parameter_2_19 ? phv_data_26 : _GEN_1539; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1541 = 14'h1b == parameter_2_19 ? phv_data_27 : _GEN_1540; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1542 = 14'h1c == parameter_2_19 ? phv_data_28 : _GEN_1541; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1543 = 14'h1d == parameter_2_19 ? phv_data_29 : _GEN_1542; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1544 = 14'h1e == parameter_2_19 ? phv_data_30 : _GEN_1543; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1545 = 14'h1f == parameter_2_19 ? phv_data_31 : _GEN_1544; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1546 = 14'h20 == parameter_2_19 ? phv_data_32 : _GEN_1545; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1547 = 14'h21 == parameter_2_19 ? phv_data_33 : _GEN_1546; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1548 = 14'h22 == parameter_2_19 ? phv_data_34 : _GEN_1547; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1549 = 14'h23 == parameter_2_19 ? phv_data_35 : _GEN_1548; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1550 = 14'h24 == parameter_2_19 ? phv_data_36 : _GEN_1549; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1551 = 14'h25 == parameter_2_19 ? phv_data_37 : _GEN_1550; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1552 = 14'h26 == parameter_2_19 ? phv_data_38 : _GEN_1551; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1553 = 14'h27 == parameter_2_19 ? phv_data_39 : _GEN_1552; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1554 = 14'h28 == parameter_2_19 ? phv_data_40 : _GEN_1553; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1555 = 14'h29 == parameter_2_19 ? phv_data_41 : _GEN_1554; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1556 = 14'h2a == parameter_2_19 ? phv_data_42 : _GEN_1555; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1557 = 14'h2b == parameter_2_19 ? phv_data_43 : _GEN_1556; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1558 = 14'h2c == parameter_2_19 ? phv_data_44 : _GEN_1557; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1559 = 14'h2d == parameter_2_19 ? phv_data_45 : _GEN_1558; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1560 = 14'h2e == parameter_2_19 ? phv_data_46 : _GEN_1559; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1561 = 14'h2f == parameter_2_19 ? phv_data_47 : _GEN_1560; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1562 = 14'h30 == parameter_2_19 ? phv_data_48 : _GEN_1561; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1563 = 14'h31 == parameter_2_19 ? phv_data_49 : _GEN_1562; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1564 = 14'h32 == parameter_2_19 ? phv_data_50 : _GEN_1563; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1565 = 14'h33 == parameter_2_19 ? phv_data_51 : _GEN_1564; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1566 = 14'h34 == parameter_2_19 ? phv_data_52 : _GEN_1565; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1567 = 14'h35 == parameter_2_19 ? phv_data_53 : _GEN_1566; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1568 = 14'h36 == parameter_2_19 ? phv_data_54 : _GEN_1567; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1569 = 14'h37 == parameter_2_19 ? phv_data_55 : _GEN_1568; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1570 = 14'h38 == parameter_2_19 ? phv_data_56 : _GEN_1569; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1571 = 14'h39 == parameter_2_19 ? phv_data_57 : _GEN_1570; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1572 = 14'h3a == parameter_2_19 ? phv_data_58 : _GEN_1571; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1573 = 14'h3b == parameter_2_19 ? phv_data_59 : _GEN_1572; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1574 = 14'h3c == parameter_2_19 ? phv_data_60 : _GEN_1573; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1575 = 14'h3d == parameter_2_19 ? phv_data_61 : _GEN_1574; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1576 = 14'h3e == parameter_2_19 ? phv_data_62 : _GEN_1575; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1577 = 14'h3f == parameter_2_19 ? phv_data_63 : _GEN_1576; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_20 = vliw_20[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_20 = vliw_20[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_20 = parameter_2_20[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_20 = parameter_2_20[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_20 = {{1'd0}, args_offset_20}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_20 = _total_offset_T_20[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1581 = 3'h1 == total_offset_20 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1582 = 3'h2 == total_offset_20 ? args_2 : _GEN_1581; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1583 = 3'h3 == total_offset_20 ? args_3 : _GEN_1582; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1584 = 3'h4 == total_offset_20 ? args_4 : _GEN_1583; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1585 = 3'h5 == total_offset_20 ? args_5 : _GEN_1584; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1586 = 3'h6 == total_offset_20 ? args_6 : _GEN_1585; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1587 = total_offset_20 < 3'h7 ? _GEN_1586 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_20_0 = 3'h0 < args_length_20 ? _GEN_1587 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_1589 = opcode_20 == 4'ha ? field_bytes_20_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1590 = opcode_20 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1423 = opcode_20 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_41 = _T_1423 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_1591 = opcode_20 == 4'h8 | opcode_20 == 4'hb ? parameter_2_20[7:0] : _GEN_1589; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_1592 = opcode_20 == 4'h8 | opcode_20 == 4'hb ? _field_tag_T_41 : _GEN_1590; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_1593 = 14'h0 == parameter_2_20 ? phv_data_0 : _GEN_1591; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1594 = 14'h1 == parameter_2_20 ? phv_data_1 : _GEN_1593; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1595 = 14'h2 == parameter_2_20 ? phv_data_2 : _GEN_1594; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1596 = 14'h3 == parameter_2_20 ? phv_data_3 : _GEN_1595; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1597 = 14'h4 == parameter_2_20 ? phv_data_4 : _GEN_1596; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1598 = 14'h5 == parameter_2_20 ? phv_data_5 : _GEN_1597; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1599 = 14'h6 == parameter_2_20 ? phv_data_6 : _GEN_1598; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1600 = 14'h7 == parameter_2_20 ? phv_data_7 : _GEN_1599; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1601 = 14'h8 == parameter_2_20 ? phv_data_8 : _GEN_1600; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1602 = 14'h9 == parameter_2_20 ? phv_data_9 : _GEN_1601; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1603 = 14'ha == parameter_2_20 ? phv_data_10 : _GEN_1602; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1604 = 14'hb == parameter_2_20 ? phv_data_11 : _GEN_1603; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1605 = 14'hc == parameter_2_20 ? phv_data_12 : _GEN_1604; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1606 = 14'hd == parameter_2_20 ? phv_data_13 : _GEN_1605; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1607 = 14'he == parameter_2_20 ? phv_data_14 : _GEN_1606; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1608 = 14'hf == parameter_2_20 ? phv_data_15 : _GEN_1607; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1609 = 14'h10 == parameter_2_20 ? phv_data_16 : _GEN_1608; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1610 = 14'h11 == parameter_2_20 ? phv_data_17 : _GEN_1609; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1611 = 14'h12 == parameter_2_20 ? phv_data_18 : _GEN_1610; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1612 = 14'h13 == parameter_2_20 ? phv_data_19 : _GEN_1611; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1613 = 14'h14 == parameter_2_20 ? phv_data_20 : _GEN_1612; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1614 = 14'h15 == parameter_2_20 ? phv_data_21 : _GEN_1613; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1615 = 14'h16 == parameter_2_20 ? phv_data_22 : _GEN_1614; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1616 = 14'h17 == parameter_2_20 ? phv_data_23 : _GEN_1615; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1617 = 14'h18 == parameter_2_20 ? phv_data_24 : _GEN_1616; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1618 = 14'h19 == parameter_2_20 ? phv_data_25 : _GEN_1617; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1619 = 14'h1a == parameter_2_20 ? phv_data_26 : _GEN_1618; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1620 = 14'h1b == parameter_2_20 ? phv_data_27 : _GEN_1619; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1621 = 14'h1c == parameter_2_20 ? phv_data_28 : _GEN_1620; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1622 = 14'h1d == parameter_2_20 ? phv_data_29 : _GEN_1621; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1623 = 14'h1e == parameter_2_20 ? phv_data_30 : _GEN_1622; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1624 = 14'h1f == parameter_2_20 ? phv_data_31 : _GEN_1623; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1625 = 14'h20 == parameter_2_20 ? phv_data_32 : _GEN_1624; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1626 = 14'h21 == parameter_2_20 ? phv_data_33 : _GEN_1625; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1627 = 14'h22 == parameter_2_20 ? phv_data_34 : _GEN_1626; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1628 = 14'h23 == parameter_2_20 ? phv_data_35 : _GEN_1627; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1629 = 14'h24 == parameter_2_20 ? phv_data_36 : _GEN_1628; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1630 = 14'h25 == parameter_2_20 ? phv_data_37 : _GEN_1629; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1631 = 14'h26 == parameter_2_20 ? phv_data_38 : _GEN_1630; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1632 = 14'h27 == parameter_2_20 ? phv_data_39 : _GEN_1631; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1633 = 14'h28 == parameter_2_20 ? phv_data_40 : _GEN_1632; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1634 = 14'h29 == parameter_2_20 ? phv_data_41 : _GEN_1633; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1635 = 14'h2a == parameter_2_20 ? phv_data_42 : _GEN_1634; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1636 = 14'h2b == parameter_2_20 ? phv_data_43 : _GEN_1635; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1637 = 14'h2c == parameter_2_20 ? phv_data_44 : _GEN_1636; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1638 = 14'h2d == parameter_2_20 ? phv_data_45 : _GEN_1637; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1639 = 14'h2e == parameter_2_20 ? phv_data_46 : _GEN_1638; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1640 = 14'h2f == parameter_2_20 ? phv_data_47 : _GEN_1639; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1641 = 14'h30 == parameter_2_20 ? phv_data_48 : _GEN_1640; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1642 = 14'h31 == parameter_2_20 ? phv_data_49 : _GEN_1641; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1643 = 14'h32 == parameter_2_20 ? phv_data_50 : _GEN_1642; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1644 = 14'h33 == parameter_2_20 ? phv_data_51 : _GEN_1643; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1645 = 14'h34 == parameter_2_20 ? phv_data_52 : _GEN_1644; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1646 = 14'h35 == parameter_2_20 ? phv_data_53 : _GEN_1645; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1647 = 14'h36 == parameter_2_20 ? phv_data_54 : _GEN_1646; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1648 = 14'h37 == parameter_2_20 ? phv_data_55 : _GEN_1647; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1649 = 14'h38 == parameter_2_20 ? phv_data_56 : _GEN_1648; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1650 = 14'h39 == parameter_2_20 ? phv_data_57 : _GEN_1649; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1651 = 14'h3a == parameter_2_20 ? phv_data_58 : _GEN_1650; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1652 = 14'h3b == parameter_2_20 ? phv_data_59 : _GEN_1651; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1653 = 14'h3c == parameter_2_20 ? phv_data_60 : _GEN_1652; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1654 = 14'h3d == parameter_2_20 ? phv_data_61 : _GEN_1653; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1655 = 14'h3e == parameter_2_20 ? phv_data_62 : _GEN_1654; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1656 = 14'h3f == parameter_2_20 ? phv_data_63 : _GEN_1655; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_21 = vliw_21[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_21 = vliw_21[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_21 = parameter_2_21[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_21 = parameter_2_21[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_21 = {{1'd0}, args_offset_21}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_21 = _total_offset_T_21[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1660 = 3'h1 == total_offset_21 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1661 = 3'h2 == total_offset_21 ? args_2 : _GEN_1660; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1662 = 3'h3 == total_offset_21 ? args_3 : _GEN_1661; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1663 = 3'h4 == total_offset_21 ? args_4 : _GEN_1662; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1664 = 3'h5 == total_offset_21 ? args_5 : _GEN_1663; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1665 = 3'h6 == total_offset_21 ? args_6 : _GEN_1664; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1666 = total_offset_21 < 3'h7 ? _GEN_1665 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_21_0 = 3'h0 < args_length_21 ? _GEN_1666 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_1668 = opcode_21 == 4'ha ? field_bytes_21_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1669 = opcode_21 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1494 = opcode_21 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_43 = _T_1494 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_1670 = opcode_21 == 4'h8 | opcode_21 == 4'hb ? parameter_2_21[7:0] : _GEN_1668; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_1671 = opcode_21 == 4'h8 | opcode_21 == 4'hb ? _field_tag_T_43 : _GEN_1669; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_1672 = 14'h0 == parameter_2_21 ? phv_data_0 : _GEN_1670; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1673 = 14'h1 == parameter_2_21 ? phv_data_1 : _GEN_1672; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1674 = 14'h2 == parameter_2_21 ? phv_data_2 : _GEN_1673; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1675 = 14'h3 == parameter_2_21 ? phv_data_3 : _GEN_1674; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1676 = 14'h4 == parameter_2_21 ? phv_data_4 : _GEN_1675; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1677 = 14'h5 == parameter_2_21 ? phv_data_5 : _GEN_1676; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1678 = 14'h6 == parameter_2_21 ? phv_data_6 : _GEN_1677; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1679 = 14'h7 == parameter_2_21 ? phv_data_7 : _GEN_1678; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1680 = 14'h8 == parameter_2_21 ? phv_data_8 : _GEN_1679; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1681 = 14'h9 == parameter_2_21 ? phv_data_9 : _GEN_1680; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1682 = 14'ha == parameter_2_21 ? phv_data_10 : _GEN_1681; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1683 = 14'hb == parameter_2_21 ? phv_data_11 : _GEN_1682; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1684 = 14'hc == parameter_2_21 ? phv_data_12 : _GEN_1683; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1685 = 14'hd == parameter_2_21 ? phv_data_13 : _GEN_1684; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1686 = 14'he == parameter_2_21 ? phv_data_14 : _GEN_1685; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1687 = 14'hf == parameter_2_21 ? phv_data_15 : _GEN_1686; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1688 = 14'h10 == parameter_2_21 ? phv_data_16 : _GEN_1687; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1689 = 14'h11 == parameter_2_21 ? phv_data_17 : _GEN_1688; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1690 = 14'h12 == parameter_2_21 ? phv_data_18 : _GEN_1689; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1691 = 14'h13 == parameter_2_21 ? phv_data_19 : _GEN_1690; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1692 = 14'h14 == parameter_2_21 ? phv_data_20 : _GEN_1691; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1693 = 14'h15 == parameter_2_21 ? phv_data_21 : _GEN_1692; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1694 = 14'h16 == parameter_2_21 ? phv_data_22 : _GEN_1693; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1695 = 14'h17 == parameter_2_21 ? phv_data_23 : _GEN_1694; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1696 = 14'h18 == parameter_2_21 ? phv_data_24 : _GEN_1695; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1697 = 14'h19 == parameter_2_21 ? phv_data_25 : _GEN_1696; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1698 = 14'h1a == parameter_2_21 ? phv_data_26 : _GEN_1697; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1699 = 14'h1b == parameter_2_21 ? phv_data_27 : _GEN_1698; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1700 = 14'h1c == parameter_2_21 ? phv_data_28 : _GEN_1699; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1701 = 14'h1d == parameter_2_21 ? phv_data_29 : _GEN_1700; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1702 = 14'h1e == parameter_2_21 ? phv_data_30 : _GEN_1701; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1703 = 14'h1f == parameter_2_21 ? phv_data_31 : _GEN_1702; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1704 = 14'h20 == parameter_2_21 ? phv_data_32 : _GEN_1703; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1705 = 14'h21 == parameter_2_21 ? phv_data_33 : _GEN_1704; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1706 = 14'h22 == parameter_2_21 ? phv_data_34 : _GEN_1705; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1707 = 14'h23 == parameter_2_21 ? phv_data_35 : _GEN_1706; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1708 = 14'h24 == parameter_2_21 ? phv_data_36 : _GEN_1707; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1709 = 14'h25 == parameter_2_21 ? phv_data_37 : _GEN_1708; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1710 = 14'h26 == parameter_2_21 ? phv_data_38 : _GEN_1709; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1711 = 14'h27 == parameter_2_21 ? phv_data_39 : _GEN_1710; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1712 = 14'h28 == parameter_2_21 ? phv_data_40 : _GEN_1711; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1713 = 14'h29 == parameter_2_21 ? phv_data_41 : _GEN_1712; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1714 = 14'h2a == parameter_2_21 ? phv_data_42 : _GEN_1713; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1715 = 14'h2b == parameter_2_21 ? phv_data_43 : _GEN_1714; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1716 = 14'h2c == parameter_2_21 ? phv_data_44 : _GEN_1715; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1717 = 14'h2d == parameter_2_21 ? phv_data_45 : _GEN_1716; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1718 = 14'h2e == parameter_2_21 ? phv_data_46 : _GEN_1717; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1719 = 14'h2f == parameter_2_21 ? phv_data_47 : _GEN_1718; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1720 = 14'h30 == parameter_2_21 ? phv_data_48 : _GEN_1719; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1721 = 14'h31 == parameter_2_21 ? phv_data_49 : _GEN_1720; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1722 = 14'h32 == parameter_2_21 ? phv_data_50 : _GEN_1721; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1723 = 14'h33 == parameter_2_21 ? phv_data_51 : _GEN_1722; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1724 = 14'h34 == parameter_2_21 ? phv_data_52 : _GEN_1723; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1725 = 14'h35 == parameter_2_21 ? phv_data_53 : _GEN_1724; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1726 = 14'h36 == parameter_2_21 ? phv_data_54 : _GEN_1725; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1727 = 14'h37 == parameter_2_21 ? phv_data_55 : _GEN_1726; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1728 = 14'h38 == parameter_2_21 ? phv_data_56 : _GEN_1727; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1729 = 14'h39 == parameter_2_21 ? phv_data_57 : _GEN_1728; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1730 = 14'h3a == parameter_2_21 ? phv_data_58 : _GEN_1729; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1731 = 14'h3b == parameter_2_21 ? phv_data_59 : _GEN_1730; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1732 = 14'h3c == parameter_2_21 ? phv_data_60 : _GEN_1731; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1733 = 14'h3d == parameter_2_21 ? phv_data_61 : _GEN_1732; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1734 = 14'h3e == parameter_2_21 ? phv_data_62 : _GEN_1733; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1735 = 14'h3f == parameter_2_21 ? phv_data_63 : _GEN_1734; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_22 = vliw_22[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_22 = vliw_22[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_22 = parameter_2_22[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_22 = parameter_2_22[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_22 = {{1'd0}, args_offset_22}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_22 = _total_offset_T_22[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1739 = 3'h1 == total_offset_22 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1740 = 3'h2 == total_offset_22 ? args_2 : _GEN_1739; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1741 = 3'h3 == total_offset_22 ? args_3 : _GEN_1740; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1742 = 3'h4 == total_offset_22 ? args_4 : _GEN_1741; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1743 = 3'h5 == total_offset_22 ? args_5 : _GEN_1742; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1744 = 3'h6 == total_offset_22 ? args_6 : _GEN_1743; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1745 = total_offset_22 < 3'h7 ? _GEN_1744 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_22_0 = 3'h0 < args_length_22 ? _GEN_1745 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_1747 = opcode_22 == 4'ha ? field_bytes_22_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1748 = opcode_22 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1565 = opcode_22 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_45 = _T_1565 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_1749 = opcode_22 == 4'h8 | opcode_22 == 4'hb ? parameter_2_22[7:0] : _GEN_1747; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_1750 = opcode_22 == 4'h8 | opcode_22 == 4'hb ? _field_tag_T_45 : _GEN_1748; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_1751 = 14'h0 == parameter_2_22 ? phv_data_0 : _GEN_1749; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1752 = 14'h1 == parameter_2_22 ? phv_data_1 : _GEN_1751; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1753 = 14'h2 == parameter_2_22 ? phv_data_2 : _GEN_1752; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1754 = 14'h3 == parameter_2_22 ? phv_data_3 : _GEN_1753; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1755 = 14'h4 == parameter_2_22 ? phv_data_4 : _GEN_1754; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1756 = 14'h5 == parameter_2_22 ? phv_data_5 : _GEN_1755; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1757 = 14'h6 == parameter_2_22 ? phv_data_6 : _GEN_1756; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1758 = 14'h7 == parameter_2_22 ? phv_data_7 : _GEN_1757; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1759 = 14'h8 == parameter_2_22 ? phv_data_8 : _GEN_1758; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1760 = 14'h9 == parameter_2_22 ? phv_data_9 : _GEN_1759; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1761 = 14'ha == parameter_2_22 ? phv_data_10 : _GEN_1760; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1762 = 14'hb == parameter_2_22 ? phv_data_11 : _GEN_1761; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1763 = 14'hc == parameter_2_22 ? phv_data_12 : _GEN_1762; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1764 = 14'hd == parameter_2_22 ? phv_data_13 : _GEN_1763; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1765 = 14'he == parameter_2_22 ? phv_data_14 : _GEN_1764; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1766 = 14'hf == parameter_2_22 ? phv_data_15 : _GEN_1765; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1767 = 14'h10 == parameter_2_22 ? phv_data_16 : _GEN_1766; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1768 = 14'h11 == parameter_2_22 ? phv_data_17 : _GEN_1767; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1769 = 14'h12 == parameter_2_22 ? phv_data_18 : _GEN_1768; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1770 = 14'h13 == parameter_2_22 ? phv_data_19 : _GEN_1769; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1771 = 14'h14 == parameter_2_22 ? phv_data_20 : _GEN_1770; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1772 = 14'h15 == parameter_2_22 ? phv_data_21 : _GEN_1771; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1773 = 14'h16 == parameter_2_22 ? phv_data_22 : _GEN_1772; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1774 = 14'h17 == parameter_2_22 ? phv_data_23 : _GEN_1773; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1775 = 14'h18 == parameter_2_22 ? phv_data_24 : _GEN_1774; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1776 = 14'h19 == parameter_2_22 ? phv_data_25 : _GEN_1775; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1777 = 14'h1a == parameter_2_22 ? phv_data_26 : _GEN_1776; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1778 = 14'h1b == parameter_2_22 ? phv_data_27 : _GEN_1777; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1779 = 14'h1c == parameter_2_22 ? phv_data_28 : _GEN_1778; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1780 = 14'h1d == parameter_2_22 ? phv_data_29 : _GEN_1779; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1781 = 14'h1e == parameter_2_22 ? phv_data_30 : _GEN_1780; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1782 = 14'h1f == parameter_2_22 ? phv_data_31 : _GEN_1781; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1783 = 14'h20 == parameter_2_22 ? phv_data_32 : _GEN_1782; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1784 = 14'h21 == parameter_2_22 ? phv_data_33 : _GEN_1783; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1785 = 14'h22 == parameter_2_22 ? phv_data_34 : _GEN_1784; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1786 = 14'h23 == parameter_2_22 ? phv_data_35 : _GEN_1785; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1787 = 14'h24 == parameter_2_22 ? phv_data_36 : _GEN_1786; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1788 = 14'h25 == parameter_2_22 ? phv_data_37 : _GEN_1787; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1789 = 14'h26 == parameter_2_22 ? phv_data_38 : _GEN_1788; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1790 = 14'h27 == parameter_2_22 ? phv_data_39 : _GEN_1789; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1791 = 14'h28 == parameter_2_22 ? phv_data_40 : _GEN_1790; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1792 = 14'h29 == parameter_2_22 ? phv_data_41 : _GEN_1791; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1793 = 14'h2a == parameter_2_22 ? phv_data_42 : _GEN_1792; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1794 = 14'h2b == parameter_2_22 ? phv_data_43 : _GEN_1793; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1795 = 14'h2c == parameter_2_22 ? phv_data_44 : _GEN_1794; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1796 = 14'h2d == parameter_2_22 ? phv_data_45 : _GEN_1795; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1797 = 14'h2e == parameter_2_22 ? phv_data_46 : _GEN_1796; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1798 = 14'h2f == parameter_2_22 ? phv_data_47 : _GEN_1797; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1799 = 14'h30 == parameter_2_22 ? phv_data_48 : _GEN_1798; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1800 = 14'h31 == parameter_2_22 ? phv_data_49 : _GEN_1799; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1801 = 14'h32 == parameter_2_22 ? phv_data_50 : _GEN_1800; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1802 = 14'h33 == parameter_2_22 ? phv_data_51 : _GEN_1801; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1803 = 14'h34 == parameter_2_22 ? phv_data_52 : _GEN_1802; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1804 = 14'h35 == parameter_2_22 ? phv_data_53 : _GEN_1803; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1805 = 14'h36 == parameter_2_22 ? phv_data_54 : _GEN_1804; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1806 = 14'h37 == parameter_2_22 ? phv_data_55 : _GEN_1805; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1807 = 14'h38 == parameter_2_22 ? phv_data_56 : _GEN_1806; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1808 = 14'h39 == parameter_2_22 ? phv_data_57 : _GEN_1807; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1809 = 14'h3a == parameter_2_22 ? phv_data_58 : _GEN_1808; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1810 = 14'h3b == parameter_2_22 ? phv_data_59 : _GEN_1809; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1811 = 14'h3c == parameter_2_22 ? phv_data_60 : _GEN_1810; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1812 = 14'h3d == parameter_2_22 ? phv_data_61 : _GEN_1811; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1813 = 14'h3e == parameter_2_22 ? phv_data_62 : _GEN_1812; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1814 = 14'h3f == parameter_2_22 ? phv_data_63 : _GEN_1813; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_23 = vliw_23[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_23 = vliw_23[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_23 = parameter_2_23[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_23 = parameter_2_23[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_23 = {{1'd0}, args_offset_23}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_23 = _total_offset_T_23[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1818 = 3'h1 == total_offset_23 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1819 = 3'h2 == total_offset_23 ? args_2 : _GEN_1818; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1820 = 3'h3 == total_offset_23 ? args_3 : _GEN_1819; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1821 = 3'h4 == total_offset_23 ? args_4 : _GEN_1820; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1822 = 3'h5 == total_offset_23 ? args_5 : _GEN_1821; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1823 = 3'h6 == total_offset_23 ? args_6 : _GEN_1822; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1824 = total_offset_23 < 3'h7 ? _GEN_1823 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_23_0 = 3'h0 < args_length_23 ? _GEN_1824 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_1826 = opcode_23 == 4'ha ? field_bytes_23_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1827 = opcode_23 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1636 = opcode_23 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_47 = _T_1636 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_1828 = opcode_23 == 4'h8 | opcode_23 == 4'hb ? parameter_2_23[7:0] : _GEN_1826; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_1829 = opcode_23 == 4'h8 | opcode_23 == 4'hb ? _field_tag_T_47 : _GEN_1827; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_1830 = 14'h0 == parameter_2_23 ? phv_data_0 : _GEN_1828; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1831 = 14'h1 == parameter_2_23 ? phv_data_1 : _GEN_1830; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1832 = 14'h2 == parameter_2_23 ? phv_data_2 : _GEN_1831; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1833 = 14'h3 == parameter_2_23 ? phv_data_3 : _GEN_1832; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1834 = 14'h4 == parameter_2_23 ? phv_data_4 : _GEN_1833; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1835 = 14'h5 == parameter_2_23 ? phv_data_5 : _GEN_1834; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1836 = 14'h6 == parameter_2_23 ? phv_data_6 : _GEN_1835; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1837 = 14'h7 == parameter_2_23 ? phv_data_7 : _GEN_1836; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1838 = 14'h8 == parameter_2_23 ? phv_data_8 : _GEN_1837; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1839 = 14'h9 == parameter_2_23 ? phv_data_9 : _GEN_1838; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1840 = 14'ha == parameter_2_23 ? phv_data_10 : _GEN_1839; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1841 = 14'hb == parameter_2_23 ? phv_data_11 : _GEN_1840; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1842 = 14'hc == parameter_2_23 ? phv_data_12 : _GEN_1841; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1843 = 14'hd == parameter_2_23 ? phv_data_13 : _GEN_1842; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1844 = 14'he == parameter_2_23 ? phv_data_14 : _GEN_1843; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1845 = 14'hf == parameter_2_23 ? phv_data_15 : _GEN_1844; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1846 = 14'h10 == parameter_2_23 ? phv_data_16 : _GEN_1845; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1847 = 14'h11 == parameter_2_23 ? phv_data_17 : _GEN_1846; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1848 = 14'h12 == parameter_2_23 ? phv_data_18 : _GEN_1847; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1849 = 14'h13 == parameter_2_23 ? phv_data_19 : _GEN_1848; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1850 = 14'h14 == parameter_2_23 ? phv_data_20 : _GEN_1849; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1851 = 14'h15 == parameter_2_23 ? phv_data_21 : _GEN_1850; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1852 = 14'h16 == parameter_2_23 ? phv_data_22 : _GEN_1851; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1853 = 14'h17 == parameter_2_23 ? phv_data_23 : _GEN_1852; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1854 = 14'h18 == parameter_2_23 ? phv_data_24 : _GEN_1853; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1855 = 14'h19 == parameter_2_23 ? phv_data_25 : _GEN_1854; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1856 = 14'h1a == parameter_2_23 ? phv_data_26 : _GEN_1855; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1857 = 14'h1b == parameter_2_23 ? phv_data_27 : _GEN_1856; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1858 = 14'h1c == parameter_2_23 ? phv_data_28 : _GEN_1857; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1859 = 14'h1d == parameter_2_23 ? phv_data_29 : _GEN_1858; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1860 = 14'h1e == parameter_2_23 ? phv_data_30 : _GEN_1859; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1861 = 14'h1f == parameter_2_23 ? phv_data_31 : _GEN_1860; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1862 = 14'h20 == parameter_2_23 ? phv_data_32 : _GEN_1861; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1863 = 14'h21 == parameter_2_23 ? phv_data_33 : _GEN_1862; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1864 = 14'h22 == parameter_2_23 ? phv_data_34 : _GEN_1863; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1865 = 14'h23 == parameter_2_23 ? phv_data_35 : _GEN_1864; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1866 = 14'h24 == parameter_2_23 ? phv_data_36 : _GEN_1865; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1867 = 14'h25 == parameter_2_23 ? phv_data_37 : _GEN_1866; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1868 = 14'h26 == parameter_2_23 ? phv_data_38 : _GEN_1867; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1869 = 14'h27 == parameter_2_23 ? phv_data_39 : _GEN_1868; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1870 = 14'h28 == parameter_2_23 ? phv_data_40 : _GEN_1869; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1871 = 14'h29 == parameter_2_23 ? phv_data_41 : _GEN_1870; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1872 = 14'h2a == parameter_2_23 ? phv_data_42 : _GEN_1871; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1873 = 14'h2b == parameter_2_23 ? phv_data_43 : _GEN_1872; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1874 = 14'h2c == parameter_2_23 ? phv_data_44 : _GEN_1873; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1875 = 14'h2d == parameter_2_23 ? phv_data_45 : _GEN_1874; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1876 = 14'h2e == parameter_2_23 ? phv_data_46 : _GEN_1875; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1877 = 14'h2f == parameter_2_23 ? phv_data_47 : _GEN_1876; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1878 = 14'h30 == parameter_2_23 ? phv_data_48 : _GEN_1877; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1879 = 14'h31 == parameter_2_23 ? phv_data_49 : _GEN_1878; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1880 = 14'h32 == parameter_2_23 ? phv_data_50 : _GEN_1879; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1881 = 14'h33 == parameter_2_23 ? phv_data_51 : _GEN_1880; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1882 = 14'h34 == parameter_2_23 ? phv_data_52 : _GEN_1881; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1883 = 14'h35 == parameter_2_23 ? phv_data_53 : _GEN_1882; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1884 = 14'h36 == parameter_2_23 ? phv_data_54 : _GEN_1883; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1885 = 14'h37 == parameter_2_23 ? phv_data_55 : _GEN_1884; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1886 = 14'h38 == parameter_2_23 ? phv_data_56 : _GEN_1885; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1887 = 14'h39 == parameter_2_23 ? phv_data_57 : _GEN_1886; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1888 = 14'h3a == parameter_2_23 ? phv_data_58 : _GEN_1887; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1889 = 14'h3b == parameter_2_23 ? phv_data_59 : _GEN_1888; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1890 = 14'h3c == parameter_2_23 ? phv_data_60 : _GEN_1889; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1891 = 14'h3d == parameter_2_23 ? phv_data_61 : _GEN_1890; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1892 = 14'h3e == parameter_2_23 ? phv_data_62 : _GEN_1891; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1893 = 14'h3f == parameter_2_23 ? phv_data_63 : _GEN_1892; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_24 = vliw_24[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_24 = vliw_24[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_24 = parameter_2_24[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_24 = parameter_2_24[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_24 = {{1'd0}, args_offset_24}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_24 = _total_offset_T_24[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1897 = 3'h1 == total_offset_24 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1898 = 3'h2 == total_offset_24 ? args_2 : _GEN_1897; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1899 = 3'h3 == total_offset_24 ? args_3 : _GEN_1898; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1900 = 3'h4 == total_offset_24 ? args_4 : _GEN_1899; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1901 = 3'h5 == total_offset_24 ? args_5 : _GEN_1900; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1902 = 3'h6 == total_offset_24 ? args_6 : _GEN_1901; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1903 = total_offset_24 < 3'h7 ? _GEN_1902 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_24_0 = 3'h0 < args_length_24 ? _GEN_1903 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_1905 = opcode_24 == 4'ha ? field_bytes_24_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1906 = opcode_24 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1707 = opcode_24 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_49 = _T_1707 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_1907 = opcode_24 == 4'h8 | opcode_24 == 4'hb ? parameter_2_24[7:0] : _GEN_1905; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_1908 = opcode_24 == 4'h8 | opcode_24 == 4'hb ? _field_tag_T_49 : _GEN_1906; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_1909 = 14'h0 == parameter_2_24 ? phv_data_0 : _GEN_1907; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1910 = 14'h1 == parameter_2_24 ? phv_data_1 : _GEN_1909; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1911 = 14'h2 == parameter_2_24 ? phv_data_2 : _GEN_1910; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1912 = 14'h3 == parameter_2_24 ? phv_data_3 : _GEN_1911; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1913 = 14'h4 == parameter_2_24 ? phv_data_4 : _GEN_1912; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1914 = 14'h5 == parameter_2_24 ? phv_data_5 : _GEN_1913; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1915 = 14'h6 == parameter_2_24 ? phv_data_6 : _GEN_1914; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1916 = 14'h7 == parameter_2_24 ? phv_data_7 : _GEN_1915; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1917 = 14'h8 == parameter_2_24 ? phv_data_8 : _GEN_1916; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1918 = 14'h9 == parameter_2_24 ? phv_data_9 : _GEN_1917; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1919 = 14'ha == parameter_2_24 ? phv_data_10 : _GEN_1918; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1920 = 14'hb == parameter_2_24 ? phv_data_11 : _GEN_1919; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1921 = 14'hc == parameter_2_24 ? phv_data_12 : _GEN_1920; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1922 = 14'hd == parameter_2_24 ? phv_data_13 : _GEN_1921; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1923 = 14'he == parameter_2_24 ? phv_data_14 : _GEN_1922; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1924 = 14'hf == parameter_2_24 ? phv_data_15 : _GEN_1923; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1925 = 14'h10 == parameter_2_24 ? phv_data_16 : _GEN_1924; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1926 = 14'h11 == parameter_2_24 ? phv_data_17 : _GEN_1925; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1927 = 14'h12 == parameter_2_24 ? phv_data_18 : _GEN_1926; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1928 = 14'h13 == parameter_2_24 ? phv_data_19 : _GEN_1927; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1929 = 14'h14 == parameter_2_24 ? phv_data_20 : _GEN_1928; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1930 = 14'h15 == parameter_2_24 ? phv_data_21 : _GEN_1929; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1931 = 14'h16 == parameter_2_24 ? phv_data_22 : _GEN_1930; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1932 = 14'h17 == parameter_2_24 ? phv_data_23 : _GEN_1931; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1933 = 14'h18 == parameter_2_24 ? phv_data_24 : _GEN_1932; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1934 = 14'h19 == parameter_2_24 ? phv_data_25 : _GEN_1933; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1935 = 14'h1a == parameter_2_24 ? phv_data_26 : _GEN_1934; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1936 = 14'h1b == parameter_2_24 ? phv_data_27 : _GEN_1935; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1937 = 14'h1c == parameter_2_24 ? phv_data_28 : _GEN_1936; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1938 = 14'h1d == parameter_2_24 ? phv_data_29 : _GEN_1937; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1939 = 14'h1e == parameter_2_24 ? phv_data_30 : _GEN_1938; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1940 = 14'h1f == parameter_2_24 ? phv_data_31 : _GEN_1939; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1941 = 14'h20 == parameter_2_24 ? phv_data_32 : _GEN_1940; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1942 = 14'h21 == parameter_2_24 ? phv_data_33 : _GEN_1941; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1943 = 14'h22 == parameter_2_24 ? phv_data_34 : _GEN_1942; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1944 = 14'h23 == parameter_2_24 ? phv_data_35 : _GEN_1943; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1945 = 14'h24 == parameter_2_24 ? phv_data_36 : _GEN_1944; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1946 = 14'h25 == parameter_2_24 ? phv_data_37 : _GEN_1945; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1947 = 14'h26 == parameter_2_24 ? phv_data_38 : _GEN_1946; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1948 = 14'h27 == parameter_2_24 ? phv_data_39 : _GEN_1947; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1949 = 14'h28 == parameter_2_24 ? phv_data_40 : _GEN_1948; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1950 = 14'h29 == parameter_2_24 ? phv_data_41 : _GEN_1949; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1951 = 14'h2a == parameter_2_24 ? phv_data_42 : _GEN_1950; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1952 = 14'h2b == parameter_2_24 ? phv_data_43 : _GEN_1951; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1953 = 14'h2c == parameter_2_24 ? phv_data_44 : _GEN_1952; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1954 = 14'h2d == parameter_2_24 ? phv_data_45 : _GEN_1953; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1955 = 14'h2e == parameter_2_24 ? phv_data_46 : _GEN_1954; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1956 = 14'h2f == parameter_2_24 ? phv_data_47 : _GEN_1955; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1957 = 14'h30 == parameter_2_24 ? phv_data_48 : _GEN_1956; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1958 = 14'h31 == parameter_2_24 ? phv_data_49 : _GEN_1957; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1959 = 14'h32 == parameter_2_24 ? phv_data_50 : _GEN_1958; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1960 = 14'h33 == parameter_2_24 ? phv_data_51 : _GEN_1959; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1961 = 14'h34 == parameter_2_24 ? phv_data_52 : _GEN_1960; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1962 = 14'h35 == parameter_2_24 ? phv_data_53 : _GEN_1961; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1963 = 14'h36 == parameter_2_24 ? phv_data_54 : _GEN_1962; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1964 = 14'h37 == parameter_2_24 ? phv_data_55 : _GEN_1963; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1965 = 14'h38 == parameter_2_24 ? phv_data_56 : _GEN_1964; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1966 = 14'h39 == parameter_2_24 ? phv_data_57 : _GEN_1965; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1967 = 14'h3a == parameter_2_24 ? phv_data_58 : _GEN_1966; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1968 = 14'h3b == parameter_2_24 ? phv_data_59 : _GEN_1967; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1969 = 14'h3c == parameter_2_24 ? phv_data_60 : _GEN_1968; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1970 = 14'h3d == parameter_2_24 ? phv_data_61 : _GEN_1969; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1971 = 14'h3e == parameter_2_24 ? phv_data_62 : _GEN_1970; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1972 = 14'h3f == parameter_2_24 ? phv_data_63 : _GEN_1971; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_25 = vliw_25[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_25 = vliw_25[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_25 = parameter_2_25[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_25 = parameter_2_25[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_25 = {{1'd0}, args_offset_25}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_25 = _total_offset_T_25[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1976 = 3'h1 == total_offset_25 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1977 = 3'h2 == total_offset_25 ? args_2 : _GEN_1976; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1978 = 3'h3 == total_offset_25 ? args_3 : _GEN_1977; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1979 = 3'h4 == total_offset_25 ? args_4 : _GEN_1978; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1980 = 3'h5 == total_offset_25 ? args_5 : _GEN_1979; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1981 = 3'h6 == total_offset_25 ? args_6 : _GEN_1980; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1982 = total_offset_25 < 3'h7 ? _GEN_1981 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_25_0 = 3'h0 < args_length_25 ? _GEN_1982 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_1984 = opcode_25 == 4'ha ? field_bytes_25_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1985 = opcode_25 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1778 = opcode_25 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_51 = _T_1778 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_1986 = opcode_25 == 4'h8 | opcode_25 == 4'hb ? parameter_2_25[7:0] : _GEN_1984; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_1987 = opcode_25 == 4'h8 | opcode_25 == 4'hb ? _field_tag_T_51 : _GEN_1985; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_1988 = 14'h0 == parameter_2_25 ? phv_data_0 : _GEN_1986; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1989 = 14'h1 == parameter_2_25 ? phv_data_1 : _GEN_1988; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1990 = 14'h2 == parameter_2_25 ? phv_data_2 : _GEN_1989; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1991 = 14'h3 == parameter_2_25 ? phv_data_3 : _GEN_1990; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1992 = 14'h4 == parameter_2_25 ? phv_data_4 : _GEN_1991; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1993 = 14'h5 == parameter_2_25 ? phv_data_5 : _GEN_1992; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1994 = 14'h6 == parameter_2_25 ? phv_data_6 : _GEN_1993; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1995 = 14'h7 == parameter_2_25 ? phv_data_7 : _GEN_1994; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1996 = 14'h8 == parameter_2_25 ? phv_data_8 : _GEN_1995; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1997 = 14'h9 == parameter_2_25 ? phv_data_9 : _GEN_1996; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1998 = 14'ha == parameter_2_25 ? phv_data_10 : _GEN_1997; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1999 = 14'hb == parameter_2_25 ? phv_data_11 : _GEN_1998; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2000 = 14'hc == parameter_2_25 ? phv_data_12 : _GEN_1999; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2001 = 14'hd == parameter_2_25 ? phv_data_13 : _GEN_2000; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2002 = 14'he == parameter_2_25 ? phv_data_14 : _GEN_2001; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2003 = 14'hf == parameter_2_25 ? phv_data_15 : _GEN_2002; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2004 = 14'h10 == parameter_2_25 ? phv_data_16 : _GEN_2003; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2005 = 14'h11 == parameter_2_25 ? phv_data_17 : _GEN_2004; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2006 = 14'h12 == parameter_2_25 ? phv_data_18 : _GEN_2005; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2007 = 14'h13 == parameter_2_25 ? phv_data_19 : _GEN_2006; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2008 = 14'h14 == parameter_2_25 ? phv_data_20 : _GEN_2007; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2009 = 14'h15 == parameter_2_25 ? phv_data_21 : _GEN_2008; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2010 = 14'h16 == parameter_2_25 ? phv_data_22 : _GEN_2009; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2011 = 14'h17 == parameter_2_25 ? phv_data_23 : _GEN_2010; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2012 = 14'h18 == parameter_2_25 ? phv_data_24 : _GEN_2011; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2013 = 14'h19 == parameter_2_25 ? phv_data_25 : _GEN_2012; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2014 = 14'h1a == parameter_2_25 ? phv_data_26 : _GEN_2013; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2015 = 14'h1b == parameter_2_25 ? phv_data_27 : _GEN_2014; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2016 = 14'h1c == parameter_2_25 ? phv_data_28 : _GEN_2015; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2017 = 14'h1d == parameter_2_25 ? phv_data_29 : _GEN_2016; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2018 = 14'h1e == parameter_2_25 ? phv_data_30 : _GEN_2017; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2019 = 14'h1f == parameter_2_25 ? phv_data_31 : _GEN_2018; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2020 = 14'h20 == parameter_2_25 ? phv_data_32 : _GEN_2019; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2021 = 14'h21 == parameter_2_25 ? phv_data_33 : _GEN_2020; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2022 = 14'h22 == parameter_2_25 ? phv_data_34 : _GEN_2021; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2023 = 14'h23 == parameter_2_25 ? phv_data_35 : _GEN_2022; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2024 = 14'h24 == parameter_2_25 ? phv_data_36 : _GEN_2023; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2025 = 14'h25 == parameter_2_25 ? phv_data_37 : _GEN_2024; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2026 = 14'h26 == parameter_2_25 ? phv_data_38 : _GEN_2025; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2027 = 14'h27 == parameter_2_25 ? phv_data_39 : _GEN_2026; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2028 = 14'h28 == parameter_2_25 ? phv_data_40 : _GEN_2027; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2029 = 14'h29 == parameter_2_25 ? phv_data_41 : _GEN_2028; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2030 = 14'h2a == parameter_2_25 ? phv_data_42 : _GEN_2029; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2031 = 14'h2b == parameter_2_25 ? phv_data_43 : _GEN_2030; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2032 = 14'h2c == parameter_2_25 ? phv_data_44 : _GEN_2031; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2033 = 14'h2d == parameter_2_25 ? phv_data_45 : _GEN_2032; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2034 = 14'h2e == parameter_2_25 ? phv_data_46 : _GEN_2033; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2035 = 14'h2f == parameter_2_25 ? phv_data_47 : _GEN_2034; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2036 = 14'h30 == parameter_2_25 ? phv_data_48 : _GEN_2035; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2037 = 14'h31 == parameter_2_25 ? phv_data_49 : _GEN_2036; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2038 = 14'h32 == parameter_2_25 ? phv_data_50 : _GEN_2037; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2039 = 14'h33 == parameter_2_25 ? phv_data_51 : _GEN_2038; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2040 = 14'h34 == parameter_2_25 ? phv_data_52 : _GEN_2039; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2041 = 14'h35 == parameter_2_25 ? phv_data_53 : _GEN_2040; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2042 = 14'h36 == parameter_2_25 ? phv_data_54 : _GEN_2041; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2043 = 14'h37 == parameter_2_25 ? phv_data_55 : _GEN_2042; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2044 = 14'h38 == parameter_2_25 ? phv_data_56 : _GEN_2043; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2045 = 14'h39 == parameter_2_25 ? phv_data_57 : _GEN_2044; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2046 = 14'h3a == parameter_2_25 ? phv_data_58 : _GEN_2045; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2047 = 14'h3b == parameter_2_25 ? phv_data_59 : _GEN_2046; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2048 = 14'h3c == parameter_2_25 ? phv_data_60 : _GEN_2047; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2049 = 14'h3d == parameter_2_25 ? phv_data_61 : _GEN_2048; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2050 = 14'h3e == parameter_2_25 ? phv_data_62 : _GEN_2049; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2051 = 14'h3f == parameter_2_25 ? phv_data_63 : _GEN_2050; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_26 = vliw_26[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_26 = vliw_26[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_26 = parameter_2_26[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_26 = parameter_2_26[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_26 = {{1'd0}, args_offset_26}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_26 = _total_offset_T_26[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2055 = 3'h1 == total_offset_26 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2056 = 3'h2 == total_offset_26 ? args_2 : _GEN_2055; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2057 = 3'h3 == total_offset_26 ? args_3 : _GEN_2056; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2058 = 3'h4 == total_offset_26 ? args_4 : _GEN_2057; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2059 = 3'h5 == total_offset_26 ? args_5 : _GEN_2058; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2060 = 3'h6 == total_offset_26 ? args_6 : _GEN_2059; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2061 = total_offset_26 < 3'h7 ? _GEN_2060 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_26_0 = 3'h0 < args_length_26 ? _GEN_2061 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_2063 = opcode_26 == 4'ha ? field_bytes_26_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2064 = opcode_26 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1849 = opcode_26 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_53 = _T_1849 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_2065 = opcode_26 == 4'h8 | opcode_26 == 4'hb ? parameter_2_26[7:0] : _GEN_2063; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_2066 = opcode_26 == 4'h8 | opcode_26 == 4'hb ? _field_tag_T_53 : _GEN_2064; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_2067 = 14'h0 == parameter_2_26 ? phv_data_0 : _GEN_2065; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2068 = 14'h1 == parameter_2_26 ? phv_data_1 : _GEN_2067; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2069 = 14'h2 == parameter_2_26 ? phv_data_2 : _GEN_2068; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2070 = 14'h3 == parameter_2_26 ? phv_data_3 : _GEN_2069; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2071 = 14'h4 == parameter_2_26 ? phv_data_4 : _GEN_2070; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2072 = 14'h5 == parameter_2_26 ? phv_data_5 : _GEN_2071; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2073 = 14'h6 == parameter_2_26 ? phv_data_6 : _GEN_2072; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2074 = 14'h7 == parameter_2_26 ? phv_data_7 : _GEN_2073; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2075 = 14'h8 == parameter_2_26 ? phv_data_8 : _GEN_2074; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2076 = 14'h9 == parameter_2_26 ? phv_data_9 : _GEN_2075; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2077 = 14'ha == parameter_2_26 ? phv_data_10 : _GEN_2076; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2078 = 14'hb == parameter_2_26 ? phv_data_11 : _GEN_2077; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2079 = 14'hc == parameter_2_26 ? phv_data_12 : _GEN_2078; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2080 = 14'hd == parameter_2_26 ? phv_data_13 : _GEN_2079; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2081 = 14'he == parameter_2_26 ? phv_data_14 : _GEN_2080; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2082 = 14'hf == parameter_2_26 ? phv_data_15 : _GEN_2081; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2083 = 14'h10 == parameter_2_26 ? phv_data_16 : _GEN_2082; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2084 = 14'h11 == parameter_2_26 ? phv_data_17 : _GEN_2083; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2085 = 14'h12 == parameter_2_26 ? phv_data_18 : _GEN_2084; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2086 = 14'h13 == parameter_2_26 ? phv_data_19 : _GEN_2085; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2087 = 14'h14 == parameter_2_26 ? phv_data_20 : _GEN_2086; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2088 = 14'h15 == parameter_2_26 ? phv_data_21 : _GEN_2087; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2089 = 14'h16 == parameter_2_26 ? phv_data_22 : _GEN_2088; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2090 = 14'h17 == parameter_2_26 ? phv_data_23 : _GEN_2089; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2091 = 14'h18 == parameter_2_26 ? phv_data_24 : _GEN_2090; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2092 = 14'h19 == parameter_2_26 ? phv_data_25 : _GEN_2091; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2093 = 14'h1a == parameter_2_26 ? phv_data_26 : _GEN_2092; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2094 = 14'h1b == parameter_2_26 ? phv_data_27 : _GEN_2093; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2095 = 14'h1c == parameter_2_26 ? phv_data_28 : _GEN_2094; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2096 = 14'h1d == parameter_2_26 ? phv_data_29 : _GEN_2095; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2097 = 14'h1e == parameter_2_26 ? phv_data_30 : _GEN_2096; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2098 = 14'h1f == parameter_2_26 ? phv_data_31 : _GEN_2097; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2099 = 14'h20 == parameter_2_26 ? phv_data_32 : _GEN_2098; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2100 = 14'h21 == parameter_2_26 ? phv_data_33 : _GEN_2099; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2101 = 14'h22 == parameter_2_26 ? phv_data_34 : _GEN_2100; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2102 = 14'h23 == parameter_2_26 ? phv_data_35 : _GEN_2101; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2103 = 14'h24 == parameter_2_26 ? phv_data_36 : _GEN_2102; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2104 = 14'h25 == parameter_2_26 ? phv_data_37 : _GEN_2103; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2105 = 14'h26 == parameter_2_26 ? phv_data_38 : _GEN_2104; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2106 = 14'h27 == parameter_2_26 ? phv_data_39 : _GEN_2105; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2107 = 14'h28 == parameter_2_26 ? phv_data_40 : _GEN_2106; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2108 = 14'h29 == parameter_2_26 ? phv_data_41 : _GEN_2107; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2109 = 14'h2a == parameter_2_26 ? phv_data_42 : _GEN_2108; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2110 = 14'h2b == parameter_2_26 ? phv_data_43 : _GEN_2109; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2111 = 14'h2c == parameter_2_26 ? phv_data_44 : _GEN_2110; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2112 = 14'h2d == parameter_2_26 ? phv_data_45 : _GEN_2111; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2113 = 14'h2e == parameter_2_26 ? phv_data_46 : _GEN_2112; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2114 = 14'h2f == parameter_2_26 ? phv_data_47 : _GEN_2113; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2115 = 14'h30 == parameter_2_26 ? phv_data_48 : _GEN_2114; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2116 = 14'h31 == parameter_2_26 ? phv_data_49 : _GEN_2115; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2117 = 14'h32 == parameter_2_26 ? phv_data_50 : _GEN_2116; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2118 = 14'h33 == parameter_2_26 ? phv_data_51 : _GEN_2117; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2119 = 14'h34 == parameter_2_26 ? phv_data_52 : _GEN_2118; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2120 = 14'h35 == parameter_2_26 ? phv_data_53 : _GEN_2119; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2121 = 14'h36 == parameter_2_26 ? phv_data_54 : _GEN_2120; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2122 = 14'h37 == parameter_2_26 ? phv_data_55 : _GEN_2121; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2123 = 14'h38 == parameter_2_26 ? phv_data_56 : _GEN_2122; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2124 = 14'h39 == parameter_2_26 ? phv_data_57 : _GEN_2123; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2125 = 14'h3a == parameter_2_26 ? phv_data_58 : _GEN_2124; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2126 = 14'h3b == parameter_2_26 ? phv_data_59 : _GEN_2125; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2127 = 14'h3c == parameter_2_26 ? phv_data_60 : _GEN_2126; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2128 = 14'h3d == parameter_2_26 ? phv_data_61 : _GEN_2127; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2129 = 14'h3e == parameter_2_26 ? phv_data_62 : _GEN_2128; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2130 = 14'h3f == parameter_2_26 ? phv_data_63 : _GEN_2129; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_27 = vliw_27[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_27 = vliw_27[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_27 = parameter_2_27[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_27 = parameter_2_27[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_27 = {{1'd0}, args_offset_27}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_27 = _total_offset_T_27[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2134 = 3'h1 == total_offset_27 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2135 = 3'h2 == total_offset_27 ? args_2 : _GEN_2134; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2136 = 3'h3 == total_offset_27 ? args_3 : _GEN_2135; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2137 = 3'h4 == total_offset_27 ? args_4 : _GEN_2136; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2138 = 3'h5 == total_offset_27 ? args_5 : _GEN_2137; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2139 = 3'h6 == total_offset_27 ? args_6 : _GEN_2138; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2140 = total_offset_27 < 3'h7 ? _GEN_2139 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_27_0 = 3'h0 < args_length_27 ? _GEN_2140 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_2142 = opcode_27 == 4'ha ? field_bytes_27_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2143 = opcode_27 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1920 = opcode_27 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_55 = _T_1920 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_2144 = opcode_27 == 4'h8 | opcode_27 == 4'hb ? parameter_2_27[7:0] : _GEN_2142; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_2145 = opcode_27 == 4'h8 | opcode_27 == 4'hb ? _field_tag_T_55 : _GEN_2143; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_2146 = 14'h0 == parameter_2_27 ? phv_data_0 : _GEN_2144; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2147 = 14'h1 == parameter_2_27 ? phv_data_1 : _GEN_2146; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2148 = 14'h2 == parameter_2_27 ? phv_data_2 : _GEN_2147; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2149 = 14'h3 == parameter_2_27 ? phv_data_3 : _GEN_2148; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2150 = 14'h4 == parameter_2_27 ? phv_data_4 : _GEN_2149; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2151 = 14'h5 == parameter_2_27 ? phv_data_5 : _GEN_2150; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2152 = 14'h6 == parameter_2_27 ? phv_data_6 : _GEN_2151; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2153 = 14'h7 == parameter_2_27 ? phv_data_7 : _GEN_2152; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2154 = 14'h8 == parameter_2_27 ? phv_data_8 : _GEN_2153; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2155 = 14'h9 == parameter_2_27 ? phv_data_9 : _GEN_2154; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2156 = 14'ha == parameter_2_27 ? phv_data_10 : _GEN_2155; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2157 = 14'hb == parameter_2_27 ? phv_data_11 : _GEN_2156; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2158 = 14'hc == parameter_2_27 ? phv_data_12 : _GEN_2157; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2159 = 14'hd == parameter_2_27 ? phv_data_13 : _GEN_2158; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2160 = 14'he == parameter_2_27 ? phv_data_14 : _GEN_2159; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2161 = 14'hf == parameter_2_27 ? phv_data_15 : _GEN_2160; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2162 = 14'h10 == parameter_2_27 ? phv_data_16 : _GEN_2161; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2163 = 14'h11 == parameter_2_27 ? phv_data_17 : _GEN_2162; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2164 = 14'h12 == parameter_2_27 ? phv_data_18 : _GEN_2163; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2165 = 14'h13 == parameter_2_27 ? phv_data_19 : _GEN_2164; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2166 = 14'h14 == parameter_2_27 ? phv_data_20 : _GEN_2165; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2167 = 14'h15 == parameter_2_27 ? phv_data_21 : _GEN_2166; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2168 = 14'h16 == parameter_2_27 ? phv_data_22 : _GEN_2167; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2169 = 14'h17 == parameter_2_27 ? phv_data_23 : _GEN_2168; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2170 = 14'h18 == parameter_2_27 ? phv_data_24 : _GEN_2169; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2171 = 14'h19 == parameter_2_27 ? phv_data_25 : _GEN_2170; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2172 = 14'h1a == parameter_2_27 ? phv_data_26 : _GEN_2171; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2173 = 14'h1b == parameter_2_27 ? phv_data_27 : _GEN_2172; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2174 = 14'h1c == parameter_2_27 ? phv_data_28 : _GEN_2173; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2175 = 14'h1d == parameter_2_27 ? phv_data_29 : _GEN_2174; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2176 = 14'h1e == parameter_2_27 ? phv_data_30 : _GEN_2175; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2177 = 14'h1f == parameter_2_27 ? phv_data_31 : _GEN_2176; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2178 = 14'h20 == parameter_2_27 ? phv_data_32 : _GEN_2177; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2179 = 14'h21 == parameter_2_27 ? phv_data_33 : _GEN_2178; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2180 = 14'h22 == parameter_2_27 ? phv_data_34 : _GEN_2179; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2181 = 14'h23 == parameter_2_27 ? phv_data_35 : _GEN_2180; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2182 = 14'h24 == parameter_2_27 ? phv_data_36 : _GEN_2181; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2183 = 14'h25 == parameter_2_27 ? phv_data_37 : _GEN_2182; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2184 = 14'h26 == parameter_2_27 ? phv_data_38 : _GEN_2183; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2185 = 14'h27 == parameter_2_27 ? phv_data_39 : _GEN_2184; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2186 = 14'h28 == parameter_2_27 ? phv_data_40 : _GEN_2185; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2187 = 14'h29 == parameter_2_27 ? phv_data_41 : _GEN_2186; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2188 = 14'h2a == parameter_2_27 ? phv_data_42 : _GEN_2187; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2189 = 14'h2b == parameter_2_27 ? phv_data_43 : _GEN_2188; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2190 = 14'h2c == parameter_2_27 ? phv_data_44 : _GEN_2189; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2191 = 14'h2d == parameter_2_27 ? phv_data_45 : _GEN_2190; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2192 = 14'h2e == parameter_2_27 ? phv_data_46 : _GEN_2191; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2193 = 14'h2f == parameter_2_27 ? phv_data_47 : _GEN_2192; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2194 = 14'h30 == parameter_2_27 ? phv_data_48 : _GEN_2193; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2195 = 14'h31 == parameter_2_27 ? phv_data_49 : _GEN_2194; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2196 = 14'h32 == parameter_2_27 ? phv_data_50 : _GEN_2195; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2197 = 14'h33 == parameter_2_27 ? phv_data_51 : _GEN_2196; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2198 = 14'h34 == parameter_2_27 ? phv_data_52 : _GEN_2197; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2199 = 14'h35 == parameter_2_27 ? phv_data_53 : _GEN_2198; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2200 = 14'h36 == parameter_2_27 ? phv_data_54 : _GEN_2199; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2201 = 14'h37 == parameter_2_27 ? phv_data_55 : _GEN_2200; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2202 = 14'h38 == parameter_2_27 ? phv_data_56 : _GEN_2201; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2203 = 14'h39 == parameter_2_27 ? phv_data_57 : _GEN_2202; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2204 = 14'h3a == parameter_2_27 ? phv_data_58 : _GEN_2203; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2205 = 14'h3b == parameter_2_27 ? phv_data_59 : _GEN_2204; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2206 = 14'h3c == parameter_2_27 ? phv_data_60 : _GEN_2205; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2207 = 14'h3d == parameter_2_27 ? phv_data_61 : _GEN_2206; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2208 = 14'h3e == parameter_2_27 ? phv_data_62 : _GEN_2207; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2209 = 14'h3f == parameter_2_27 ? phv_data_63 : _GEN_2208; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_28 = vliw_28[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_28 = vliw_28[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_28 = parameter_2_28[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_28 = parameter_2_28[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_28 = {{1'd0}, args_offset_28}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_28 = _total_offset_T_28[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2213 = 3'h1 == total_offset_28 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2214 = 3'h2 == total_offset_28 ? args_2 : _GEN_2213; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2215 = 3'h3 == total_offset_28 ? args_3 : _GEN_2214; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2216 = 3'h4 == total_offset_28 ? args_4 : _GEN_2215; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2217 = 3'h5 == total_offset_28 ? args_5 : _GEN_2216; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2218 = 3'h6 == total_offset_28 ? args_6 : _GEN_2217; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2219 = total_offset_28 < 3'h7 ? _GEN_2218 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_28_0 = 3'h0 < args_length_28 ? _GEN_2219 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_2221 = opcode_28 == 4'ha ? field_bytes_28_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2222 = opcode_28 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1991 = opcode_28 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_57 = _T_1991 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_2223 = opcode_28 == 4'h8 | opcode_28 == 4'hb ? parameter_2_28[7:0] : _GEN_2221; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_2224 = opcode_28 == 4'h8 | opcode_28 == 4'hb ? _field_tag_T_57 : _GEN_2222; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_2225 = 14'h0 == parameter_2_28 ? phv_data_0 : _GEN_2223; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2226 = 14'h1 == parameter_2_28 ? phv_data_1 : _GEN_2225; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2227 = 14'h2 == parameter_2_28 ? phv_data_2 : _GEN_2226; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2228 = 14'h3 == parameter_2_28 ? phv_data_3 : _GEN_2227; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2229 = 14'h4 == parameter_2_28 ? phv_data_4 : _GEN_2228; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2230 = 14'h5 == parameter_2_28 ? phv_data_5 : _GEN_2229; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2231 = 14'h6 == parameter_2_28 ? phv_data_6 : _GEN_2230; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2232 = 14'h7 == parameter_2_28 ? phv_data_7 : _GEN_2231; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2233 = 14'h8 == parameter_2_28 ? phv_data_8 : _GEN_2232; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2234 = 14'h9 == parameter_2_28 ? phv_data_9 : _GEN_2233; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2235 = 14'ha == parameter_2_28 ? phv_data_10 : _GEN_2234; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2236 = 14'hb == parameter_2_28 ? phv_data_11 : _GEN_2235; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2237 = 14'hc == parameter_2_28 ? phv_data_12 : _GEN_2236; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2238 = 14'hd == parameter_2_28 ? phv_data_13 : _GEN_2237; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2239 = 14'he == parameter_2_28 ? phv_data_14 : _GEN_2238; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2240 = 14'hf == parameter_2_28 ? phv_data_15 : _GEN_2239; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2241 = 14'h10 == parameter_2_28 ? phv_data_16 : _GEN_2240; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2242 = 14'h11 == parameter_2_28 ? phv_data_17 : _GEN_2241; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2243 = 14'h12 == parameter_2_28 ? phv_data_18 : _GEN_2242; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2244 = 14'h13 == parameter_2_28 ? phv_data_19 : _GEN_2243; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2245 = 14'h14 == parameter_2_28 ? phv_data_20 : _GEN_2244; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2246 = 14'h15 == parameter_2_28 ? phv_data_21 : _GEN_2245; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2247 = 14'h16 == parameter_2_28 ? phv_data_22 : _GEN_2246; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2248 = 14'h17 == parameter_2_28 ? phv_data_23 : _GEN_2247; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2249 = 14'h18 == parameter_2_28 ? phv_data_24 : _GEN_2248; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2250 = 14'h19 == parameter_2_28 ? phv_data_25 : _GEN_2249; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2251 = 14'h1a == parameter_2_28 ? phv_data_26 : _GEN_2250; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2252 = 14'h1b == parameter_2_28 ? phv_data_27 : _GEN_2251; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2253 = 14'h1c == parameter_2_28 ? phv_data_28 : _GEN_2252; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2254 = 14'h1d == parameter_2_28 ? phv_data_29 : _GEN_2253; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2255 = 14'h1e == parameter_2_28 ? phv_data_30 : _GEN_2254; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2256 = 14'h1f == parameter_2_28 ? phv_data_31 : _GEN_2255; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2257 = 14'h20 == parameter_2_28 ? phv_data_32 : _GEN_2256; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2258 = 14'h21 == parameter_2_28 ? phv_data_33 : _GEN_2257; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2259 = 14'h22 == parameter_2_28 ? phv_data_34 : _GEN_2258; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2260 = 14'h23 == parameter_2_28 ? phv_data_35 : _GEN_2259; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2261 = 14'h24 == parameter_2_28 ? phv_data_36 : _GEN_2260; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2262 = 14'h25 == parameter_2_28 ? phv_data_37 : _GEN_2261; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2263 = 14'h26 == parameter_2_28 ? phv_data_38 : _GEN_2262; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2264 = 14'h27 == parameter_2_28 ? phv_data_39 : _GEN_2263; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2265 = 14'h28 == parameter_2_28 ? phv_data_40 : _GEN_2264; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2266 = 14'h29 == parameter_2_28 ? phv_data_41 : _GEN_2265; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2267 = 14'h2a == parameter_2_28 ? phv_data_42 : _GEN_2266; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2268 = 14'h2b == parameter_2_28 ? phv_data_43 : _GEN_2267; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2269 = 14'h2c == parameter_2_28 ? phv_data_44 : _GEN_2268; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2270 = 14'h2d == parameter_2_28 ? phv_data_45 : _GEN_2269; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2271 = 14'h2e == parameter_2_28 ? phv_data_46 : _GEN_2270; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2272 = 14'h2f == parameter_2_28 ? phv_data_47 : _GEN_2271; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2273 = 14'h30 == parameter_2_28 ? phv_data_48 : _GEN_2272; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2274 = 14'h31 == parameter_2_28 ? phv_data_49 : _GEN_2273; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2275 = 14'h32 == parameter_2_28 ? phv_data_50 : _GEN_2274; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2276 = 14'h33 == parameter_2_28 ? phv_data_51 : _GEN_2275; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2277 = 14'h34 == parameter_2_28 ? phv_data_52 : _GEN_2276; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2278 = 14'h35 == parameter_2_28 ? phv_data_53 : _GEN_2277; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2279 = 14'h36 == parameter_2_28 ? phv_data_54 : _GEN_2278; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2280 = 14'h37 == parameter_2_28 ? phv_data_55 : _GEN_2279; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2281 = 14'h38 == parameter_2_28 ? phv_data_56 : _GEN_2280; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2282 = 14'h39 == parameter_2_28 ? phv_data_57 : _GEN_2281; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2283 = 14'h3a == parameter_2_28 ? phv_data_58 : _GEN_2282; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2284 = 14'h3b == parameter_2_28 ? phv_data_59 : _GEN_2283; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2285 = 14'h3c == parameter_2_28 ? phv_data_60 : _GEN_2284; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2286 = 14'h3d == parameter_2_28 ? phv_data_61 : _GEN_2285; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2287 = 14'h3e == parameter_2_28 ? phv_data_62 : _GEN_2286; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2288 = 14'h3f == parameter_2_28 ? phv_data_63 : _GEN_2287; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_29 = vliw_29[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_29 = vliw_29[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_29 = parameter_2_29[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_29 = parameter_2_29[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_29 = {{1'd0}, args_offset_29}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_29 = _total_offset_T_29[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2292 = 3'h1 == total_offset_29 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2293 = 3'h2 == total_offset_29 ? args_2 : _GEN_2292; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2294 = 3'h3 == total_offset_29 ? args_3 : _GEN_2293; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2295 = 3'h4 == total_offset_29 ? args_4 : _GEN_2294; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2296 = 3'h5 == total_offset_29 ? args_5 : _GEN_2295; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2297 = 3'h6 == total_offset_29 ? args_6 : _GEN_2296; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2298 = total_offset_29 < 3'h7 ? _GEN_2297 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_29_0 = 3'h0 < args_length_29 ? _GEN_2298 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_2300 = opcode_29 == 4'ha ? field_bytes_29_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2301 = opcode_29 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2062 = opcode_29 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_59 = _T_2062 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_2302 = opcode_29 == 4'h8 | opcode_29 == 4'hb ? parameter_2_29[7:0] : _GEN_2300; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_2303 = opcode_29 == 4'h8 | opcode_29 == 4'hb ? _field_tag_T_59 : _GEN_2301; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_2304 = 14'h0 == parameter_2_29 ? phv_data_0 : _GEN_2302; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2305 = 14'h1 == parameter_2_29 ? phv_data_1 : _GEN_2304; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2306 = 14'h2 == parameter_2_29 ? phv_data_2 : _GEN_2305; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2307 = 14'h3 == parameter_2_29 ? phv_data_3 : _GEN_2306; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2308 = 14'h4 == parameter_2_29 ? phv_data_4 : _GEN_2307; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2309 = 14'h5 == parameter_2_29 ? phv_data_5 : _GEN_2308; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2310 = 14'h6 == parameter_2_29 ? phv_data_6 : _GEN_2309; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2311 = 14'h7 == parameter_2_29 ? phv_data_7 : _GEN_2310; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2312 = 14'h8 == parameter_2_29 ? phv_data_8 : _GEN_2311; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2313 = 14'h9 == parameter_2_29 ? phv_data_9 : _GEN_2312; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2314 = 14'ha == parameter_2_29 ? phv_data_10 : _GEN_2313; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2315 = 14'hb == parameter_2_29 ? phv_data_11 : _GEN_2314; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2316 = 14'hc == parameter_2_29 ? phv_data_12 : _GEN_2315; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2317 = 14'hd == parameter_2_29 ? phv_data_13 : _GEN_2316; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2318 = 14'he == parameter_2_29 ? phv_data_14 : _GEN_2317; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2319 = 14'hf == parameter_2_29 ? phv_data_15 : _GEN_2318; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2320 = 14'h10 == parameter_2_29 ? phv_data_16 : _GEN_2319; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2321 = 14'h11 == parameter_2_29 ? phv_data_17 : _GEN_2320; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2322 = 14'h12 == parameter_2_29 ? phv_data_18 : _GEN_2321; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2323 = 14'h13 == parameter_2_29 ? phv_data_19 : _GEN_2322; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2324 = 14'h14 == parameter_2_29 ? phv_data_20 : _GEN_2323; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2325 = 14'h15 == parameter_2_29 ? phv_data_21 : _GEN_2324; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2326 = 14'h16 == parameter_2_29 ? phv_data_22 : _GEN_2325; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2327 = 14'h17 == parameter_2_29 ? phv_data_23 : _GEN_2326; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2328 = 14'h18 == parameter_2_29 ? phv_data_24 : _GEN_2327; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2329 = 14'h19 == parameter_2_29 ? phv_data_25 : _GEN_2328; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2330 = 14'h1a == parameter_2_29 ? phv_data_26 : _GEN_2329; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2331 = 14'h1b == parameter_2_29 ? phv_data_27 : _GEN_2330; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2332 = 14'h1c == parameter_2_29 ? phv_data_28 : _GEN_2331; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2333 = 14'h1d == parameter_2_29 ? phv_data_29 : _GEN_2332; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2334 = 14'h1e == parameter_2_29 ? phv_data_30 : _GEN_2333; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2335 = 14'h1f == parameter_2_29 ? phv_data_31 : _GEN_2334; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2336 = 14'h20 == parameter_2_29 ? phv_data_32 : _GEN_2335; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2337 = 14'h21 == parameter_2_29 ? phv_data_33 : _GEN_2336; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2338 = 14'h22 == parameter_2_29 ? phv_data_34 : _GEN_2337; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2339 = 14'h23 == parameter_2_29 ? phv_data_35 : _GEN_2338; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2340 = 14'h24 == parameter_2_29 ? phv_data_36 : _GEN_2339; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2341 = 14'h25 == parameter_2_29 ? phv_data_37 : _GEN_2340; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2342 = 14'h26 == parameter_2_29 ? phv_data_38 : _GEN_2341; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2343 = 14'h27 == parameter_2_29 ? phv_data_39 : _GEN_2342; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2344 = 14'h28 == parameter_2_29 ? phv_data_40 : _GEN_2343; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2345 = 14'h29 == parameter_2_29 ? phv_data_41 : _GEN_2344; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2346 = 14'h2a == parameter_2_29 ? phv_data_42 : _GEN_2345; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2347 = 14'h2b == parameter_2_29 ? phv_data_43 : _GEN_2346; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2348 = 14'h2c == parameter_2_29 ? phv_data_44 : _GEN_2347; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2349 = 14'h2d == parameter_2_29 ? phv_data_45 : _GEN_2348; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2350 = 14'h2e == parameter_2_29 ? phv_data_46 : _GEN_2349; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2351 = 14'h2f == parameter_2_29 ? phv_data_47 : _GEN_2350; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2352 = 14'h30 == parameter_2_29 ? phv_data_48 : _GEN_2351; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2353 = 14'h31 == parameter_2_29 ? phv_data_49 : _GEN_2352; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2354 = 14'h32 == parameter_2_29 ? phv_data_50 : _GEN_2353; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2355 = 14'h33 == parameter_2_29 ? phv_data_51 : _GEN_2354; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2356 = 14'h34 == parameter_2_29 ? phv_data_52 : _GEN_2355; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2357 = 14'h35 == parameter_2_29 ? phv_data_53 : _GEN_2356; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2358 = 14'h36 == parameter_2_29 ? phv_data_54 : _GEN_2357; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2359 = 14'h37 == parameter_2_29 ? phv_data_55 : _GEN_2358; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2360 = 14'h38 == parameter_2_29 ? phv_data_56 : _GEN_2359; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2361 = 14'h39 == parameter_2_29 ? phv_data_57 : _GEN_2360; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2362 = 14'h3a == parameter_2_29 ? phv_data_58 : _GEN_2361; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2363 = 14'h3b == parameter_2_29 ? phv_data_59 : _GEN_2362; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2364 = 14'h3c == parameter_2_29 ? phv_data_60 : _GEN_2363; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2365 = 14'h3d == parameter_2_29 ? phv_data_61 : _GEN_2364; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2366 = 14'h3e == parameter_2_29 ? phv_data_62 : _GEN_2365; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2367 = 14'h3f == parameter_2_29 ? phv_data_63 : _GEN_2366; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_30 = vliw_30[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_30 = vliw_30[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_30 = parameter_2_30[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_30 = parameter_2_30[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_30 = {{1'd0}, args_offset_30}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_30 = _total_offset_T_30[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2371 = 3'h1 == total_offset_30 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2372 = 3'h2 == total_offset_30 ? args_2 : _GEN_2371; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2373 = 3'h3 == total_offset_30 ? args_3 : _GEN_2372; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2374 = 3'h4 == total_offset_30 ? args_4 : _GEN_2373; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2375 = 3'h5 == total_offset_30 ? args_5 : _GEN_2374; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2376 = 3'h6 == total_offset_30 ? args_6 : _GEN_2375; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2377 = total_offset_30 < 3'h7 ? _GEN_2376 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_30_0 = 3'h0 < args_length_30 ? _GEN_2377 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_2379 = opcode_30 == 4'ha ? field_bytes_30_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2380 = opcode_30 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2133 = opcode_30 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_61 = _T_2133 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_2381 = opcode_30 == 4'h8 | opcode_30 == 4'hb ? parameter_2_30[7:0] : _GEN_2379; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_2382 = opcode_30 == 4'h8 | opcode_30 == 4'hb ? _field_tag_T_61 : _GEN_2380; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_2383 = 14'h0 == parameter_2_30 ? phv_data_0 : _GEN_2381; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2384 = 14'h1 == parameter_2_30 ? phv_data_1 : _GEN_2383; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2385 = 14'h2 == parameter_2_30 ? phv_data_2 : _GEN_2384; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2386 = 14'h3 == parameter_2_30 ? phv_data_3 : _GEN_2385; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2387 = 14'h4 == parameter_2_30 ? phv_data_4 : _GEN_2386; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2388 = 14'h5 == parameter_2_30 ? phv_data_5 : _GEN_2387; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2389 = 14'h6 == parameter_2_30 ? phv_data_6 : _GEN_2388; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2390 = 14'h7 == parameter_2_30 ? phv_data_7 : _GEN_2389; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2391 = 14'h8 == parameter_2_30 ? phv_data_8 : _GEN_2390; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2392 = 14'h9 == parameter_2_30 ? phv_data_9 : _GEN_2391; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2393 = 14'ha == parameter_2_30 ? phv_data_10 : _GEN_2392; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2394 = 14'hb == parameter_2_30 ? phv_data_11 : _GEN_2393; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2395 = 14'hc == parameter_2_30 ? phv_data_12 : _GEN_2394; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2396 = 14'hd == parameter_2_30 ? phv_data_13 : _GEN_2395; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2397 = 14'he == parameter_2_30 ? phv_data_14 : _GEN_2396; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2398 = 14'hf == parameter_2_30 ? phv_data_15 : _GEN_2397; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2399 = 14'h10 == parameter_2_30 ? phv_data_16 : _GEN_2398; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2400 = 14'h11 == parameter_2_30 ? phv_data_17 : _GEN_2399; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2401 = 14'h12 == parameter_2_30 ? phv_data_18 : _GEN_2400; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2402 = 14'h13 == parameter_2_30 ? phv_data_19 : _GEN_2401; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2403 = 14'h14 == parameter_2_30 ? phv_data_20 : _GEN_2402; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2404 = 14'h15 == parameter_2_30 ? phv_data_21 : _GEN_2403; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2405 = 14'h16 == parameter_2_30 ? phv_data_22 : _GEN_2404; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2406 = 14'h17 == parameter_2_30 ? phv_data_23 : _GEN_2405; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2407 = 14'h18 == parameter_2_30 ? phv_data_24 : _GEN_2406; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2408 = 14'h19 == parameter_2_30 ? phv_data_25 : _GEN_2407; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2409 = 14'h1a == parameter_2_30 ? phv_data_26 : _GEN_2408; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2410 = 14'h1b == parameter_2_30 ? phv_data_27 : _GEN_2409; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2411 = 14'h1c == parameter_2_30 ? phv_data_28 : _GEN_2410; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2412 = 14'h1d == parameter_2_30 ? phv_data_29 : _GEN_2411; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2413 = 14'h1e == parameter_2_30 ? phv_data_30 : _GEN_2412; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2414 = 14'h1f == parameter_2_30 ? phv_data_31 : _GEN_2413; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2415 = 14'h20 == parameter_2_30 ? phv_data_32 : _GEN_2414; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2416 = 14'h21 == parameter_2_30 ? phv_data_33 : _GEN_2415; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2417 = 14'h22 == parameter_2_30 ? phv_data_34 : _GEN_2416; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2418 = 14'h23 == parameter_2_30 ? phv_data_35 : _GEN_2417; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2419 = 14'h24 == parameter_2_30 ? phv_data_36 : _GEN_2418; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2420 = 14'h25 == parameter_2_30 ? phv_data_37 : _GEN_2419; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2421 = 14'h26 == parameter_2_30 ? phv_data_38 : _GEN_2420; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2422 = 14'h27 == parameter_2_30 ? phv_data_39 : _GEN_2421; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2423 = 14'h28 == parameter_2_30 ? phv_data_40 : _GEN_2422; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2424 = 14'h29 == parameter_2_30 ? phv_data_41 : _GEN_2423; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2425 = 14'h2a == parameter_2_30 ? phv_data_42 : _GEN_2424; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2426 = 14'h2b == parameter_2_30 ? phv_data_43 : _GEN_2425; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2427 = 14'h2c == parameter_2_30 ? phv_data_44 : _GEN_2426; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2428 = 14'h2d == parameter_2_30 ? phv_data_45 : _GEN_2427; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2429 = 14'h2e == parameter_2_30 ? phv_data_46 : _GEN_2428; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2430 = 14'h2f == parameter_2_30 ? phv_data_47 : _GEN_2429; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2431 = 14'h30 == parameter_2_30 ? phv_data_48 : _GEN_2430; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2432 = 14'h31 == parameter_2_30 ? phv_data_49 : _GEN_2431; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2433 = 14'h32 == parameter_2_30 ? phv_data_50 : _GEN_2432; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2434 = 14'h33 == parameter_2_30 ? phv_data_51 : _GEN_2433; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2435 = 14'h34 == parameter_2_30 ? phv_data_52 : _GEN_2434; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2436 = 14'h35 == parameter_2_30 ? phv_data_53 : _GEN_2435; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2437 = 14'h36 == parameter_2_30 ? phv_data_54 : _GEN_2436; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2438 = 14'h37 == parameter_2_30 ? phv_data_55 : _GEN_2437; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2439 = 14'h38 == parameter_2_30 ? phv_data_56 : _GEN_2438; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2440 = 14'h39 == parameter_2_30 ? phv_data_57 : _GEN_2439; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2441 = 14'h3a == parameter_2_30 ? phv_data_58 : _GEN_2440; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2442 = 14'h3b == parameter_2_30 ? phv_data_59 : _GEN_2441; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2443 = 14'h3c == parameter_2_30 ? phv_data_60 : _GEN_2442; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2444 = 14'h3d == parameter_2_30 ? phv_data_61 : _GEN_2443; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2445 = 14'h3e == parameter_2_30 ? phv_data_62 : _GEN_2444; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2446 = 14'h3f == parameter_2_30 ? phv_data_63 : _GEN_2445; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_31 = vliw_31[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_31 = vliw_31[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_31 = parameter_2_31[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_31 = parameter_2_31[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_31 = {{1'd0}, args_offset_31}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_31 = _total_offset_T_31[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2450 = 3'h1 == total_offset_31 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2451 = 3'h2 == total_offset_31 ? args_2 : _GEN_2450; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2452 = 3'h3 == total_offset_31 ? args_3 : _GEN_2451; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2453 = 3'h4 == total_offset_31 ? args_4 : _GEN_2452; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2454 = 3'h5 == total_offset_31 ? args_5 : _GEN_2453; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2455 = 3'h6 == total_offset_31 ? args_6 : _GEN_2454; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2456 = total_offset_31 < 3'h7 ? _GEN_2455 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_31_0 = 3'h0 < args_length_31 ? _GEN_2456 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_2458 = opcode_31 == 4'ha ? field_bytes_31_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2459 = opcode_31 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2204 = opcode_31 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_63 = _T_2204 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_2460 = opcode_31 == 4'h8 | opcode_31 == 4'hb ? parameter_2_31[7:0] : _GEN_2458; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_2461 = opcode_31 == 4'h8 | opcode_31 == 4'hb ? _field_tag_T_63 : _GEN_2459; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_2462 = 14'h0 == parameter_2_31 ? phv_data_0 : _GEN_2460; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2463 = 14'h1 == parameter_2_31 ? phv_data_1 : _GEN_2462; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2464 = 14'h2 == parameter_2_31 ? phv_data_2 : _GEN_2463; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2465 = 14'h3 == parameter_2_31 ? phv_data_3 : _GEN_2464; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2466 = 14'h4 == parameter_2_31 ? phv_data_4 : _GEN_2465; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2467 = 14'h5 == parameter_2_31 ? phv_data_5 : _GEN_2466; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2468 = 14'h6 == parameter_2_31 ? phv_data_6 : _GEN_2467; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2469 = 14'h7 == parameter_2_31 ? phv_data_7 : _GEN_2468; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2470 = 14'h8 == parameter_2_31 ? phv_data_8 : _GEN_2469; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2471 = 14'h9 == parameter_2_31 ? phv_data_9 : _GEN_2470; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2472 = 14'ha == parameter_2_31 ? phv_data_10 : _GEN_2471; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2473 = 14'hb == parameter_2_31 ? phv_data_11 : _GEN_2472; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2474 = 14'hc == parameter_2_31 ? phv_data_12 : _GEN_2473; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2475 = 14'hd == parameter_2_31 ? phv_data_13 : _GEN_2474; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2476 = 14'he == parameter_2_31 ? phv_data_14 : _GEN_2475; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2477 = 14'hf == parameter_2_31 ? phv_data_15 : _GEN_2476; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2478 = 14'h10 == parameter_2_31 ? phv_data_16 : _GEN_2477; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2479 = 14'h11 == parameter_2_31 ? phv_data_17 : _GEN_2478; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2480 = 14'h12 == parameter_2_31 ? phv_data_18 : _GEN_2479; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2481 = 14'h13 == parameter_2_31 ? phv_data_19 : _GEN_2480; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2482 = 14'h14 == parameter_2_31 ? phv_data_20 : _GEN_2481; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2483 = 14'h15 == parameter_2_31 ? phv_data_21 : _GEN_2482; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2484 = 14'h16 == parameter_2_31 ? phv_data_22 : _GEN_2483; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2485 = 14'h17 == parameter_2_31 ? phv_data_23 : _GEN_2484; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2486 = 14'h18 == parameter_2_31 ? phv_data_24 : _GEN_2485; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2487 = 14'h19 == parameter_2_31 ? phv_data_25 : _GEN_2486; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2488 = 14'h1a == parameter_2_31 ? phv_data_26 : _GEN_2487; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2489 = 14'h1b == parameter_2_31 ? phv_data_27 : _GEN_2488; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2490 = 14'h1c == parameter_2_31 ? phv_data_28 : _GEN_2489; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2491 = 14'h1d == parameter_2_31 ? phv_data_29 : _GEN_2490; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2492 = 14'h1e == parameter_2_31 ? phv_data_30 : _GEN_2491; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2493 = 14'h1f == parameter_2_31 ? phv_data_31 : _GEN_2492; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2494 = 14'h20 == parameter_2_31 ? phv_data_32 : _GEN_2493; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2495 = 14'h21 == parameter_2_31 ? phv_data_33 : _GEN_2494; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2496 = 14'h22 == parameter_2_31 ? phv_data_34 : _GEN_2495; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2497 = 14'h23 == parameter_2_31 ? phv_data_35 : _GEN_2496; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2498 = 14'h24 == parameter_2_31 ? phv_data_36 : _GEN_2497; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2499 = 14'h25 == parameter_2_31 ? phv_data_37 : _GEN_2498; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2500 = 14'h26 == parameter_2_31 ? phv_data_38 : _GEN_2499; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2501 = 14'h27 == parameter_2_31 ? phv_data_39 : _GEN_2500; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2502 = 14'h28 == parameter_2_31 ? phv_data_40 : _GEN_2501; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2503 = 14'h29 == parameter_2_31 ? phv_data_41 : _GEN_2502; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2504 = 14'h2a == parameter_2_31 ? phv_data_42 : _GEN_2503; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2505 = 14'h2b == parameter_2_31 ? phv_data_43 : _GEN_2504; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2506 = 14'h2c == parameter_2_31 ? phv_data_44 : _GEN_2505; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2507 = 14'h2d == parameter_2_31 ? phv_data_45 : _GEN_2506; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2508 = 14'h2e == parameter_2_31 ? phv_data_46 : _GEN_2507; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2509 = 14'h2f == parameter_2_31 ? phv_data_47 : _GEN_2508; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2510 = 14'h30 == parameter_2_31 ? phv_data_48 : _GEN_2509; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2511 = 14'h31 == parameter_2_31 ? phv_data_49 : _GEN_2510; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2512 = 14'h32 == parameter_2_31 ? phv_data_50 : _GEN_2511; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2513 = 14'h33 == parameter_2_31 ? phv_data_51 : _GEN_2512; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2514 = 14'h34 == parameter_2_31 ? phv_data_52 : _GEN_2513; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2515 = 14'h35 == parameter_2_31 ? phv_data_53 : _GEN_2514; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2516 = 14'h36 == parameter_2_31 ? phv_data_54 : _GEN_2515; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2517 = 14'h37 == parameter_2_31 ? phv_data_55 : _GEN_2516; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2518 = 14'h38 == parameter_2_31 ? phv_data_56 : _GEN_2517; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2519 = 14'h39 == parameter_2_31 ? phv_data_57 : _GEN_2518; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2520 = 14'h3a == parameter_2_31 ? phv_data_58 : _GEN_2519; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2521 = 14'h3b == parameter_2_31 ? phv_data_59 : _GEN_2520; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2522 = 14'h3c == parameter_2_31 ? phv_data_60 : _GEN_2521; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2523 = 14'h3d == parameter_2_31 ? phv_data_61 : _GEN_2522; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2524 = 14'h3e == parameter_2_31 ? phv_data_62 : _GEN_2523; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2525 = 14'h3f == parameter_2_31 ? phv_data_63 : _GEN_2524; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_32 = vliw_32[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_32 = vliw_32[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_32 = parameter_2_32[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_32 = parameter_2_32[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_32 = {{1'd0}, args_offset_32}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_32 = _total_offset_T_32[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2529 = 3'h1 == total_offset_32 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2530 = 3'h2 == total_offset_32 ? args_2 : _GEN_2529; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2531 = 3'h3 == total_offset_32 ? args_3 : _GEN_2530; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2532 = 3'h4 == total_offset_32 ? args_4 : _GEN_2531; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2533 = 3'h5 == total_offset_32 ? args_5 : _GEN_2532; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2534 = 3'h6 == total_offset_32 ? args_6 : _GEN_2533; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2535 = total_offset_32 < 3'h7 ? _GEN_2534 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_32_0 = 3'h0 < args_length_32 ? _GEN_2535 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_2537 = opcode_32 == 4'ha ? field_bytes_32_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2538 = opcode_32 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2275 = opcode_32 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_65 = _T_2275 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_2539 = opcode_32 == 4'h8 | opcode_32 == 4'hb ? parameter_2_32[7:0] : _GEN_2537; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_2540 = opcode_32 == 4'h8 | opcode_32 == 4'hb ? _field_tag_T_65 : _GEN_2538; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_2541 = 14'h0 == parameter_2_32 ? phv_data_0 : _GEN_2539; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2542 = 14'h1 == parameter_2_32 ? phv_data_1 : _GEN_2541; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2543 = 14'h2 == parameter_2_32 ? phv_data_2 : _GEN_2542; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2544 = 14'h3 == parameter_2_32 ? phv_data_3 : _GEN_2543; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2545 = 14'h4 == parameter_2_32 ? phv_data_4 : _GEN_2544; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2546 = 14'h5 == parameter_2_32 ? phv_data_5 : _GEN_2545; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2547 = 14'h6 == parameter_2_32 ? phv_data_6 : _GEN_2546; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2548 = 14'h7 == parameter_2_32 ? phv_data_7 : _GEN_2547; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2549 = 14'h8 == parameter_2_32 ? phv_data_8 : _GEN_2548; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2550 = 14'h9 == parameter_2_32 ? phv_data_9 : _GEN_2549; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2551 = 14'ha == parameter_2_32 ? phv_data_10 : _GEN_2550; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2552 = 14'hb == parameter_2_32 ? phv_data_11 : _GEN_2551; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2553 = 14'hc == parameter_2_32 ? phv_data_12 : _GEN_2552; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2554 = 14'hd == parameter_2_32 ? phv_data_13 : _GEN_2553; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2555 = 14'he == parameter_2_32 ? phv_data_14 : _GEN_2554; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2556 = 14'hf == parameter_2_32 ? phv_data_15 : _GEN_2555; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2557 = 14'h10 == parameter_2_32 ? phv_data_16 : _GEN_2556; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2558 = 14'h11 == parameter_2_32 ? phv_data_17 : _GEN_2557; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2559 = 14'h12 == parameter_2_32 ? phv_data_18 : _GEN_2558; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2560 = 14'h13 == parameter_2_32 ? phv_data_19 : _GEN_2559; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2561 = 14'h14 == parameter_2_32 ? phv_data_20 : _GEN_2560; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2562 = 14'h15 == parameter_2_32 ? phv_data_21 : _GEN_2561; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2563 = 14'h16 == parameter_2_32 ? phv_data_22 : _GEN_2562; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2564 = 14'h17 == parameter_2_32 ? phv_data_23 : _GEN_2563; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2565 = 14'h18 == parameter_2_32 ? phv_data_24 : _GEN_2564; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2566 = 14'h19 == parameter_2_32 ? phv_data_25 : _GEN_2565; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2567 = 14'h1a == parameter_2_32 ? phv_data_26 : _GEN_2566; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2568 = 14'h1b == parameter_2_32 ? phv_data_27 : _GEN_2567; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2569 = 14'h1c == parameter_2_32 ? phv_data_28 : _GEN_2568; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2570 = 14'h1d == parameter_2_32 ? phv_data_29 : _GEN_2569; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2571 = 14'h1e == parameter_2_32 ? phv_data_30 : _GEN_2570; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2572 = 14'h1f == parameter_2_32 ? phv_data_31 : _GEN_2571; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2573 = 14'h20 == parameter_2_32 ? phv_data_32 : _GEN_2572; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2574 = 14'h21 == parameter_2_32 ? phv_data_33 : _GEN_2573; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2575 = 14'h22 == parameter_2_32 ? phv_data_34 : _GEN_2574; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2576 = 14'h23 == parameter_2_32 ? phv_data_35 : _GEN_2575; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2577 = 14'h24 == parameter_2_32 ? phv_data_36 : _GEN_2576; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2578 = 14'h25 == parameter_2_32 ? phv_data_37 : _GEN_2577; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2579 = 14'h26 == parameter_2_32 ? phv_data_38 : _GEN_2578; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2580 = 14'h27 == parameter_2_32 ? phv_data_39 : _GEN_2579; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2581 = 14'h28 == parameter_2_32 ? phv_data_40 : _GEN_2580; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2582 = 14'h29 == parameter_2_32 ? phv_data_41 : _GEN_2581; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2583 = 14'h2a == parameter_2_32 ? phv_data_42 : _GEN_2582; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2584 = 14'h2b == parameter_2_32 ? phv_data_43 : _GEN_2583; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2585 = 14'h2c == parameter_2_32 ? phv_data_44 : _GEN_2584; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2586 = 14'h2d == parameter_2_32 ? phv_data_45 : _GEN_2585; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2587 = 14'h2e == parameter_2_32 ? phv_data_46 : _GEN_2586; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2588 = 14'h2f == parameter_2_32 ? phv_data_47 : _GEN_2587; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2589 = 14'h30 == parameter_2_32 ? phv_data_48 : _GEN_2588; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2590 = 14'h31 == parameter_2_32 ? phv_data_49 : _GEN_2589; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2591 = 14'h32 == parameter_2_32 ? phv_data_50 : _GEN_2590; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2592 = 14'h33 == parameter_2_32 ? phv_data_51 : _GEN_2591; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2593 = 14'h34 == parameter_2_32 ? phv_data_52 : _GEN_2592; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2594 = 14'h35 == parameter_2_32 ? phv_data_53 : _GEN_2593; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2595 = 14'h36 == parameter_2_32 ? phv_data_54 : _GEN_2594; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2596 = 14'h37 == parameter_2_32 ? phv_data_55 : _GEN_2595; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2597 = 14'h38 == parameter_2_32 ? phv_data_56 : _GEN_2596; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2598 = 14'h39 == parameter_2_32 ? phv_data_57 : _GEN_2597; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2599 = 14'h3a == parameter_2_32 ? phv_data_58 : _GEN_2598; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2600 = 14'h3b == parameter_2_32 ? phv_data_59 : _GEN_2599; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2601 = 14'h3c == parameter_2_32 ? phv_data_60 : _GEN_2600; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2602 = 14'h3d == parameter_2_32 ? phv_data_61 : _GEN_2601; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2603 = 14'h3e == parameter_2_32 ? phv_data_62 : _GEN_2602; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2604 = 14'h3f == parameter_2_32 ? phv_data_63 : _GEN_2603; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_33 = vliw_33[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_33 = vliw_33[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_33 = parameter_2_33[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_33 = parameter_2_33[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_33 = {{1'd0}, args_offset_33}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_33 = _total_offset_T_33[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2608 = 3'h1 == total_offset_33 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2609 = 3'h2 == total_offset_33 ? args_2 : _GEN_2608; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2610 = 3'h3 == total_offset_33 ? args_3 : _GEN_2609; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2611 = 3'h4 == total_offset_33 ? args_4 : _GEN_2610; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2612 = 3'h5 == total_offset_33 ? args_5 : _GEN_2611; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2613 = 3'h6 == total_offset_33 ? args_6 : _GEN_2612; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2614 = total_offset_33 < 3'h7 ? _GEN_2613 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_33_0 = 3'h0 < args_length_33 ? _GEN_2614 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_2616 = opcode_33 == 4'ha ? field_bytes_33_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2617 = opcode_33 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2346 = opcode_33 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_67 = _T_2346 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_2618 = opcode_33 == 4'h8 | opcode_33 == 4'hb ? parameter_2_33[7:0] : _GEN_2616; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_2619 = opcode_33 == 4'h8 | opcode_33 == 4'hb ? _field_tag_T_67 : _GEN_2617; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_2620 = 14'h0 == parameter_2_33 ? phv_data_0 : _GEN_2618; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2621 = 14'h1 == parameter_2_33 ? phv_data_1 : _GEN_2620; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2622 = 14'h2 == parameter_2_33 ? phv_data_2 : _GEN_2621; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2623 = 14'h3 == parameter_2_33 ? phv_data_3 : _GEN_2622; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2624 = 14'h4 == parameter_2_33 ? phv_data_4 : _GEN_2623; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2625 = 14'h5 == parameter_2_33 ? phv_data_5 : _GEN_2624; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2626 = 14'h6 == parameter_2_33 ? phv_data_6 : _GEN_2625; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2627 = 14'h7 == parameter_2_33 ? phv_data_7 : _GEN_2626; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2628 = 14'h8 == parameter_2_33 ? phv_data_8 : _GEN_2627; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2629 = 14'h9 == parameter_2_33 ? phv_data_9 : _GEN_2628; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2630 = 14'ha == parameter_2_33 ? phv_data_10 : _GEN_2629; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2631 = 14'hb == parameter_2_33 ? phv_data_11 : _GEN_2630; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2632 = 14'hc == parameter_2_33 ? phv_data_12 : _GEN_2631; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2633 = 14'hd == parameter_2_33 ? phv_data_13 : _GEN_2632; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2634 = 14'he == parameter_2_33 ? phv_data_14 : _GEN_2633; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2635 = 14'hf == parameter_2_33 ? phv_data_15 : _GEN_2634; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2636 = 14'h10 == parameter_2_33 ? phv_data_16 : _GEN_2635; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2637 = 14'h11 == parameter_2_33 ? phv_data_17 : _GEN_2636; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2638 = 14'h12 == parameter_2_33 ? phv_data_18 : _GEN_2637; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2639 = 14'h13 == parameter_2_33 ? phv_data_19 : _GEN_2638; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2640 = 14'h14 == parameter_2_33 ? phv_data_20 : _GEN_2639; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2641 = 14'h15 == parameter_2_33 ? phv_data_21 : _GEN_2640; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2642 = 14'h16 == parameter_2_33 ? phv_data_22 : _GEN_2641; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2643 = 14'h17 == parameter_2_33 ? phv_data_23 : _GEN_2642; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2644 = 14'h18 == parameter_2_33 ? phv_data_24 : _GEN_2643; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2645 = 14'h19 == parameter_2_33 ? phv_data_25 : _GEN_2644; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2646 = 14'h1a == parameter_2_33 ? phv_data_26 : _GEN_2645; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2647 = 14'h1b == parameter_2_33 ? phv_data_27 : _GEN_2646; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2648 = 14'h1c == parameter_2_33 ? phv_data_28 : _GEN_2647; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2649 = 14'h1d == parameter_2_33 ? phv_data_29 : _GEN_2648; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2650 = 14'h1e == parameter_2_33 ? phv_data_30 : _GEN_2649; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2651 = 14'h1f == parameter_2_33 ? phv_data_31 : _GEN_2650; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2652 = 14'h20 == parameter_2_33 ? phv_data_32 : _GEN_2651; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2653 = 14'h21 == parameter_2_33 ? phv_data_33 : _GEN_2652; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2654 = 14'h22 == parameter_2_33 ? phv_data_34 : _GEN_2653; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2655 = 14'h23 == parameter_2_33 ? phv_data_35 : _GEN_2654; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2656 = 14'h24 == parameter_2_33 ? phv_data_36 : _GEN_2655; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2657 = 14'h25 == parameter_2_33 ? phv_data_37 : _GEN_2656; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2658 = 14'h26 == parameter_2_33 ? phv_data_38 : _GEN_2657; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2659 = 14'h27 == parameter_2_33 ? phv_data_39 : _GEN_2658; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2660 = 14'h28 == parameter_2_33 ? phv_data_40 : _GEN_2659; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2661 = 14'h29 == parameter_2_33 ? phv_data_41 : _GEN_2660; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2662 = 14'h2a == parameter_2_33 ? phv_data_42 : _GEN_2661; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2663 = 14'h2b == parameter_2_33 ? phv_data_43 : _GEN_2662; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2664 = 14'h2c == parameter_2_33 ? phv_data_44 : _GEN_2663; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2665 = 14'h2d == parameter_2_33 ? phv_data_45 : _GEN_2664; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2666 = 14'h2e == parameter_2_33 ? phv_data_46 : _GEN_2665; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2667 = 14'h2f == parameter_2_33 ? phv_data_47 : _GEN_2666; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2668 = 14'h30 == parameter_2_33 ? phv_data_48 : _GEN_2667; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2669 = 14'h31 == parameter_2_33 ? phv_data_49 : _GEN_2668; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2670 = 14'h32 == parameter_2_33 ? phv_data_50 : _GEN_2669; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2671 = 14'h33 == parameter_2_33 ? phv_data_51 : _GEN_2670; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2672 = 14'h34 == parameter_2_33 ? phv_data_52 : _GEN_2671; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2673 = 14'h35 == parameter_2_33 ? phv_data_53 : _GEN_2672; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2674 = 14'h36 == parameter_2_33 ? phv_data_54 : _GEN_2673; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2675 = 14'h37 == parameter_2_33 ? phv_data_55 : _GEN_2674; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2676 = 14'h38 == parameter_2_33 ? phv_data_56 : _GEN_2675; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2677 = 14'h39 == parameter_2_33 ? phv_data_57 : _GEN_2676; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2678 = 14'h3a == parameter_2_33 ? phv_data_58 : _GEN_2677; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2679 = 14'h3b == parameter_2_33 ? phv_data_59 : _GEN_2678; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2680 = 14'h3c == parameter_2_33 ? phv_data_60 : _GEN_2679; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2681 = 14'h3d == parameter_2_33 ? phv_data_61 : _GEN_2680; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2682 = 14'h3e == parameter_2_33 ? phv_data_62 : _GEN_2681; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2683 = 14'h3f == parameter_2_33 ? phv_data_63 : _GEN_2682; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_34 = vliw_34[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_34 = vliw_34[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_34 = parameter_2_34[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_34 = parameter_2_34[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_34 = {{1'd0}, args_offset_34}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_34 = _total_offset_T_34[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2687 = 3'h1 == total_offset_34 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2688 = 3'h2 == total_offset_34 ? args_2 : _GEN_2687; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2689 = 3'h3 == total_offset_34 ? args_3 : _GEN_2688; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2690 = 3'h4 == total_offset_34 ? args_4 : _GEN_2689; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2691 = 3'h5 == total_offset_34 ? args_5 : _GEN_2690; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2692 = 3'h6 == total_offset_34 ? args_6 : _GEN_2691; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2693 = total_offset_34 < 3'h7 ? _GEN_2692 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_34_0 = 3'h0 < args_length_34 ? _GEN_2693 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_2695 = opcode_34 == 4'ha ? field_bytes_34_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2696 = opcode_34 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2417 = opcode_34 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_69 = _T_2417 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_2697 = opcode_34 == 4'h8 | opcode_34 == 4'hb ? parameter_2_34[7:0] : _GEN_2695; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_2698 = opcode_34 == 4'h8 | opcode_34 == 4'hb ? _field_tag_T_69 : _GEN_2696; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_2699 = 14'h0 == parameter_2_34 ? phv_data_0 : _GEN_2697; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2700 = 14'h1 == parameter_2_34 ? phv_data_1 : _GEN_2699; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2701 = 14'h2 == parameter_2_34 ? phv_data_2 : _GEN_2700; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2702 = 14'h3 == parameter_2_34 ? phv_data_3 : _GEN_2701; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2703 = 14'h4 == parameter_2_34 ? phv_data_4 : _GEN_2702; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2704 = 14'h5 == parameter_2_34 ? phv_data_5 : _GEN_2703; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2705 = 14'h6 == parameter_2_34 ? phv_data_6 : _GEN_2704; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2706 = 14'h7 == parameter_2_34 ? phv_data_7 : _GEN_2705; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2707 = 14'h8 == parameter_2_34 ? phv_data_8 : _GEN_2706; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2708 = 14'h9 == parameter_2_34 ? phv_data_9 : _GEN_2707; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2709 = 14'ha == parameter_2_34 ? phv_data_10 : _GEN_2708; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2710 = 14'hb == parameter_2_34 ? phv_data_11 : _GEN_2709; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2711 = 14'hc == parameter_2_34 ? phv_data_12 : _GEN_2710; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2712 = 14'hd == parameter_2_34 ? phv_data_13 : _GEN_2711; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2713 = 14'he == parameter_2_34 ? phv_data_14 : _GEN_2712; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2714 = 14'hf == parameter_2_34 ? phv_data_15 : _GEN_2713; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2715 = 14'h10 == parameter_2_34 ? phv_data_16 : _GEN_2714; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2716 = 14'h11 == parameter_2_34 ? phv_data_17 : _GEN_2715; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2717 = 14'h12 == parameter_2_34 ? phv_data_18 : _GEN_2716; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2718 = 14'h13 == parameter_2_34 ? phv_data_19 : _GEN_2717; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2719 = 14'h14 == parameter_2_34 ? phv_data_20 : _GEN_2718; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2720 = 14'h15 == parameter_2_34 ? phv_data_21 : _GEN_2719; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2721 = 14'h16 == parameter_2_34 ? phv_data_22 : _GEN_2720; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2722 = 14'h17 == parameter_2_34 ? phv_data_23 : _GEN_2721; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2723 = 14'h18 == parameter_2_34 ? phv_data_24 : _GEN_2722; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2724 = 14'h19 == parameter_2_34 ? phv_data_25 : _GEN_2723; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2725 = 14'h1a == parameter_2_34 ? phv_data_26 : _GEN_2724; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2726 = 14'h1b == parameter_2_34 ? phv_data_27 : _GEN_2725; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2727 = 14'h1c == parameter_2_34 ? phv_data_28 : _GEN_2726; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2728 = 14'h1d == parameter_2_34 ? phv_data_29 : _GEN_2727; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2729 = 14'h1e == parameter_2_34 ? phv_data_30 : _GEN_2728; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2730 = 14'h1f == parameter_2_34 ? phv_data_31 : _GEN_2729; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2731 = 14'h20 == parameter_2_34 ? phv_data_32 : _GEN_2730; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2732 = 14'h21 == parameter_2_34 ? phv_data_33 : _GEN_2731; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2733 = 14'h22 == parameter_2_34 ? phv_data_34 : _GEN_2732; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2734 = 14'h23 == parameter_2_34 ? phv_data_35 : _GEN_2733; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2735 = 14'h24 == parameter_2_34 ? phv_data_36 : _GEN_2734; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2736 = 14'h25 == parameter_2_34 ? phv_data_37 : _GEN_2735; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2737 = 14'h26 == parameter_2_34 ? phv_data_38 : _GEN_2736; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2738 = 14'h27 == parameter_2_34 ? phv_data_39 : _GEN_2737; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2739 = 14'h28 == parameter_2_34 ? phv_data_40 : _GEN_2738; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2740 = 14'h29 == parameter_2_34 ? phv_data_41 : _GEN_2739; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2741 = 14'h2a == parameter_2_34 ? phv_data_42 : _GEN_2740; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2742 = 14'h2b == parameter_2_34 ? phv_data_43 : _GEN_2741; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2743 = 14'h2c == parameter_2_34 ? phv_data_44 : _GEN_2742; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2744 = 14'h2d == parameter_2_34 ? phv_data_45 : _GEN_2743; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2745 = 14'h2e == parameter_2_34 ? phv_data_46 : _GEN_2744; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2746 = 14'h2f == parameter_2_34 ? phv_data_47 : _GEN_2745; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2747 = 14'h30 == parameter_2_34 ? phv_data_48 : _GEN_2746; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2748 = 14'h31 == parameter_2_34 ? phv_data_49 : _GEN_2747; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2749 = 14'h32 == parameter_2_34 ? phv_data_50 : _GEN_2748; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2750 = 14'h33 == parameter_2_34 ? phv_data_51 : _GEN_2749; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2751 = 14'h34 == parameter_2_34 ? phv_data_52 : _GEN_2750; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2752 = 14'h35 == parameter_2_34 ? phv_data_53 : _GEN_2751; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2753 = 14'h36 == parameter_2_34 ? phv_data_54 : _GEN_2752; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2754 = 14'h37 == parameter_2_34 ? phv_data_55 : _GEN_2753; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2755 = 14'h38 == parameter_2_34 ? phv_data_56 : _GEN_2754; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2756 = 14'h39 == parameter_2_34 ? phv_data_57 : _GEN_2755; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2757 = 14'h3a == parameter_2_34 ? phv_data_58 : _GEN_2756; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2758 = 14'h3b == parameter_2_34 ? phv_data_59 : _GEN_2757; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2759 = 14'h3c == parameter_2_34 ? phv_data_60 : _GEN_2758; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2760 = 14'h3d == parameter_2_34 ? phv_data_61 : _GEN_2759; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2761 = 14'h3e == parameter_2_34 ? phv_data_62 : _GEN_2760; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2762 = 14'h3f == parameter_2_34 ? phv_data_63 : _GEN_2761; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_35 = vliw_35[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_35 = vliw_35[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_35 = parameter_2_35[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_35 = parameter_2_35[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_35 = {{1'd0}, args_offset_35}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_35 = _total_offset_T_35[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2766 = 3'h1 == total_offset_35 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2767 = 3'h2 == total_offset_35 ? args_2 : _GEN_2766; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2768 = 3'h3 == total_offset_35 ? args_3 : _GEN_2767; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2769 = 3'h4 == total_offset_35 ? args_4 : _GEN_2768; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2770 = 3'h5 == total_offset_35 ? args_5 : _GEN_2769; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2771 = 3'h6 == total_offset_35 ? args_6 : _GEN_2770; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2772 = total_offset_35 < 3'h7 ? _GEN_2771 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_35_0 = 3'h0 < args_length_35 ? _GEN_2772 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_2774 = opcode_35 == 4'ha ? field_bytes_35_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2775 = opcode_35 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2488 = opcode_35 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_71 = _T_2488 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_2776 = opcode_35 == 4'h8 | opcode_35 == 4'hb ? parameter_2_35[7:0] : _GEN_2774; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_2777 = opcode_35 == 4'h8 | opcode_35 == 4'hb ? _field_tag_T_71 : _GEN_2775; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_2778 = 14'h0 == parameter_2_35 ? phv_data_0 : _GEN_2776; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2779 = 14'h1 == parameter_2_35 ? phv_data_1 : _GEN_2778; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2780 = 14'h2 == parameter_2_35 ? phv_data_2 : _GEN_2779; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2781 = 14'h3 == parameter_2_35 ? phv_data_3 : _GEN_2780; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2782 = 14'h4 == parameter_2_35 ? phv_data_4 : _GEN_2781; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2783 = 14'h5 == parameter_2_35 ? phv_data_5 : _GEN_2782; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2784 = 14'h6 == parameter_2_35 ? phv_data_6 : _GEN_2783; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2785 = 14'h7 == parameter_2_35 ? phv_data_7 : _GEN_2784; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2786 = 14'h8 == parameter_2_35 ? phv_data_8 : _GEN_2785; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2787 = 14'h9 == parameter_2_35 ? phv_data_9 : _GEN_2786; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2788 = 14'ha == parameter_2_35 ? phv_data_10 : _GEN_2787; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2789 = 14'hb == parameter_2_35 ? phv_data_11 : _GEN_2788; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2790 = 14'hc == parameter_2_35 ? phv_data_12 : _GEN_2789; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2791 = 14'hd == parameter_2_35 ? phv_data_13 : _GEN_2790; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2792 = 14'he == parameter_2_35 ? phv_data_14 : _GEN_2791; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2793 = 14'hf == parameter_2_35 ? phv_data_15 : _GEN_2792; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2794 = 14'h10 == parameter_2_35 ? phv_data_16 : _GEN_2793; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2795 = 14'h11 == parameter_2_35 ? phv_data_17 : _GEN_2794; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2796 = 14'h12 == parameter_2_35 ? phv_data_18 : _GEN_2795; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2797 = 14'h13 == parameter_2_35 ? phv_data_19 : _GEN_2796; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2798 = 14'h14 == parameter_2_35 ? phv_data_20 : _GEN_2797; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2799 = 14'h15 == parameter_2_35 ? phv_data_21 : _GEN_2798; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2800 = 14'h16 == parameter_2_35 ? phv_data_22 : _GEN_2799; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2801 = 14'h17 == parameter_2_35 ? phv_data_23 : _GEN_2800; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2802 = 14'h18 == parameter_2_35 ? phv_data_24 : _GEN_2801; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2803 = 14'h19 == parameter_2_35 ? phv_data_25 : _GEN_2802; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2804 = 14'h1a == parameter_2_35 ? phv_data_26 : _GEN_2803; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2805 = 14'h1b == parameter_2_35 ? phv_data_27 : _GEN_2804; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2806 = 14'h1c == parameter_2_35 ? phv_data_28 : _GEN_2805; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2807 = 14'h1d == parameter_2_35 ? phv_data_29 : _GEN_2806; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2808 = 14'h1e == parameter_2_35 ? phv_data_30 : _GEN_2807; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2809 = 14'h1f == parameter_2_35 ? phv_data_31 : _GEN_2808; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2810 = 14'h20 == parameter_2_35 ? phv_data_32 : _GEN_2809; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2811 = 14'h21 == parameter_2_35 ? phv_data_33 : _GEN_2810; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2812 = 14'h22 == parameter_2_35 ? phv_data_34 : _GEN_2811; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2813 = 14'h23 == parameter_2_35 ? phv_data_35 : _GEN_2812; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2814 = 14'h24 == parameter_2_35 ? phv_data_36 : _GEN_2813; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2815 = 14'h25 == parameter_2_35 ? phv_data_37 : _GEN_2814; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2816 = 14'h26 == parameter_2_35 ? phv_data_38 : _GEN_2815; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2817 = 14'h27 == parameter_2_35 ? phv_data_39 : _GEN_2816; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2818 = 14'h28 == parameter_2_35 ? phv_data_40 : _GEN_2817; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2819 = 14'h29 == parameter_2_35 ? phv_data_41 : _GEN_2818; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2820 = 14'h2a == parameter_2_35 ? phv_data_42 : _GEN_2819; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2821 = 14'h2b == parameter_2_35 ? phv_data_43 : _GEN_2820; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2822 = 14'h2c == parameter_2_35 ? phv_data_44 : _GEN_2821; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2823 = 14'h2d == parameter_2_35 ? phv_data_45 : _GEN_2822; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2824 = 14'h2e == parameter_2_35 ? phv_data_46 : _GEN_2823; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2825 = 14'h2f == parameter_2_35 ? phv_data_47 : _GEN_2824; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2826 = 14'h30 == parameter_2_35 ? phv_data_48 : _GEN_2825; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2827 = 14'h31 == parameter_2_35 ? phv_data_49 : _GEN_2826; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2828 = 14'h32 == parameter_2_35 ? phv_data_50 : _GEN_2827; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2829 = 14'h33 == parameter_2_35 ? phv_data_51 : _GEN_2828; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2830 = 14'h34 == parameter_2_35 ? phv_data_52 : _GEN_2829; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2831 = 14'h35 == parameter_2_35 ? phv_data_53 : _GEN_2830; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2832 = 14'h36 == parameter_2_35 ? phv_data_54 : _GEN_2831; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2833 = 14'h37 == parameter_2_35 ? phv_data_55 : _GEN_2832; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2834 = 14'h38 == parameter_2_35 ? phv_data_56 : _GEN_2833; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2835 = 14'h39 == parameter_2_35 ? phv_data_57 : _GEN_2834; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2836 = 14'h3a == parameter_2_35 ? phv_data_58 : _GEN_2835; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2837 = 14'h3b == parameter_2_35 ? phv_data_59 : _GEN_2836; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2838 = 14'h3c == parameter_2_35 ? phv_data_60 : _GEN_2837; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2839 = 14'h3d == parameter_2_35 ? phv_data_61 : _GEN_2838; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2840 = 14'h3e == parameter_2_35 ? phv_data_62 : _GEN_2839; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2841 = 14'h3f == parameter_2_35 ? phv_data_63 : _GEN_2840; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_36 = vliw_36[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_36 = vliw_36[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_36 = parameter_2_36[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_36 = parameter_2_36[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_36 = {{1'd0}, args_offset_36}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_36 = _total_offset_T_36[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2845 = 3'h1 == total_offset_36 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2846 = 3'h2 == total_offset_36 ? args_2 : _GEN_2845; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2847 = 3'h3 == total_offset_36 ? args_3 : _GEN_2846; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2848 = 3'h4 == total_offset_36 ? args_4 : _GEN_2847; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2849 = 3'h5 == total_offset_36 ? args_5 : _GEN_2848; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2850 = 3'h6 == total_offset_36 ? args_6 : _GEN_2849; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2851 = total_offset_36 < 3'h7 ? _GEN_2850 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_36_0 = 3'h0 < args_length_36 ? _GEN_2851 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_2853 = opcode_36 == 4'ha ? field_bytes_36_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2854 = opcode_36 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2559 = opcode_36 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_73 = _T_2559 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_2855 = opcode_36 == 4'h8 | opcode_36 == 4'hb ? parameter_2_36[7:0] : _GEN_2853; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_2856 = opcode_36 == 4'h8 | opcode_36 == 4'hb ? _field_tag_T_73 : _GEN_2854; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_2857 = 14'h0 == parameter_2_36 ? phv_data_0 : _GEN_2855; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2858 = 14'h1 == parameter_2_36 ? phv_data_1 : _GEN_2857; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2859 = 14'h2 == parameter_2_36 ? phv_data_2 : _GEN_2858; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2860 = 14'h3 == parameter_2_36 ? phv_data_3 : _GEN_2859; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2861 = 14'h4 == parameter_2_36 ? phv_data_4 : _GEN_2860; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2862 = 14'h5 == parameter_2_36 ? phv_data_5 : _GEN_2861; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2863 = 14'h6 == parameter_2_36 ? phv_data_6 : _GEN_2862; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2864 = 14'h7 == parameter_2_36 ? phv_data_7 : _GEN_2863; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2865 = 14'h8 == parameter_2_36 ? phv_data_8 : _GEN_2864; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2866 = 14'h9 == parameter_2_36 ? phv_data_9 : _GEN_2865; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2867 = 14'ha == parameter_2_36 ? phv_data_10 : _GEN_2866; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2868 = 14'hb == parameter_2_36 ? phv_data_11 : _GEN_2867; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2869 = 14'hc == parameter_2_36 ? phv_data_12 : _GEN_2868; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2870 = 14'hd == parameter_2_36 ? phv_data_13 : _GEN_2869; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2871 = 14'he == parameter_2_36 ? phv_data_14 : _GEN_2870; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2872 = 14'hf == parameter_2_36 ? phv_data_15 : _GEN_2871; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2873 = 14'h10 == parameter_2_36 ? phv_data_16 : _GEN_2872; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2874 = 14'h11 == parameter_2_36 ? phv_data_17 : _GEN_2873; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2875 = 14'h12 == parameter_2_36 ? phv_data_18 : _GEN_2874; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2876 = 14'h13 == parameter_2_36 ? phv_data_19 : _GEN_2875; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2877 = 14'h14 == parameter_2_36 ? phv_data_20 : _GEN_2876; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2878 = 14'h15 == parameter_2_36 ? phv_data_21 : _GEN_2877; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2879 = 14'h16 == parameter_2_36 ? phv_data_22 : _GEN_2878; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2880 = 14'h17 == parameter_2_36 ? phv_data_23 : _GEN_2879; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2881 = 14'h18 == parameter_2_36 ? phv_data_24 : _GEN_2880; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2882 = 14'h19 == parameter_2_36 ? phv_data_25 : _GEN_2881; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2883 = 14'h1a == parameter_2_36 ? phv_data_26 : _GEN_2882; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2884 = 14'h1b == parameter_2_36 ? phv_data_27 : _GEN_2883; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2885 = 14'h1c == parameter_2_36 ? phv_data_28 : _GEN_2884; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2886 = 14'h1d == parameter_2_36 ? phv_data_29 : _GEN_2885; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2887 = 14'h1e == parameter_2_36 ? phv_data_30 : _GEN_2886; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2888 = 14'h1f == parameter_2_36 ? phv_data_31 : _GEN_2887; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2889 = 14'h20 == parameter_2_36 ? phv_data_32 : _GEN_2888; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2890 = 14'h21 == parameter_2_36 ? phv_data_33 : _GEN_2889; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2891 = 14'h22 == parameter_2_36 ? phv_data_34 : _GEN_2890; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2892 = 14'h23 == parameter_2_36 ? phv_data_35 : _GEN_2891; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2893 = 14'h24 == parameter_2_36 ? phv_data_36 : _GEN_2892; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2894 = 14'h25 == parameter_2_36 ? phv_data_37 : _GEN_2893; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2895 = 14'h26 == parameter_2_36 ? phv_data_38 : _GEN_2894; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2896 = 14'h27 == parameter_2_36 ? phv_data_39 : _GEN_2895; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2897 = 14'h28 == parameter_2_36 ? phv_data_40 : _GEN_2896; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2898 = 14'h29 == parameter_2_36 ? phv_data_41 : _GEN_2897; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2899 = 14'h2a == parameter_2_36 ? phv_data_42 : _GEN_2898; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2900 = 14'h2b == parameter_2_36 ? phv_data_43 : _GEN_2899; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2901 = 14'h2c == parameter_2_36 ? phv_data_44 : _GEN_2900; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2902 = 14'h2d == parameter_2_36 ? phv_data_45 : _GEN_2901; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2903 = 14'h2e == parameter_2_36 ? phv_data_46 : _GEN_2902; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2904 = 14'h2f == parameter_2_36 ? phv_data_47 : _GEN_2903; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2905 = 14'h30 == parameter_2_36 ? phv_data_48 : _GEN_2904; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2906 = 14'h31 == parameter_2_36 ? phv_data_49 : _GEN_2905; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2907 = 14'h32 == parameter_2_36 ? phv_data_50 : _GEN_2906; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2908 = 14'h33 == parameter_2_36 ? phv_data_51 : _GEN_2907; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2909 = 14'h34 == parameter_2_36 ? phv_data_52 : _GEN_2908; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2910 = 14'h35 == parameter_2_36 ? phv_data_53 : _GEN_2909; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2911 = 14'h36 == parameter_2_36 ? phv_data_54 : _GEN_2910; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2912 = 14'h37 == parameter_2_36 ? phv_data_55 : _GEN_2911; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2913 = 14'h38 == parameter_2_36 ? phv_data_56 : _GEN_2912; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2914 = 14'h39 == parameter_2_36 ? phv_data_57 : _GEN_2913; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2915 = 14'h3a == parameter_2_36 ? phv_data_58 : _GEN_2914; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2916 = 14'h3b == parameter_2_36 ? phv_data_59 : _GEN_2915; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2917 = 14'h3c == parameter_2_36 ? phv_data_60 : _GEN_2916; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2918 = 14'h3d == parameter_2_36 ? phv_data_61 : _GEN_2917; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2919 = 14'h3e == parameter_2_36 ? phv_data_62 : _GEN_2918; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2920 = 14'h3f == parameter_2_36 ? phv_data_63 : _GEN_2919; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_37 = vliw_37[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_37 = vliw_37[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_37 = parameter_2_37[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_37 = parameter_2_37[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_37 = {{1'd0}, args_offset_37}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_37 = _total_offset_T_37[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2924 = 3'h1 == total_offset_37 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2925 = 3'h2 == total_offset_37 ? args_2 : _GEN_2924; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2926 = 3'h3 == total_offset_37 ? args_3 : _GEN_2925; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2927 = 3'h4 == total_offset_37 ? args_4 : _GEN_2926; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2928 = 3'h5 == total_offset_37 ? args_5 : _GEN_2927; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2929 = 3'h6 == total_offset_37 ? args_6 : _GEN_2928; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2930 = total_offset_37 < 3'h7 ? _GEN_2929 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_37_0 = 3'h0 < args_length_37 ? _GEN_2930 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_2932 = opcode_37 == 4'ha ? field_bytes_37_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2933 = opcode_37 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2630 = opcode_37 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_75 = _T_2630 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_2934 = opcode_37 == 4'h8 | opcode_37 == 4'hb ? parameter_2_37[7:0] : _GEN_2932; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_2935 = opcode_37 == 4'h8 | opcode_37 == 4'hb ? _field_tag_T_75 : _GEN_2933; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_2936 = 14'h0 == parameter_2_37 ? phv_data_0 : _GEN_2934; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2937 = 14'h1 == parameter_2_37 ? phv_data_1 : _GEN_2936; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2938 = 14'h2 == parameter_2_37 ? phv_data_2 : _GEN_2937; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2939 = 14'h3 == parameter_2_37 ? phv_data_3 : _GEN_2938; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2940 = 14'h4 == parameter_2_37 ? phv_data_4 : _GEN_2939; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2941 = 14'h5 == parameter_2_37 ? phv_data_5 : _GEN_2940; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2942 = 14'h6 == parameter_2_37 ? phv_data_6 : _GEN_2941; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2943 = 14'h7 == parameter_2_37 ? phv_data_7 : _GEN_2942; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2944 = 14'h8 == parameter_2_37 ? phv_data_8 : _GEN_2943; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2945 = 14'h9 == parameter_2_37 ? phv_data_9 : _GEN_2944; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2946 = 14'ha == parameter_2_37 ? phv_data_10 : _GEN_2945; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2947 = 14'hb == parameter_2_37 ? phv_data_11 : _GEN_2946; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2948 = 14'hc == parameter_2_37 ? phv_data_12 : _GEN_2947; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2949 = 14'hd == parameter_2_37 ? phv_data_13 : _GEN_2948; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2950 = 14'he == parameter_2_37 ? phv_data_14 : _GEN_2949; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2951 = 14'hf == parameter_2_37 ? phv_data_15 : _GEN_2950; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2952 = 14'h10 == parameter_2_37 ? phv_data_16 : _GEN_2951; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2953 = 14'h11 == parameter_2_37 ? phv_data_17 : _GEN_2952; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2954 = 14'h12 == parameter_2_37 ? phv_data_18 : _GEN_2953; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2955 = 14'h13 == parameter_2_37 ? phv_data_19 : _GEN_2954; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2956 = 14'h14 == parameter_2_37 ? phv_data_20 : _GEN_2955; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2957 = 14'h15 == parameter_2_37 ? phv_data_21 : _GEN_2956; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2958 = 14'h16 == parameter_2_37 ? phv_data_22 : _GEN_2957; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2959 = 14'h17 == parameter_2_37 ? phv_data_23 : _GEN_2958; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2960 = 14'h18 == parameter_2_37 ? phv_data_24 : _GEN_2959; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2961 = 14'h19 == parameter_2_37 ? phv_data_25 : _GEN_2960; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2962 = 14'h1a == parameter_2_37 ? phv_data_26 : _GEN_2961; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2963 = 14'h1b == parameter_2_37 ? phv_data_27 : _GEN_2962; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2964 = 14'h1c == parameter_2_37 ? phv_data_28 : _GEN_2963; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2965 = 14'h1d == parameter_2_37 ? phv_data_29 : _GEN_2964; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2966 = 14'h1e == parameter_2_37 ? phv_data_30 : _GEN_2965; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2967 = 14'h1f == parameter_2_37 ? phv_data_31 : _GEN_2966; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2968 = 14'h20 == parameter_2_37 ? phv_data_32 : _GEN_2967; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2969 = 14'h21 == parameter_2_37 ? phv_data_33 : _GEN_2968; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2970 = 14'h22 == parameter_2_37 ? phv_data_34 : _GEN_2969; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2971 = 14'h23 == parameter_2_37 ? phv_data_35 : _GEN_2970; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2972 = 14'h24 == parameter_2_37 ? phv_data_36 : _GEN_2971; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2973 = 14'h25 == parameter_2_37 ? phv_data_37 : _GEN_2972; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2974 = 14'h26 == parameter_2_37 ? phv_data_38 : _GEN_2973; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2975 = 14'h27 == parameter_2_37 ? phv_data_39 : _GEN_2974; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2976 = 14'h28 == parameter_2_37 ? phv_data_40 : _GEN_2975; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2977 = 14'h29 == parameter_2_37 ? phv_data_41 : _GEN_2976; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2978 = 14'h2a == parameter_2_37 ? phv_data_42 : _GEN_2977; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2979 = 14'h2b == parameter_2_37 ? phv_data_43 : _GEN_2978; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2980 = 14'h2c == parameter_2_37 ? phv_data_44 : _GEN_2979; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2981 = 14'h2d == parameter_2_37 ? phv_data_45 : _GEN_2980; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2982 = 14'h2e == parameter_2_37 ? phv_data_46 : _GEN_2981; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2983 = 14'h2f == parameter_2_37 ? phv_data_47 : _GEN_2982; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2984 = 14'h30 == parameter_2_37 ? phv_data_48 : _GEN_2983; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2985 = 14'h31 == parameter_2_37 ? phv_data_49 : _GEN_2984; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2986 = 14'h32 == parameter_2_37 ? phv_data_50 : _GEN_2985; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2987 = 14'h33 == parameter_2_37 ? phv_data_51 : _GEN_2986; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2988 = 14'h34 == parameter_2_37 ? phv_data_52 : _GEN_2987; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2989 = 14'h35 == parameter_2_37 ? phv_data_53 : _GEN_2988; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2990 = 14'h36 == parameter_2_37 ? phv_data_54 : _GEN_2989; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2991 = 14'h37 == parameter_2_37 ? phv_data_55 : _GEN_2990; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2992 = 14'h38 == parameter_2_37 ? phv_data_56 : _GEN_2991; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2993 = 14'h39 == parameter_2_37 ? phv_data_57 : _GEN_2992; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2994 = 14'h3a == parameter_2_37 ? phv_data_58 : _GEN_2993; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2995 = 14'h3b == parameter_2_37 ? phv_data_59 : _GEN_2994; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2996 = 14'h3c == parameter_2_37 ? phv_data_60 : _GEN_2995; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2997 = 14'h3d == parameter_2_37 ? phv_data_61 : _GEN_2996; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2998 = 14'h3e == parameter_2_37 ? phv_data_62 : _GEN_2997; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_2999 = 14'h3f == parameter_2_37 ? phv_data_63 : _GEN_2998; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_38 = vliw_38[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_38 = vliw_38[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_38 = parameter_2_38[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_38 = parameter_2_38[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_38 = {{1'd0}, args_offset_38}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_38 = _total_offset_T_38[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3003 = 3'h1 == total_offset_38 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3004 = 3'h2 == total_offset_38 ? args_2 : _GEN_3003; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3005 = 3'h3 == total_offset_38 ? args_3 : _GEN_3004; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3006 = 3'h4 == total_offset_38 ? args_4 : _GEN_3005; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3007 = 3'h5 == total_offset_38 ? args_5 : _GEN_3006; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3008 = 3'h6 == total_offset_38 ? args_6 : _GEN_3007; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3009 = total_offset_38 < 3'h7 ? _GEN_3008 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_38_0 = 3'h0 < args_length_38 ? _GEN_3009 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_3011 = opcode_38 == 4'ha ? field_bytes_38_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3012 = opcode_38 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2701 = opcode_38 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_77 = _T_2701 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_3013 = opcode_38 == 4'h8 | opcode_38 == 4'hb ? parameter_2_38[7:0] : _GEN_3011; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_3014 = opcode_38 == 4'h8 | opcode_38 == 4'hb ? _field_tag_T_77 : _GEN_3012; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_3015 = 14'h0 == parameter_2_38 ? phv_data_0 : _GEN_3013; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3016 = 14'h1 == parameter_2_38 ? phv_data_1 : _GEN_3015; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3017 = 14'h2 == parameter_2_38 ? phv_data_2 : _GEN_3016; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3018 = 14'h3 == parameter_2_38 ? phv_data_3 : _GEN_3017; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3019 = 14'h4 == parameter_2_38 ? phv_data_4 : _GEN_3018; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3020 = 14'h5 == parameter_2_38 ? phv_data_5 : _GEN_3019; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3021 = 14'h6 == parameter_2_38 ? phv_data_6 : _GEN_3020; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3022 = 14'h7 == parameter_2_38 ? phv_data_7 : _GEN_3021; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3023 = 14'h8 == parameter_2_38 ? phv_data_8 : _GEN_3022; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3024 = 14'h9 == parameter_2_38 ? phv_data_9 : _GEN_3023; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3025 = 14'ha == parameter_2_38 ? phv_data_10 : _GEN_3024; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3026 = 14'hb == parameter_2_38 ? phv_data_11 : _GEN_3025; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3027 = 14'hc == parameter_2_38 ? phv_data_12 : _GEN_3026; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3028 = 14'hd == parameter_2_38 ? phv_data_13 : _GEN_3027; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3029 = 14'he == parameter_2_38 ? phv_data_14 : _GEN_3028; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3030 = 14'hf == parameter_2_38 ? phv_data_15 : _GEN_3029; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3031 = 14'h10 == parameter_2_38 ? phv_data_16 : _GEN_3030; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3032 = 14'h11 == parameter_2_38 ? phv_data_17 : _GEN_3031; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3033 = 14'h12 == parameter_2_38 ? phv_data_18 : _GEN_3032; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3034 = 14'h13 == parameter_2_38 ? phv_data_19 : _GEN_3033; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3035 = 14'h14 == parameter_2_38 ? phv_data_20 : _GEN_3034; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3036 = 14'h15 == parameter_2_38 ? phv_data_21 : _GEN_3035; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3037 = 14'h16 == parameter_2_38 ? phv_data_22 : _GEN_3036; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3038 = 14'h17 == parameter_2_38 ? phv_data_23 : _GEN_3037; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3039 = 14'h18 == parameter_2_38 ? phv_data_24 : _GEN_3038; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3040 = 14'h19 == parameter_2_38 ? phv_data_25 : _GEN_3039; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3041 = 14'h1a == parameter_2_38 ? phv_data_26 : _GEN_3040; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3042 = 14'h1b == parameter_2_38 ? phv_data_27 : _GEN_3041; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3043 = 14'h1c == parameter_2_38 ? phv_data_28 : _GEN_3042; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3044 = 14'h1d == parameter_2_38 ? phv_data_29 : _GEN_3043; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3045 = 14'h1e == parameter_2_38 ? phv_data_30 : _GEN_3044; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3046 = 14'h1f == parameter_2_38 ? phv_data_31 : _GEN_3045; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3047 = 14'h20 == parameter_2_38 ? phv_data_32 : _GEN_3046; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3048 = 14'h21 == parameter_2_38 ? phv_data_33 : _GEN_3047; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3049 = 14'h22 == parameter_2_38 ? phv_data_34 : _GEN_3048; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3050 = 14'h23 == parameter_2_38 ? phv_data_35 : _GEN_3049; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3051 = 14'h24 == parameter_2_38 ? phv_data_36 : _GEN_3050; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3052 = 14'h25 == parameter_2_38 ? phv_data_37 : _GEN_3051; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3053 = 14'h26 == parameter_2_38 ? phv_data_38 : _GEN_3052; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3054 = 14'h27 == parameter_2_38 ? phv_data_39 : _GEN_3053; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3055 = 14'h28 == parameter_2_38 ? phv_data_40 : _GEN_3054; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3056 = 14'h29 == parameter_2_38 ? phv_data_41 : _GEN_3055; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3057 = 14'h2a == parameter_2_38 ? phv_data_42 : _GEN_3056; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3058 = 14'h2b == parameter_2_38 ? phv_data_43 : _GEN_3057; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3059 = 14'h2c == parameter_2_38 ? phv_data_44 : _GEN_3058; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3060 = 14'h2d == parameter_2_38 ? phv_data_45 : _GEN_3059; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3061 = 14'h2e == parameter_2_38 ? phv_data_46 : _GEN_3060; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3062 = 14'h2f == parameter_2_38 ? phv_data_47 : _GEN_3061; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3063 = 14'h30 == parameter_2_38 ? phv_data_48 : _GEN_3062; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3064 = 14'h31 == parameter_2_38 ? phv_data_49 : _GEN_3063; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3065 = 14'h32 == parameter_2_38 ? phv_data_50 : _GEN_3064; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3066 = 14'h33 == parameter_2_38 ? phv_data_51 : _GEN_3065; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3067 = 14'h34 == parameter_2_38 ? phv_data_52 : _GEN_3066; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3068 = 14'h35 == parameter_2_38 ? phv_data_53 : _GEN_3067; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3069 = 14'h36 == parameter_2_38 ? phv_data_54 : _GEN_3068; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3070 = 14'h37 == parameter_2_38 ? phv_data_55 : _GEN_3069; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3071 = 14'h38 == parameter_2_38 ? phv_data_56 : _GEN_3070; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3072 = 14'h39 == parameter_2_38 ? phv_data_57 : _GEN_3071; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3073 = 14'h3a == parameter_2_38 ? phv_data_58 : _GEN_3072; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3074 = 14'h3b == parameter_2_38 ? phv_data_59 : _GEN_3073; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3075 = 14'h3c == parameter_2_38 ? phv_data_60 : _GEN_3074; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3076 = 14'h3d == parameter_2_38 ? phv_data_61 : _GEN_3075; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3077 = 14'h3e == parameter_2_38 ? phv_data_62 : _GEN_3076; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3078 = 14'h3f == parameter_2_38 ? phv_data_63 : _GEN_3077; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_39 = vliw_39[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_39 = vliw_39[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_39 = parameter_2_39[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_39 = parameter_2_39[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_39 = {{1'd0}, args_offset_39}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_39 = _total_offset_T_39[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3082 = 3'h1 == total_offset_39 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3083 = 3'h2 == total_offset_39 ? args_2 : _GEN_3082; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3084 = 3'h3 == total_offset_39 ? args_3 : _GEN_3083; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3085 = 3'h4 == total_offset_39 ? args_4 : _GEN_3084; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3086 = 3'h5 == total_offset_39 ? args_5 : _GEN_3085; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3087 = 3'h6 == total_offset_39 ? args_6 : _GEN_3086; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3088 = total_offset_39 < 3'h7 ? _GEN_3087 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_39_0 = 3'h0 < args_length_39 ? _GEN_3088 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_3090 = opcode_39 == 4'ha ? field_bytes_39_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3091 = opcode_39 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2772 = opcode_39 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_79 = _T_2772 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_3092 = opcode_39 == 4'h8 | opcode_39 == 4'hb ? parameter_2_39[7:0] : _GEN_3090; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_3093 = opcode_39 == 4'h8 | opcode_39 == 4'hb ? _field_tag_T_79 : _GEN_3091; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_3094 = 14'h0 == parameter_2_39 ? phv_data_0 : _GEN_3092; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3095 = 14'h1 == parameter_2_39 ? phv_data_1 : _GEN_3094; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3096 = 14'h2 == parameter_2_39 ? phv_data_2 : _GEN_3095; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3097 = 14'h3 == parameter_2_39 ? phv_data_3 : _GEN_3096; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3098 = 14'h4 == parameter_2_39 ? phv_data_4 : _GEN_3097; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3099 = 14'h5 == parameter_2_39 ? phv_data_5 : _GEN_3098; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3100 = 14'h6 == parameter_2_39 ? phv_data_6 : _GEN_3099; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3101 = 14'h7 == parameter_2_39 ? phv_data_7 : _GEN_3100; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3102 = 14'h8 == parameter_2_39 ? phv_data_8 : _GEN_3101; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3103 = 14'h9 == parameter_2_39 ? phv_data_9 : _GEN_3102; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3104 = 14'ha == parameter_2_39 ? phv_data_10 : _GEN_3103; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3105 = 14'hb == parameter_2_39 ? phv_data_11 : _GEN_3104; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3106 = 14'hc == parameter_2_39 ? phv_data_12 : _GEN_3105; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3107 = 14'hd == parameter_2_39 ? phv_data_13 : _GEN_3106; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3108 = 14'he == parameter_2_39 ? phv_data_14 : _GEN_3107; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3109 = 14'hf == parameter_2_39 ? phv_data_15 : _GEN_3108; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3110 = 14'h10 == parameter_2_39 ? phv_data_16 : _GEN_3109; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3111 = 14'h11 == parameter_2_39 ? phv_data_17 : _GEN_3110; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3112 = 14'h12 == parameter_2_39 ? phv_data_18 : _GEN_3111; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3113 = 14'h13 == parameter_2_39 ? phv_data_19 : _GEN_3112; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3114 = 14'h14 == parameter_2_39 ? phv_data_20 : _GEN_3113; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3115 = 14'h15 == parameter_2_39 ? phv_data_21 : _GEN_3114; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3116 = 14'h16 == parameter_2_39 ? phv_data_22 : _GEN_3115; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3117 = 14'h17 == parameter_2_39 ? phv_data_23 : _GEN_3116; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3118 = 14'h18 == parameter_2_39 ? phv_data_24 : _GEN_3117; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3119 = 14'h19 == parameter_2_39 ? phv_data_25 : _GEN_3118; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3120 = 14'h1a == parameter_2_39 ? phv_data_26 : _GEN_3119; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3121 = 14'h1b == parameter_2_39 ? phv_data_27 : _GEN_3120; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3122 = 14'h1c == parameter_2_39 ? phv_data_28 : _GEN_3121; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3123 = 14'h1d == parameter_2_39 ? phv_data_29 : _GEN_3122; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3124 = 14'h1e == parameter_2_39 ? phv_data_30 : _GEN_3123; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3125 = 14'h1f == parameter_2_39 ? phv_data_31 : _GEN_3124; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3126 = 14'h20 == parameter_2_39 ? phv_data_32 : _GEN_3125; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3127 = 14'h21 == parameter_2_39 ? phv_data_33 : _GEN_3126; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3128 = 14'h22 == parameter_2_39 ? phv_data_34 : _GEN_3127; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3129 = 14'h23 == parameter_2_39 ? phv_data_35 : _GEN_3128; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3130 = 14'h24 == parameter_2_39 ? phv_data_36 : _GEN_3129; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3131 = 14'h25 == parameter_2_39 ? phv_data_37 : _GEN_3130; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3132 = 14'h26 == parameter_2_39 ? phv_data_38 : _GEN_3131; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3133 = 14'h27 == parameter_2_39 ? phv_data_39 : _GEN_3132; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3134 = 14'h28 == parameter_2_39 ? phv_data_40 : _GEN_3133; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3135 = 14'h29 == parameter_2_39 ? phv_data_41 : _GEN_3134; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3136 = 14'h2a == parameter_2_39 ? phv_data_42 : _GEN_3135; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3137 = 14'h2b == parameter_2_39 ? phv_data_43 : _GEN_3136; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3138 = 14'h2c == parameter_2_39 ? phv_data_44 : _GEN_3137; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3139 = 14'h2d == parameter_2_39 ? phv_data_45 : _GEN_3138; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3140 = 14'h2e == parameter_2_39 ? phv_data_46 : _GEN_3139; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3141 = 14'h2f == parameter_2_39 ? phv_data_47 : _GEN_3140; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3142 = 14'h30 == parameter_2_39 ? phv_data_48 : _GEN_3141; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3143 = 14'h31 == parameter_2_39 ? phv_data_49 : _GEN_3142; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3144 = 14'h32 == parameter_2_39 ? phv_data_50 : _GEN_3143; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3145 = 14'h33 == parameter_2_39 ? phv_data_51 : _GEN_3144; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3146 = 14'h34 == parameter_2_39 ? phv_data_52 : _GEN_3145; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3147 = 14'h35 == parameter_2_39 ? phv_data_53 : _GEN_3146; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3148 = 14'h36 == parameter_2_39 ? phv_data_54 : _GEN_3147; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3149 = 14'h37 == parameter_2_39 ? phv_data_55 : _GEN_3148; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3150 = 14'h38 == parameter_2_39 ? phv_data_56 : _GEN_3149; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3151 = 14'h39 == parameter_2_39 ? phv_data_57 : _GEN_3150; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3152 = 14'h3a == parameter_2_39 ? phv_data_58 : _GEN_3151; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3153 = 14'h3b == parameter_2_39 ? phv_data_59 : _GEN_3152; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3154 = 14'h3c == parameter_2_39 ? phv_data_60 : _GEN_3153; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3155 = 14'h3d == parameter_2_39 ? phv_data_61 : _GEN_3154; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3156 = 14'h3e == parameter_2_39 ? phv_data_62 : _GEN_3155; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3157 = 14'h3f == parameter_2_39 ? phv_data_63 : _GEN_3156; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_40 = vliw_40[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_40 = vliw_40[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_40 = parameter_2_40[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_40 = parameter_2_40[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_40 = {{1'd0}, args_offset_40}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_40 = _total_offset_T_40[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3161 = 3'h1 == total_offset_40 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3162 = 3'h2 == total_offset_40 ? args_2 : _GEN_3161; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3163 = 3'h3 == total_offset_40 ? args_3 : _GEN_3162; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3164 = 3'h4 == total_offset_40 ? args_4 : _GEN_3163; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3165 = 3'h5 == total_offset_40 ? args_5 : _GEN_3164; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3166 = 3'h6 == total_offset_40 ? args_6 : _GEN_3165; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3167 = total_offset_40 < 3'h7 ? _GEN_3166 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_40_0 = 3'h0 < args_length_40 ? _GEN_3167 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_3169 = opcode_40 == 4'ha ? field_bytes_40_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3170 = opcode_40 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2843 = opcode_40 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_81 = _T_2843 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_3171 = opcode_40 == 4'h8 | opcode_40 == 4'hb ? parameter_2_40[7:0] : _GEN_3169; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_3172 = opcode_40 == 4'h8 | opcode_40 == 4'hb ? _field_tag_T_81 : _GEN_3170; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_3173 = 14'h0 == parameter_2_40 ? phv_data_0 : _GEN_3171; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3174 = 14'h1 == parameter_2_40 ? phv_data_1 : _GEN_3173; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3175 = 14'h2 == parameter_2_40 ? phv_data_2 : _GEN_3174; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3176 = 14'h3 == parameter_2_40 ? phv_data_3 : _GEN_3175; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3177 = 14'h4 == parameter_2_40 ? phv_data_4 : _GEN_3176; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3178 = 14'h5 == parameter_2_40 ? phv_data_5 : _GEN_3177; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3179 = 14'h6 == parameter_2_40 ? phv_data_6 : _GEN_3178; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3180 = 14'h7 == parameter_2_40 ? phv_data_7 : _GEN_3179; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3181 = 14'h8 == parameter_2_40 ? phv_data_8 : _GEN_3180; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3182 = 14'h9 == parameter_2_40 ? phv_data_9 : _GEN_3181; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3183 = 14'ha == parameter_2_40 ? phv_data_10 : _GEN_3182; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3184 = 14'hb == parameter_2_40 ? phv_data_11 : _GEN_3183; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3185 = 14'hc == parameter_2_40 ? phv_data_12 : _GEN_3184; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3186 = 14'hd == parameter_2_40 ? phv_data_13 : _GEN_3185; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3187 = 14'he == parameter_2_40 ? phv_data_14 : _GEN_3186; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3188 = 14'hf == parameter_2_40 ? phv_data_15 : _GEN_3187; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3189 = 14'h10 == parameter_2_40 ? phv_data_16 : _GEN_3188; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3190 = 14'h11 == parameter_2_40 ? phv_data_17 : _GEN_3189; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3191 = 14'h12 == parameter_2_40 ? phv_data_18 : _GEN_3190; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3192 = 14'h13 == parameter_2_40 ? phv_data_19 : _GEN_3191; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3193 = 14'h14 == parameter_2_40 ? phv_data_20 : _GEN_3192; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3194 = 14'h15 == parameter_2_40 ? phv_data_21 : _GEN_3193; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3195 = 14'h16 == parameter_2_40 ? phv_data_22 : _GEN_3194; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3196 = 14'h17 == parameter_2_40 ? phv_data_23 : _GEN_3195; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3197 = 14'h18 == parameter_2_40 ? phv_data_24 : _GEN_3196; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3198 = 14'h19 == parameter_2_40 ? phv_data_25 : _GEN_3197; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3199 = 14'h1a == parameter_2_40 ? phv_data_26 : _GEN_3198; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3200 = 14'h1b == parameter_2_40 ? phv_data_27 : _GEN_3199; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3201 = 14'h1c == parameter_2_40 ? phv_data_28 : _GEN_3200; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3202 = 14'h1d == parameter_2_40 ? phv_data_29 : _GEN_3201; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3203 = 14'h1e == parameter_2_40 ? phv_data_30 : _GEN_3202; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3204 = 14'h1f == parameter_2_40 ? phv_data_31 : _GEN_3203; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3205 = 14'h20 == parameter_2_40 ? phv_data_32 : _GEN_3204; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3206 = 14'h21 == parameter_2_40 ? phv_data_33 : _GEN_3205; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3207 = 14'h22 == parameter_2_40 ? phv_data_34 : _GEN_3206; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3208 = 14'h23 == parameter_2_40 ? phv_data_35 : _GEN_3207; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3209 = 14'h24 == parameter_2_40 ? phv_data_36 : _GEN_3208; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3210 = 14'h25 == parameter_2_40 ? phv_data_37 : _GEN_3209; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3211 = 14'h26 == parameter_2_40 ? phv_data_38 : _GEN_3210; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3212 = 14'h27 == parameter_2_40 ? phv_data_39 : _GEN_3211; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3213 = 14'h28 == parameter_2_40 ? phv_data_40 : _GEN_3212; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3214 = 14'h29 == parameter_2_40 ? phv_data_41 : _GEN_3213; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3215 = 14'h2a == parameter_2_40 ? phv_data_42 : _GEN_3214; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3216 = 14'h2b == parameter_2_40 ? phv_data_43 : _GEN_3215; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3217 = 14'h2c == parameter_2_40 ? phv_data_44 : _GEN_3216; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3218 = 14'h2d == parameter_2_40 ? phv_data_45 : _GEN_3217; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3219 = 14'h2e == parameter_2_40 ? phv_data_46 : _GEN_3218; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3220 = 14'h2f == parameter_2_40 ? phv_data_47 : _GEN_3219; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3221 = 14'h30 == parameter_2_40 ? phv_data_48 : _GEN_3220; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3222 = 14'h31 == parameter_2_40 ? phv_data_49 : _GEN_3221; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3223 = 14'h32 == parameter_2_40 ? phv_data_50 : _GEN_3222; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3224 = 14'h33 == parameter_2_40 ? phv_data_51 : _GEN_3223; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3225 = 14'h34 == parameter_2_40 ? phv_data_52 : _GEN_3224; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3226 = 14'h35 == parameter_2_40 ? phv_data_53 : _GEN_3225; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3227 = 14'h36 == parameter_2_40 ? phv_data_54 : _GEN_3226; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3228 = 14'h37 == parameter_2_40 ? phv_data_55 : _GEN_3227; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3229 = 14'h38 == parameter_2_40 ? phv_data_56 : _GEN_3228; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3230 = 14'h39 == parameter_2_40 ? phv_data_57 : _GEN_3229; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3231 = 14'h3a == parameter_2_40 ? phv_data_58 : _GEN_3230; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3232 = 14'h3b == parameter_2_40 ? phv_data_59 : _GEN_3231; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3233 = 14'h3c == parameter_2_40 ? phv_data_60 : _GEN_3232; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3234 = 14'h3d == parameter_2_40 ? phv_data_61 : _GEN_3233; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3235 = 14'h3e == parameter_2_40 ? phv_data_62 : _GEN_3234; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3236 = 14'h3f == parameter_2_40 ? phv_data_63 : _GEN_3235; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_41 = vliw_41[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_41 = vliw_41[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_41 = parameter_2_41[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_41 = parameter_2_41[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_41 = {{1'd0}, args_offset_41}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_41 = _total_offset_T_41[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3240 = 3'h1 == total_offset_41 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3241 = 3'h2 == total_offset_41 ? args_2 : _GEN_3240; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3242 = 3'h3 == total_offset_41 ? args_3 : _GEN_3241; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3243 = 3'h4 == total_offset_41 ? args_4 : _GEN_3242; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3244 = 3'h5 == total_offset_41 ? args_5 : _GEN_3243; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3245 = 3'h6 == total_offset_41 ? args_6 : _GEN_3244; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3246 = total_offset_41 < 3'h7 ? _GEN_3245 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_41_0 = 3'h0 < args_length_41 ? _GEN_3246 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_3248 = opcode_41 == 4'ha ? field_bytes_41_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3249 = opcode_41 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2914 = opcode_41 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_83 = _T_2914 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_3250 = opcode_41 == 4'h8 | opcode_41 == 4'hb ? parameter_2_41[7:0] : _GEN_3248; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_3251 = opcode_41 == 4'h8 | opcode_41 == 4'hb ? _field_tag_T_83 : _GEN_3249; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_3252 = 14'h0 == parameter_2_41 ? phv_data_0 : _GEN_3250; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3253 = 14'h1 == parameter_2_41 ? phv_data_1 : _GEN_3252; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3254 = 14'h2 == parameter_2_41 ? phv_data_2 : _GEN_3253; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3255 = 14'h3 == parameter_2_41 ? phv_data_3 : _GEN_3254; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3256 = 14'h4 == parameter_2_41 ? phv_data_4 : _GEN_3255; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3257 = 14'h5 == parameter_2_41 ? phv_data_5 : _GEN_3256; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3258 = 14'h6 == parameter_2_41 ? phv_data_6 : _GEN_3257; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3259 = 14'h7 == parameter_2_41 ? phv_data_7 : _GEN_3258; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3260 = 14'h8 == parameter_2_41 ? phv_data_8 : _GEN_3259; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3261 = 14'h9 == parameter_2_41 ? phv_data_9 : _GEN_3260; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3262 = 14'ha == parameter_2_41 ? phv_data_10 : _GEN_3261; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3263 = 14'hb == parameter_2_41 ? phv_data_11 : _GEN_3262; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3264 = 14'hc == parameter_2_41 ? phv_data_12 : _GEN_3263; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3265 = 14'hd == parameter_2_41 ? phv_data_13 : _GEN_3264; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3266 = 14'he == parameter_2_41 ? phv_data_14 : _GEN_3265; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3267 = 14'hf == parameter_2_41 ? phv_data_15 : _GEN_3266; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3268 = 14'h10 == parameter_2_41 ? phv_data_16 : _GEN_3267; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3269 = 14'h11 == parameter_2_41 ? phv_data_17 : _GEN_3268; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3270 = 14'h12 == parameter_2_41 ? phv_data_18 : _GEN_3269; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3271 = 14'h13 == parameter_2_41 ? phv_data_19 : _GEN_3270; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3272 = 14'h14 == parameter_2_41 ? phv_data_20 : _GEN_3271; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3273 = 14'h15 == parameter_2_41 ? phv_data_21 : _GEN_3272; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3274 = 14'h16 == parameter_2_41 ? phv_data_22 : _GEN_3273; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3275 = 14'h17 == parameter_2_41 ? phv_data_23 : _GEN_3274; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3276 = 14'h18 == parameter_2_41 ? phv_data_24 : _GEN_3275; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3277 = 14'h19 == parameter_2_41 ? phv_data_25 : _GEN_3276; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3278 = 14'h1a == parameter_2_41 ? phv_data_26 : _GEN_3277; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3279 = 14'h1b == parameter_2_41 ? phv_data_27 : _GEN_3278; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3280 = 14'h1c == parameter_2_41 ? phv_data_28 : _GEN_3279; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3281 = 14'h1d == parameter_2_41 ? phv_data_29 : _GEN_3280; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3282 = 14'h1e == parameter_2_41 ? phv_data_30 : _GEN_3281; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3283 = 14'h1f == parameter_2_41 ? phv_data_31 : _GEN_3282; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3284 = 14'h20 == parameter_2_41 ? phv_data_32 : _GEN_3283; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3285 = 14'h21 == parameter_2_41 ? phv_data_33 : _GEN_3284; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3286 = 14'h22 == parameter_2_41 ? phv_data_34 : _GEN_3285; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3287 = 14'h23 == parameter_2_41 ? phv_data_35 : _GEN_3286; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3288 = 14'h24 == parameter_2_41 ? phv_data_36 : _GEN_3287; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3289 = 14'h25 == parameter_2_41 ? phv_data_37 : _GEN_3288; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3290 = 14'h26 == parameter_2_41 ? phv_data_38 : _GEN_3289; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3291 = 14'h27 == parameter_2_41 ? phv_data_39 : _GEN_3290; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3292 = 14'h28 == parameter_2_41 ? phv_data_40 : _GEN_3291; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3293 = 14'h29 == parameter_2_41 ? phv_data_41 : _GEN_3292; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3294 = 14'h2a == parameter_2_41 ? phv_data_42 : _GEN_3293; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3295 = 14'h2b == parameter_2_41 ? phv_data_43 : _GEN_3294; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3296 = 14'h2c == parameter_2_41 ? phv_data_44 : _GEN_3295; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3297 = 14'h2d == parameter_2_41 ? phv_data_45 : _GEN_3296; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3298 = 14'h2e == parameter_2_41 ? phv_data_46 : _GEN_3297; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3299 = 14'h2f == parameter_2_41 ? phv_data_47 : _GEN_3298; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3300 = 14'h30 == parameter_2_41 ? phv_data_48 : _GEN_3299; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3301 = 14'h31 == parameter_2_41 ? phv_data_49 : _GEN_3300; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3302 = 14'h32 == parameter_2_41 ? phv_data_50 : _GEN_3301; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3303 = 14'h33 == parameter_2_41 ? phv_data_51 : _GEN_3302; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3304 = 14'h34 == parameter_2_41 ? phv_data_52 : _GEN_3303; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3305 = 14'h35 == parameter_2_41 ? phv_data_53 : _GEN_3304; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3306 = 14'h36 == parameter_2_41 ? phv_data_54 : _GEN_3305; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3307 = 14'h37 == parameter_2_41 ? phv_data_55 : _GEN_3306; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3308 = 14'h38 == parameter_2_41 ? phv_data_56 : _GEN_3307; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3309 = 14'h39 == parameter_2_41 ? phv_data_57 : _GEN_3308; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3310 = 14'h3a == parameter_2_41 ? phv_data_58 : _GEN_3309; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3311 = 14'h3b == parameter_2_41 ? phv_data_59 : _GEN_3310; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3312 = 14'h3c == parameter_2_41 ? phv_data_60 : _GEN_3311; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3313 = 14'h3d == parameter_2_41 ? phv_data_61 : _GEN_3312; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3314 = 14'h3e == parameter_2_41 ? phv_data_62 : _GEN_3313; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3315 = 14'h3f == parameter_2_41 ? phv_data_63 : _GEN_3314; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_42 = vliw_42[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_42 = vliw_42[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_42 = parameter_2_42[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_42 = parameter_2_42[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_42 = {{1'd0}, args_offset_42}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_42 = _total_offset_T_42[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3319 = 3'h1 == total_offset_42 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3320 = 3'h2 == total_offset_42 ? args_2 : _GEN_3319; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3321 = 3'h3 == total_offset_42 ? args_3 : _GEN_3320; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3322 = 3'h4 == total_offset_42 ? args_4 : _GEN_3321; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3323 = 3'h5 == total_offset_42 ? args_5 : _GEN_3322; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3324 = 3'h6 == total_offset_42 ? args_6 : _GEN_3323; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3325 = total_offset_42 < 3'h7 ? _GEN_3324 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_42_0 = 3'h0 < args_length_42 ? _GEN_3325 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_3327 = opcode_42 == 4'ha ? field_bytes_42_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3328 = opcode_42 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2985 = opcode_42 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_85 = _T_2985 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_3329 = opcode_42 == 4'h8 | opcode_42 == 4'hb ? parameter_2_42[7:0] : _GEN_3327; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_3330 = opcode_42 == 4'h8 | opcode_42 == 4'hb ? _field_tag_T_85 : _GEN_3328; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_3331 = 14'h0 == parameter_2_42 ? phv_data_0 : _GEN_3329; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3332 = 14'h1 == parameter_2_42 ? phv_data_1 : _GEN_3331; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3333 = 14'h2 == parameter_2_42 ? phv_data_2 : _GEN_3332; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3334 = 14'h3 == parameter_2_42 ? phv_data_3 : _GEN_3333; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3335 = 14'h4 == parameter_2_42 ? phv_data_4 : _GEN_3334; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3336 = 14'h5 == parameter_2_42 ? phv_data_5 : _GEN_3335; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3337 = 14'h6 == parameter_2_42 ? phv_data_6 : _GEN_3336; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3338 = 14'h7 == parameter_2_42 ? phv_data_7 : _GEN_3337; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3339 = 14'h8 == parameter_2_42 ? phv_data_8 : _GEN_3338; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3340 = 14'h9 == parameter_2_42 ? phv_data_9 : _GEN_3339; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3341 = 14'ha == parameter_2_42 ? phv_data_10 : _GEN_3340; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3342 = 14'hb == parameter_2_42 ? phv_data_11 : _GEN_3341; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3343 = 14'hc == parameter_2_42 ? phv_data_12 : _GEN_3342; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3344 = 14'hd == parameter_2_42 ? phv_data_13 : _GEN_3343; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3345 = 14'he == parameter_2_42 ? phv_data_14 : _GEN_3344; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3346 = 14'hf == parameter_2_42 ? phv_data_15 : _GEN_3345; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3347 = 14'h10 == parameter_2_42 ? phv_data_16 : _GEN_3346; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3348 = 14'h11 == parameter_2_42 ? phv_data_17 : _GEN_3347; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3349 = 14'h12 == parameter_2_42 ? phv_data_18 : _GEN_3348; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3350 = 14'h13 == parameter_2_42 ? phv_data_19 : _GEN_3349; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3351 = 14'h14 == parameter_2_42 ? phv_data_20 : _GEN_3350; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3352 = 14'h15 == parameter_2_42 ? phv_data_21 : _GEN_3351; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3353 = 14'h16 == parameter_2_42 ? phv_data_22 : _GEN_3352; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3354 = 14'h17 == parameter_2_42 ? phv_data_23 : _GEN_3353; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3355 = 14'h18 == parameter_2_42 ? phv_data_24 : _GEN_3354; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3356 = 14'h19 == parameter_2_42 ? phv_data_25 : _GEN_3355; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3357 = 14'h1a == parameter_2_42 ? phv_data_26 : _GEN_3356; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3358 = 14'h1b == parameter_2_42 ? phv_data_27 : _GEN_3357; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3359 = 14'h1c == parameter_2_42 ? phv_data_28 : _GEN_3358; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3360 = 14'h1d == parameter_2_42 ? phv_data_29 : _GEN_3359; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3361 = 14'h1e == parameter_2_42 ? phv_data_30 : _GEN_3360; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3362 = 14'h1f == parameter_2_42 ? phv_data_31 : _GEN_3361; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3363 = 14'h20 == parameter_2_42 ? phv_data_32 : _GEN_3362; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3364 = 14'h21 == parameter_2_42 ? phv_data_33 : _GEN_3363; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3365 = 14'h22 == parameter_2_42 ? phv_data_34 : _GEN_3364; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3366 = 14'h23 == parameter_2_42 ? phv_data_35 : _GEN_3365; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3367 = 14'h24 == parameter_2_42 ? phv_data_36 : _GEN_3366; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3368 = 14'h25 == parameter_2_42 ? phv_data_37 : _GEN_3367; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3369 = 14'h26 == parameter_2_42 ? phv_data_38 : _GEN_3368; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3370 = 14'h27 == parameter_2_42 ? phv_data_39 : _GEN_3369; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3371 = 14'h28 == parameter_2_42 ? phv_data_40 : _GEN_3370; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3372 = 14'h29 == parameter_2_42 ? phv_data_41 : _GEN_3371; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3373 = 14'h2a == parameter_2_42 ? phv_data_42 : _GEN_3372; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3374 = 14'h2b == parameter_2_42 ? phv_data_43 : _GEN_3373; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3375 = 14'h2c == parameter_2_42 ? phv_data_44 : _GEN_3374; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3376 = 14'h2d == parameter_2_42 ? phv_data_45 : _GEN_3375; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3377 = 14'h2e == parameter_2_42 ? phv_data_46 : _GEN_3376; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3378 = 14'h2f == parameter_2_42 ? phv_data_47 : _GEN_3377; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3379 = 14'h30 == parameter_2_42 ? phv_data_48 : _GEN_3378; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3380 = 14'h31 == parameter_2_42 ? phv_data_49 : _GEN_3379; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3381 = 14'h32 == parameter_2_42 ? phv_data_50 : _GEN_3380; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3382 = 14'h33 == parameter_2_42 ? phv_data_51 : _GEN_3381; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3383 = 14'h34 == parameter_2_42 ? phv_data_52 : _GEN_3382; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3384 = 14'h35 == parameter_2_42 ? phv_data_53 : _GEN_3383; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3385 = 14'h36 == parameter_2_42 ? phv_data_54 : _GEN_3384; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3386 = 14'h37 == parameter_2_42 ? phv_data_55 : _GEN_3385; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3387 = 14'h38 == parameter_2_42 ? phv_data_56 : _GEN_3386; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3388 = 14'h39 == parameter_2_42 ? phv_data_57 : _GEN_3387; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3389 = 14'h3a == parameter_2_42 ? phv_data_58 : _GEN_3388; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3390 = 14'h3b == parameter_2_42 ? phv_data_59 : _GEN_3389; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3391 = 14'h3c == parameter_2_42 ? phv_data_60 : _GEN_3390; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3392 = 14'h3d == parameter_2_42 ? phv_data_61 : _GEN_3391; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3393 = 14'h3e == parameter_2_42 ? phv_data_62 : _GEN_3392; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3394 = 14'h3f == parameter_2_42 ? phv_data_63 : _GEN_3393; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_43 = vliw_43[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_43 = vliw_43[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_43 = parameter_2_43[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_43 = parameter_2_43[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_43 = {{1'd0}, args_offset_43}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_43 = _total_offset_T_43[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3398 = 3'h1 == total_offset_43 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3399 = 3'h2 == total_offset_43 ? args_2 : _GEN_3398; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3400 = 3'h3 == total_offset_43 ? args_3 : _GEN_3399; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3401 = 3'h4 == total_offset_43 ? args_4 : _GEN_3400; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3402 = 3'h5 == total_offset_43 ? args_5 : _GEN_3401; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3403 = 3'h6 == total_offset_43 ? args_6 : _GEN_3402; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3404 = total_offset_43 < 3'h7 ? _GEN_3403 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_43_0 = 3'h0 < args_length_43 ? _GEN_3404 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_3406 = opcode_43 == 4'ha ? field_bytes_43_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3407 = opcode_43 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_3056 = opcode_43 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_87 = _T_3056 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_3408 = opcode_43 == 4'h8 | opcode_43 == 4'hb ? parameter_2_43[7:0] : _GEN_3406; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_3409 = opcode_43 == 4'h8 | opcode_43 == 4'hb ? _field_tag_T_87 : _GEN_3407; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_3410 = 14'h0 == parameter_2_43 ? phv_data_0 : _GEN_3408; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3411 = 14'h1 == parameter_2_43 ? phv_data_1 : _GEN_3410; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3412 = 14'h2 == parameter_2_43 ? phv_data_2 : _GEN_3411; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3413 = 14'h3 == parameter_2_43 ? phv_data_3 : _GEN_3412; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3414 = 14'h4 == parameter_2_43 ? phv_data_4 : _GEN_3413; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3415 = 14'h5 == parameter_2_43 ? phv_data_5 : _GEN_3414; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3416 = 14'h6 == parameter_2_43 ? phv_data_6 : _GEN_3415; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3417 = 14'h7 == parameter_2_43 ? phv_data_7 : _GEN_3416; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3418 = 14'h8 == parameter_2_43 ? phv_data_8 : _GEN_3417; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3419 = 14'h9 == parameter_2_43 ? phv_data_9 : _GEN_3418; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3420 = 14'ha == parameter_2_43 ? phv_data_10 : _GEN_3419; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3421 = 14'hb == parameter_2_43 ? phv_data_11 : _GEN_3420; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3422 = 14'hc == parameter_2_43 ? phv_data_12 : _GEN_3421; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3423 = 14'hd == parameter_2_43 ? phv_data_13 : _GEN_3422; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3424 = 14'he == parameter_2_43 ? phv_data_14 : _GEN_3423; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3425 = 14'hf == parameter_2_43 ? phv_data_15 : _GEN_3424; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3426 = 14'h10 == parameter_2_43 ? phv_data_16 : _GEN_3425; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3427 = 14'h11 == parameter_2_43 ? phv_data_17 : _GEN_3426; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3428 = 14'h12 == parameter_2_43 ? phv_data_18 : _GEN_3427; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3429 = 14'h13 == parameter_2_43 ? phv_data_19 : _GEN_3428; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3430 = 14'h14 == parameter_2_43 ? phv_data_20 : _GEN_3429; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3431 = 14'h15 == parameter_2_43 ? phv_data_21 : _GEN_3430; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3432 = 14'h16 == parameter_2_43 ? phv_data_22 : _GEN_3431; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3433 = 14'h17 == parameter_2_43 ? phv_data_23 : _GEN_3432; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3434 = 14'h18 == parameter_2_43 ? phv_data_24 : _GEN_3433; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3435 = 14'h19 == parameter_2_43 ? phv_data_25 : _GEN_3434; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3436 = 14'h1a == parameter_2_43 ? phv_data_26 : _GEN_3435; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3437 = 14'h1b == parameter_2_43 ? phv_data_27 : _GEN_3436; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3438 = 14'h1c == parameter_2_43 ? phv_data_28 : _GEN_3437; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3439 = 14'h1d == parameter_2_43 ? phv_data_29 : _GEN_3438; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3440 = 14'h1e == parameter_2_43 ? phv_data_30 : _GEN_3439; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3441 = 14'h1f == parameter_2_43 ? phv_data_31 : _GEN_3440; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3442 = 14'h20 == parameter_2_43 ? phv_data_32 : _GEN_3441; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3443 = 14'h21 == parameter_2_43 ? phv_data_33 : _GEN_3442; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3444 = 14'h22 == parameter_2_43 ? phv_data_34 : _GEN_3443; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3445 = 14'h23 == parameter_2_43 ? phv_data_35 : _GEN_3444; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3446 = 14'h24 == parameter_2_43 ? phv_data_36 : _GEN_3445; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3447 = 14'h25 == parameter_2_43 ? phv_data_37 : _GEN_3446; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3448 = 14'h26 == parameter_2_43 ? phv_data_38 : _GEN_3447; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3449 = 14'h27 == parameter_2_43 ? phv_data_39 : _GEN_3448; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3450 = 14'h28 == parameter_2_43 ? phv_data_40 : _GEN_3449; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3451 = 14'h29 == parameter_2_43 ? phv_data_41 : _GEN_3450; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3452 = 14'h2a == parameter_2_43 ? phv_data_42 : _GEN_3451; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3453 = 14'h2b == parameter_2_43 ? phv_data_43 : _GEN_3452; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3454 = 14'h2c == parameter_2_43 ? phv_data_44 : _GEN_3453; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3455 = 14'h2d == parameter_2_43 ? phv_data_45 : _GEN_3454; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3456 = 14'h2e == parameter_2_43 ? phv_data_46 : _GEN_3455; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3457 = 14'h2f == parameter_2_43 ? phv_data_47 : _GEN_3456; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3458 = 14'h30 == parameter_2_43 ? phv_data_48 : _GEN_3457; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3459 = 14'h31 == parameter_2_43 ? phv_data_49 : _GEN_3458; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3460 = 14'h32 == parameter_2_43 ? phv_data_50 : _GEN_3459; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3461 = 14'h33 == parameter_2_43 ? phv_data_51 : _GEN_3460; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3462 = 14'h34 == parameter_2_43 ? phv_data_52 : _GEN_3461; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3463 = 14'h35 == parameter_2_43 ? phv_data_53 : _GEN_3462; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3464 = 14'h36 == parameter_2_43 ? phv_data_54 : _GEN_3463; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3465 = 14'h37 == parameter_2_43 ? phv_data_55 : _GEN_3464; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3466 = 14'h38 == parameter_2_43 ? phv_data_56 : _GEN_3465; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3467 = 14'h39 == parameter_2_43 ? phv_data_57 : _GEN_3466; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3468 = 14'h3a == parameter_2_43 ? phv_data_58 : _GEN_3467; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3469 = 14'h3b == parameter_2_43 ? phv_data_59 : _GEN_3468; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3470 = 14'h3c == parameter_2_43 ? phv_data_60 : _GEN_3469; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3471 = 14'h3d == parameter_2_43 ? phv_data_61 : _GEN_3470; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3472 = 14'h3e == parameter_2_43 ? phv_data_62 : _GEN_3471; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3473 = 14'h3f == parameter_2_43 ? phv_data_63 : _GEN_3472; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_44 = vliw_44[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_44 = vliw_44[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_44 = parameter_2_44[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_44 = parameter_2_44[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_44 = {{1'd0}, args_offset_44}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_44 = _total_offset_T_44[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3477 = 3'h1 == total_offset_44 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3478 = 3'h2 == total_offset_44 ? args_2 : _GEN_3477; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3479 = 3'h3 == total_offset_44 ? args_3 : _GEN_3478; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3480 = 3'h4 == total_offset_44 ? args_4 : _GEN_3479; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3481 = 3'h5 == total_offset_44 ? args_5 : _GEN_3480; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3482 = 3'h6 == total_offset_44 ? args_6 : _GEN_3481; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3483 = total_offset_44 < 3'h7 ? _GEN_3482 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_44_0 = 3'h0 < args_length_44 ? _GEN_3483 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_3485 = opcode_44 == 4'ha ? field_bytes_44_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3486 = opcode_44 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_3127 = opcode_44 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_89 = _T_3127 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_3487 = opcode_44 == 4'h8 | opcode_44 == 4'hb ? parameter_2_44[7:0] : _GEN_3485; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_3488 = opcode_44 == 4'h8 | opcode_44 == 4'hb ? _field_tag_T_89 : _GEN_3486; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_3489 = 14'h0 == parameter_2_44 ? phv_data_0 : _GEN_3487; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3490 = 14'h1 == parameter_2_44 ? phv_data_1 : _GEN_3489; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3491 = 14'h2 == parameter_2_44 ? phv_data_2 : _GEN_3490; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3492 = 14'h3 == parameter_2_44 ? phv_data_3 : _GEN_3491; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3493 = 14'h4 == parameter_2_44 ? phv_data_4 : _GEN_3492; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3494 = 14'h5 == parameter_2_44 ? phv_data_5 : _GEN_3493; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3495 = 14'h6 == parameter_2_44 ? phv_data_6 : _GEN_3494; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3496 = 14'h7 == parameter_2_44 ? phv_data_7 : _GEN_3495; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3497 = 14'h8 == parameter_2_44 ? phv_data_8 : _GEN_3496; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3498 = 14'h9 == parameter_2_44 ? phv_data_9 : _GEN_3497; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3499 = 14'ha == parameter_2_44 ? phv_data_10 : _GEN_3498; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3500 = 14'hb == parameter_2_44 ? phv_data_11 : _GEN_3499; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3501 = 14'hc == parameter_2_44 ? phv_data_12 : _GEN_3500; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3502 = 14'hd == parameter_2_44 ? phv_data_13 : _GEN_3501; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3503 = 14'he == parameter_2_44 ? phv_data_14 : _GEN_3502; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3504 = 14'hf == parameter_2_44 ? phv_data_15 : _GEN_3503; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3505 = 14'h10 == parameter_2_44 ? phv_data_16 : _GEN_3504; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3506 = 14'h11 == parameter_2_44 ? phv_data_17 : _GEN_3505; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3507 = 14'h12 == parameter_2_44 ? phv_data_18 : _GEN_3506; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3508 = 14'h13 == parameter_2_44 ? phv_data_19 : _GEN_3507; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3509 = 14'h14 == parameter_2_44 ? phv_data_20 : _GEN_3508; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3510 = 14'h15 == parameter_2_44 ? phv_data_21 : _GEN_3509; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3511 = 14'h16 == parameter_2_44 ? phv_data_22 : _GEN_3510; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3512 = 14'h17 == parameter_2_44 ? phv_data_23 : _GEN_3511; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3513 = 14'h18 == parameter_2_44 ? phv_data_24 : _GEN_3512; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3514 = 14'h19 == parameter_2_44 ? phv_data_25 : _GEN_3513; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3515 = 14'h1a == parameter_2_44 ? phv_data_26 : _GEN_3514; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3516 = 14'h1b == parameter_2_44 ? phv_data_27 : _GEN_3515; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3517 = 14'h1c == parameter_2_44 ? phv_data_28 : _GEN_3516; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3518 = 14'h1d == parameter_2_44 ? phv_data_29 : _GEN_3517; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3519 = 14'h1e == parameter_2_44 ? phv_data_30 : _GEN_3518; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3520 = 14'h1f == parameter_2_44 ? phv_data_31 : _GEN_3519; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3521 = 14'h20 == parameter_2_44 ? phv_data_32 : _GEN_3520; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3522 = 14'h21 == parameter_2_44 ? phv_data_33 : _GEN_3521; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3523 = 14'h22 == parameter_2_44 ? phv_data_34 : _GEN_3522; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3524 = 14'h23 == parameter_2_44 ? phv_data_35 : _GEN_3523; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3525 = 14'h24 == parameter_2_44 ? phv_data_36 : _GEN_3524; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3526 = 14'h25 == parameter_2_44 ? phv_data_37 : _GEN_3525; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3527 = 14'h26 == parameter_2_44 ? phv_data_38 : _GEN_3526; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3528 = 14'h27 == parameter_2_44 ? phv_data_39 : _GEN_3527; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3529 = 14'h28 == parameter_2_44 ? phv_data_40 : _GEN_3528; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3530 = 14'h29 == parameter_2_44 ? phv_data_41 : _GEN_3529; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3531 = 14'h2a == parameter_2_44 ? phv_data_42 : _GEN_3530; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3532 = 14'h2b == parameter_2_44 ? phv_data_43 : _GEN_3531; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3533 = 14'h2c == parameter_2_44 ? phv_data_44 : _GEN_3532; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3534 = 14'h2d == parameter_2_44 ? phv_data_45 : _GEN_3533; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3535 = 14'h2e == parameter_2_44 ? phv_data_46 : _GEN_3534; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3536 = 14'h2f == parameter_2_44 ? phv_data_47 : _GEN_3535; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3537 = 14'h30 == parameter_2_44 ? phv_data_48 : _GEN_3536; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3538 = 14'h31 == parameter_2_44 ? phv_data_49 : _GEN_3537; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3539 = 14'h32 == parameter_2_44 ? phv_data_50 : _GEN_3538; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3540 = 14'h33 == parameter_2_44 ? phv_data_51 : _GEN_3539; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3541 = 14'h34 == parameter_2_44 ? phv_data_52 : _GEN_3540; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3542 = 14'h35 == parameter_2_44 ? phv_data_53 : _GEN_3541; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3543 = 14'h36 == parameter_2_44 ? phv_data_54 : _GEN_3542; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3544 = 14'h37 == parameter_2_44 ? phv_data_55 : _GEN_3543; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3545 = 14'h38 == parameter_2_44 ? phv_data_56 : _GEN_3544; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3546 = 14'h39 == parameter_2_44 ? phv_data_57 : _GEN_3545; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3547 = 14'h3a == parameter_2_44 ? phv_data_58 : _GEN_3546; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3548 = 14'h3b == parameter_2_44 ? phv_data_59 : _GEN_3547; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3549 = 14'h3c == parameter_2_44 ? phv_data_60 : _GEN_3548; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3550 = 14'h3d == parameter_2_44 ? phv_data_61 : _GEN_3549; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3551 = 14'h3e == parameter_2_44 ? phv_data_62 : _GEN_3550; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3552 = 14'h3f == parameter_2_44 ? phv_data_63 : _GEN_3551; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_45 = vliw_45[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_45 = vliw_45[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_45 = parameter_2_45[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_45 = parameter_2_45[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_45 = {{1'd0}, args_offset_45}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_45 = _total_offset_T_45[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3556 = 3'h1 == total_offset_45 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3557 = 3'h2 == total_offset_45 ? args_2 : _GEN_3556; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3558 = 3'h3 == total_offset_45 ? args_3 : _GEN_3557; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3559 = 3'h4 == total_offset_45 ? args_4 : _GEN_3558; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3560 = 3'h5 == total_offset_45 ? args_5 : _GEN_3559; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3561 = 3'h6 == total_offset_45 ? args_6 : _GEN_3560; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3562 = total_offset_45 < 3'h7 ? _GEN_3561 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_45_0 = 3'h0 < args_length_45 ? _GEN_3562 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_3564 = opcode_45 == 4'ha ? field_bytes_45_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3565 = opcode_45 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_3198 = opcode_45 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_91 = _T_3198 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_3566 = opcode_45 == 4'h8 | opcode_45 == 4'hb ? parameter_2_45[7:0] : _GEN_3564; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_3567 = opcode_45 == 4'h8 | opcode_45 == 4'hb ? _field_tag_T_91 : _GEN_3565; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_3568 = 14'h0 == parameter_2_45 ? phv_data_0 : _GEN_3566; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3569 = 14'h1 == parameter_2_45 ? phv_data_1 : _GEN_3568; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3570 = 14'h2 == parameter_2_45 ? phv_data_2 : _GEN_3569; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3571 = 14'h3 == parameter_2_45 ? phv_data_3 : _GEN_3570; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3572 = 14'h4 == parameter_2_45 ? phv_data_4 : _GEN_3571; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3573 = 14'h5 == parameter_2_45 ? phv_data_5 : _GEN_3572; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3574 = 14'h6 == parameter_2_45 ? phv_data_6 : _GEN_3573; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3575 = 14'h7 == parameter_2_45 ? phv_data_7 : _GEN_3574; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3576 = 14'h8 == parameter_2_45 ? phv_data_8 : _GEN_3575; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3577 = 14'h9 == parameter_2_45 ? phv_data_9 : _GEN_3576; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3578 = 14'ha == parameter_2_45 ? phv_data_10 : _GEN_3577; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3579 = 14'hb == parameter_2_45 ? phv_data_11 : _GEN_3578; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3580 = 14'hc == parameter_2_45 ? phv_data_12 : _GEN_3579; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3581 = 14'hd == parameter_2_45 ? phv_data_13 : _GEN_3580; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3582 = 14'he == parameter_2_45 ? phv_data_14 : _GEN_3581; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3583 = 14'hf == parameter_2_45 ? phv_data_15 : _GEN_3582; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3584 = 14'h10 == parameter_2_45 ? phv_data_16 : _GEN_3583; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3585 = 14'h11 == parameter_2_45 ? phv_data_17 : _GEN_3584; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3586 = 14'h12 == parameter_2_45 ? phv_data_18 : _GEN_3585; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3587 = 14'h13 == parameter_2_45 ? phv_data_19 : _GEN_3586; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3588 = 14'h14 == parameter_2_45 ? phv_data_20 : _GEN_3587; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3589 = 14'h15 == parameter_2_45 ? phv_data_21 : _GEN_3588; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3590 = 14'h16 == parameter_2_45 ? phv_data_22 : _GEN_3589; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3591 = 14'h17 == parameter_2_45 ? phv_data_23 : _GEN_3590; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3592 = 14'h18 == parameter_2_45 ? phv_data_24 : _GEN_3591; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3593 = 14'h19 == parameter_2_45 ? phv_data_25 : _GEN_3592; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3594 = 14'h1a == parameter_2_45 ? phv_data_26 : _GEN_3593; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3595 = 14'h1b == parameter_2_45 ? phv_data_27 : _GEN_3594; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3596 = 14'h1c == parameter_2_45 ? phv_data_28 : _GEN_3595; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3597 = 14'h1d == parameter_2_45 ? phv_data_29 : _GEN_3596; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3598 = 14'h1e == parameter_2_45 ? phv_data_30 : _GEN_3597; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3599 = 14'h1f == parameter_2_45 ? phv_data_31 : _GEN_3598; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3600 = 14'h20 == parameter_2_45 ? phv_data_32 : _GEN_3599; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3601 = 14'h21 == parameter_2_45 ? phv_data_33 : _GEN_3600; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3602 = 14'h22 == parameter_2_45 ? phv_data_34 : _GEN_3601; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3603 = 14'h23 == parameter_2_45 ? phv_data_35 : _GEN_3602; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3604 = 14'h24 == parameter_2_45 ? phv_data_36 : _GEN_3603; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3605 = 14'h25 == parameter_2_45 ? phv_data_37 : _GEN_3604; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3606 = 14'h26 == parameter_2_45 ? phv_data_38 : _GEN_3605; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3607 = 14'h27 == parameter_2_45 ? phv_data_39 : _GEN_3606; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3608 = 14'h28 == parameter_2_45 ? phv_data_40 : _GEN_3607; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3609 = 14'h29 == parameter_2_45 ? phv_data_41 : _GEN_3608; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3610 = 14'h2a == parameter_2_45 ? phv_data_42 : _GEN_3609; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3611 = 14'h2b == parameter_2_45 ? phv_data_43 : _GEN_3610; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3612 = 14'h2c == parameter_2_45 ? phv_data_44 : _GEN_3611; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3613 = 14'h2d == parameter_2_45 ? phv_data_45 : _GEN_3612; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3614 = 14'h2e == parameter_2_45 ? phv_data_46 : _GEN_3613; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3615 = 14'h2f == parameter_2_45 ? phv_data_47 : _GEN_3614; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3616 = 14'h30 == parameter_2_45 ? phv_data_48 : _GEN_3615; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3617 = 14'h31 == parameter_2_45 ? phv_data_49 : _GEN_3616; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3618 = 14'h32 == parameter_2_45 ? phv_data_50 : _GEN_3617; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3619 = 14'h33 == parameter_2_45 ? phv_data_51 : _GEN_3618; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3620 = 14'h34 == parameter_2_45 ? phv_data_52 : _GEN_3619; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3621 = 14'h35 == parameter_2_45 ? phv_data_53 : _GEN_3620; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3622 = 14'h36 == parameter_2_45 ? phv_data_54 : _GEN_3621; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3623 = 14'h37 == parameter_2_45 ? phv_data_55 : _GEN_3622; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3624 = 14'h38 == parameter_2_45 ? phv_data_56 : _GEN_3623; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3625 = 14'h39 == parameter_2_45 ? phv_data_57 : _GEN_3624; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3626 = 14'h3a == parameter_2_45 ? phv_data_58 : _GEN_3625; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3627 = 14'h3b == parameter_2_45 ? phv_data_59 : _GEN_3626; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3628 = 14'h3c == parameter_2_45 ? phv_data_60 : _GEN_3627; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3629 = 14'h3d == parameter_2_45 ? phv_data_61 : _GEN_3628; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3630 = 14'h3e == parameter_2_45 ? phv_data_62 : _GEN_3629; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3631 = 14'h3f == parameter_2_45 ? phv_data_63 : _GEN_3630; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_46 = vliw_46[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_46 = vliw_46[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_46 = parameter_2_46[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_46 = parameter_2_46[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_46 = {{1'd0}, args_offset_46}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_46 = _total_offset_T_46[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3635 = 3'h1 == total_offset_46 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3636 = 3'h2 == total_offset_46 ? args_2 : _GEN_3635; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3637 = 3'h3 == total_offset_46 ? args_3 : _GEN_3636; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3638 = 3'h4 == total_offset_46 ? args_4 : _GEN_3637; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3639 = 3'h5 == total_offset_46 ? args_5 : _GEN_3638; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3640 = 3'h6 == total_offset_46 ? args_6 : _GEN_3639; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3641 = total_offset_46 < 3'h7 ? _GEN_3640 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_46_0 = 3'h0 < args_length_46 ? _GEN_3641 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_3643 = opcode_46 == 4'ha ? field_bytes_46_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3644 = opcode_46 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_3269 = opcode_46 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_93 = _T_3269 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_3645 = opcode_46 == 4'h8 | opcode_46 == 4'hb ? parameter_2_46[7:0] : _GEN_3643; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_3646 = opcode_46 == 4'h8 | opcode_46 == 4'hb ? _field_tag_T_93 : _GEN_3644; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_3647 = 14'h0 == parameter_2_46 ? phv_data_0 : _GEN_3645; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3648 = 14'h1 == parameter_2_46 ? phv_data_1 : _GEN_3647; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3649 = 14'h2 == parameter_2_46 ? phv_data_2 : _GEN_3648; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3650 = 14'h3 == parameter_2_46 ? phv_data_3 : _GEN_3649; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3651 = 14'h4 == parameter_2_46 ? phv_data_4 : _GEN_3650; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3652 = 14'h5 == parameter_2_46 ? phv_data_5 : _GEN_3651; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3653 = 14'h6 == parameter_2_46 ? phv_data_6 : _GEN_3652; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3654 = 14'h7 == parameter_2_46 ? phv_data_7 : _GEN_3653; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3655 = 14'h8 == parameter_2_46 ? phv_data_8 : _GEN_3654; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3656 = 14'h9 == parameter_2_46 ? phv_data_9 : _GEN_3655; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3657 = 14'ha == parameter_2_46 ? phv_data_10 : _GEN_3656; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3658 = 14'hb == parameter_2_46 ? phv_data_11 : _GEN_3657; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3659 = 14'hc == parameter_2_46 ? phv_data_12 : _GEN_3658; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3660 = 14'hd == parameter_2_46 ? phv_data_13 : _GEN_3659; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3661 = 14'he == parameter_2_46 ? phv_data_14 : _GEN_3660; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3662 = 14'hf == parameter_2_46 ? phv_data_15 : _GEN_3661; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3663 = 14'h10 == parameter_2_46 ? phv_data_16 : _GEN_3662; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3664 = 14'h11 == parameter_2_46 ? phv_data_17 : _GEN_3663; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3665 = 14'h12 == parameter_2_46 ? phv_data_18 : _GEN_3664; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3666 = 14'h13 == parameter_2_46 ? phv_data_19 : _GEN_3665; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3667 = 14'h14 == parameter_2_46 ? phv_data_20 : _GEN_3666; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3668 = 14'h15 == parameter_2_46 ? phv_data_21 : _GEN_3667; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3669 = 14'h16 == parameter_2_46 ? phv_data_22 : _GEN_3668; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3670 = 14'h17 == parameter_2_46 ? phv_data_23 : _GEN_3669; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3671 = 14'h18 == parameter_2_46 ? phv_data_24 : _GEN_3670; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3672 = 14'h19 == parameter_2_46 ? phv_data_25 : _GEN_3671; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3673 = 14'h1a == parameter_2_46 ? phv_data_26 : _GEN_3672; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3674 = 14'h1b == parameter_2_46 ? phv_data_27 : _GEN_3673; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3675 = 14'h1c == parameter_2_46 ? phv_data_28 : _GEN_3674; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3676 = 14'h1d == parameter_2_46 ? phv_data_29 : _GEN_3675; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3677 = 14'h1e == parameter_2_46 ? phv_data_30 : _GEN_3676; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3678 = 14'h1f == parameter_2_46 ? phv_data_31 : _GEN_3677; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3679 = 14'h20 == parameter_2_46 ? phv_data_32 : _GEN_3678; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3680 = 14'h21 == parameter_2_46 ? phv_data_33 : _GEN_3679; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3681 = 14'h22 == parameter_2_46 ? phv_data_34 : _GEN_3680; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3682 = 14'h23 == parameter_2_46 ? phv_data_35 : _GEN_3681; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3683 = 14'h24 == parameter_2_46 ? phv_data_36 : _GEN_3682; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3684 = 14'h25 == parameter_2_46 ? phv_data_37 : _GEN_3683; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3685 = 14'h26 == parameter_2_46 ? phv_data_38 : _GEN_3684; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3686 = 14'h27 == parameter_2_46 ? phv_data_39 : _GEN_3685; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3687 = 14'h28 == parameter_2_46 ? phv_data_40 : _GEN_3686; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3688 = 14'h29 == parameter_2_46 ? phv_data_41 : _GEN_3687; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3689 = 14'h2a == parameter_2_46 ? phv_data_42 : _GEN_3688; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3690 = 14'h2b == parameter_2_46 ? phv_data_43 : _GEN_3689; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3691 = 14'h2c == parameter_2_46 ? phv_data_44 : _GEN_3690; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3692 = 14'h2d == parameter_2_46 ? phv_data_45 : _GEN_3691; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3693 = 14'h2e == parameter_2_46 ? phv_data_46 : _GEN_3692; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3694 = 14'h2f == parameter_2_46 ? phv_data_47 : _GEN_3693; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3695 = 14'h30 == parameter_2_46 ? phv_data_48 : _GEN_3694; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3696 = 14'h31 == parameter_2_46 ? phv_data_49 : _GEN_3695; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3697 = 14'h32 == parameter_2_46 ? phv_data_50 : _GEN_3696; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3698 = 14'h33 == parameter_2_46 ? phv_data_51 : _GEN_3697; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3699 = 14'h34 == parameter_2_46 ? phv_data_52 : _GEN_3698; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3700 = 14'h35 == parameter_2_46 ? phv_data_53 : _GEN_3699; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3701 = 14'h36 == parameter_2_46 ? phv_data_54 : _GEN_3700; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3702 = 14'h37 == parameter_2_46 ? phv_data_55 : _GEN_3701; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3703 = 14'h38 == parameter_2_46 ? phv_data_56 : _GEN_3702; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3704 = 14'h39 == parameter_2_46 ? phv_data_57 : _GEN_3703; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3705 = 14'h3a == parameter_2_46 ? phv_data_58 : _GEN_3704; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3706 = 14'h3b == parameter_2_46 ? phv_data_59 : _GEN_3705; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3707 = 14'h3c == parameter_2_46 ? phv_data_60 : _GEN_3706; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3708 = 14'h3d == parameter_2_46 ? phv_data_61 : _GEN_3707; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3709 = 14'h3e == parameter_2_46 ? phv_data_62 : _GEN_3708; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3710 = 14'h3f == parameter_2_46 ? phv_data_63 : _GEN_3709; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_47 = vliw_47[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_47 = vliw_47[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_47 = parameter_2_47[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_47 = parameter_2_47[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_47 = {{1'd0}, args_offset_47}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_47 = _total_offset_T_47[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3714 = 3'h1 == total_offset_47 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3715 = 3'h2 == total_offset_47 ? args_2 : _GEN_3714; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3716 = 3'h3 == total_offset_47 ? args_3 : _GEN_3715; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3717 = 3'h4 == total_offset_47 ? args_4 : _GEN_3716; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3718 = 3'h5 == total_offset_47 ? args_5 : _GEN_3717; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3719 = 3'h6 == total_offset_47 ? args_6 : _GEN_3718; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3720 = total_offset_47 < 3'h7 ? _GEN_3719 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_47_0 = 3'h0 < args_length_47 ? _GEN_3720 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_3722 = opcode_47 == 4'ha ? field_bytes_47_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3723 = opcode_47 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_3340 = opcode_47 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_95 = _T_3340 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_3724 = opcode_47 == 4'h8 | opcode_47 == 4'hb ? parameter_2_47[7:0] : _GEN_3722; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_3725 = opcode_47 == 4'h8 | opcode_47 == 4'hb ? _field_tag_T_95 : _GEN_3723; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_3726 = 14'h0 == parameter_2_47 ? phv_data_0 : _GEN_3724; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3727 = 14'h1 == parameter_2_47 ? phv_data_1 : _GEN_3726; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3728 = 14'h2 == parameter_2_47 ? phv_data_2 : _GEN_3727; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3729 = 14'h3 == parameter_2_47 ? phv_data_3 : _GEN_3728; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3730 = 14'h4 == parameter_2_47 ? phv_data_4 : _GEN_3729; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3731 = 14'h5 == parameter_2_47 ? phv_data_5 : _GEN_3730; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3732 = 14'h6 == parameter_2_47 ? phv_data_6 : _GEN_3731; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3733 = 14'h7 == parameter_2_47 ? phv_data_7 : _GEN_3732; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3734 = 14'h8 == parameter_2_47 ? phv_data_8 : _GEN_3733; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3735 = 14'h9 == parameter_2_47 ? phv_data_9 : _GEN_3734; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3736 = 14'ha == parameter_2_47 ? phv_data_10 : _GEN_3735; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3737 = 14'hb == parameter_2_47 ? phv_data_11 : _GEN_3736; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3738 = 14'hc == parameter_2_47 ? phv_data_12 : _GEN_3737; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3739 = 14'hd == parameter_2_47 ? phv_data_13 : _GEN_3738; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3740 = 14'he == parameter_2_47 ? phv_data_14 : _GEN_3739; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3741 = 14'hf == parameter_2_47 ? phv_data_15 : _GEN_3740; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3742 = 14'h10 == parameter_2_47 ? phv_data_16 : _GEN_3741; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3743 = 14'h11 == parameter_2_47 ? phv_data_17 : _GEN_3742; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3744 = 14'h12 == parameter_2_47 ? phv_data_18 : _GEN_3743; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3745 = 14'h13 == parameter_2_47 ? phv_data_19 : _GEN_3744; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3746 = 14'h14 == parameter_2_47 ? phv_data_20 : _GEN_3745; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3747 = 14'h15 == parameter_2_47 ? phv_data_21 : _GEN_3746; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3748 = 14'h16 == parameter_2_47 ? phv_data_22 : _GEN_3747; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3749 = 14'h17 == parameter_2_47 ? phv_data_23 : _GEN_3748; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3750 = 14'h18 == parameter_2_47 ? phv_data_24 : _GEN_3749; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3751 = 14'h19 == parameter_2_47 ? phv_data_25 : _GEN_3750; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3752 = 14'h1a == parameter_2_47 ? phv_data_26 : _GEN_3751; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3753 = 14'h1b == parameter_2_47 ? phv_data_27 : _GEN_3752; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3754 = 14'h1c == parameter_2_47 ? phv_data_28 : _GEN_3753; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3755 = 14'h1d == parameter_2_47 ? phv_data_29 : _GEN_3754; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3756 = 14'h1e == parameter_2_47 ? phv_data_30 : _GEN_3755; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3757 = 14'h1f == parameter_2_47 ? phv_data_31 : _GEN_3756; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3758 = 14'h20 == parameter_2_47 ? phv_data_32 : _GEN_3757; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3759 = 14'h21 == parameter_2_47 ? phv_data_33 : _GEN_3758; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3760 = 14'h22 == parameter_2_47 ? phv_data_34 : _GEN_3759; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3761 = 14'h23 == parameter_2_47 ? phv_data_35 : _GEN_3760; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3762 = 14'h24 == parameter_2_47 ? phv_data_36 : _GEN_3761; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3763 = 14'h25 == parameter_2_47 ? phv_data_37 : _GEN_3762; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3764 = 14'h26 == parameter_2_47 ? phv_data_38 : _GEN_3763; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3765 = 14'h27 == parameter_2_47 ? phv_data_39 : _GEN_3764; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3766 = 14'h28 == parameter_2_47 ? phv_data_40 : _GEN_3765; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3767 = 14'h29 == parameter_2_47 ? phv_data_41 : _GEN_3766; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3768 = 14'h2a == parameter_2_47 ? phv_data_42 : _GEN_3767; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3769 = 14'h2b == parameter_2_47 ? phv_data_43 : _GEN_3768; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3770 = 14'h2c == parameter_2_47 ? phv_data_44 : _GEN_3769; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3771 = 14'h2d == parameter_2_47 ? phv_data_45 : _GEN_3770; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3772 = 14'h2e == parameter_2_47 ? phv_data_46 : _GEN_3771; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3773 = 14'h2f == parameter_2_47 ? phv_data_47 : _GEN_3772; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3774 = 14'h30 == parameter_2_47 ? phv_data_48 : _GEN_3773; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3775 = 14'h31 == parameter_2_47 ? phv_data_49 : _GEN_3774; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3776 = 14'h32 == parameter_2_47 ? phv_data_50 : _GEN_3775; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3777 = 14'h33 == parameter_2_47 ? phv_data_51 : _GEN_3776; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3778 = 14'h34 == parameter_2_47 ? phv_data_52 : _GEN_3777; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3779 = 14'h35 == parameter_2_47 ? phv_data_53 : _GEN_3778; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3780 = 14'h36 == parameter_2_47 ? phv_data_54 : _GEN_3779; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3781 = 14'h37 == parameter_2_47 ? phv_data_55 : _GEN_3780; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3782 = 14'h38 == parameter_2_47 ? phv_data_56 : _GEN_3781; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3783 = 14'h39 == parameter_2_47 ? phv_data_57 : _GEN_3782; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3784 = 14'h3a == parameter_2_47 ? phv_data_58 : _GEN_3783; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3785 = 14'h3b == parameter_2_47 ? phv_data_59 : _GEN_3784; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3786 = 14'h3c == parameter_2_47 ? phv_data_60 : _GEN_3785; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3787 = 14'h3d == parameter_2_47 ? phv_data_61 : _GEN_3786; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3788 = 14'h3e == parameter_2_47 ? phv_data_62 : _GEN_3787; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3789 = 14'h3f == parameter_2_47 ? phv_data_63 : _GEN_3788; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_48 = vliw_48[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_48 = vliw_48[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_48 = parameter_2_48[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_48 = parameter_2_48[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_48 = {{1'd0}, args_offset_48}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_48 = _total_offset_T_48[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3793 = 3'h1 == total_offset_48 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3794 = 3'h2 == total_offset_48 ? args_2 : _GEN_3793; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3795 = 3'h3 == total_offset_48 ? args_3 : _GEN_3794; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3796 = 3'h4 == total_offset_48 ? args_4 : _GEN_3795; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3797 = 3'h5 == total_offset_48 ? args_5 : _GEN_3796; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3798 = 3'h6 == total_offset_48 ? args_6 : _GEN_3797; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3799 = total_offset_48 < 3'h7 ? _GEN_3798 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_48_0 = 3'h0 < args_length_48 ? _GEN_3799 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_3801 = opcode_48 == 4'ha ? field_bytes_48_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3802 = opcode_48 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_3411 = opcode_48 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_97 = _T_3411 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_3803 = opcode_48 == 4'h8 | opcode_48 == 4'hb ? parameter_2_48[7:0] : _GEN_3801; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_3804 = opcode_48 == 4'h8 | opcode_48 == 4'hb ? _field_tag_T_97 : _GEN_3802; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_3805 = 14'h0 == parameter_2_48 ? phv_data_0 : _GEN_3803; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3806 = 14'h1 == parameter_2_48 ? phv_data_1 : _GEN_3805; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3807 = 14'h2 == parameter_2_48 ? phv_data_2 : _GEN_3806; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3808 = 14'h3 == parameter_2_48 ? phv_data_3 : _GEN_3807; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3809 = 14'h4 == parameter_2_48 ? phv_data_4 : _GEN_3808; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3810 = 14'h5 == parameter_2_48 ? phv_data_5 : _GEN_3809; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3811 = 14'h6 == parameter_2_48 ? phv_data_6 : _GEN_3810; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3812 = 14'h7 == parameter_2_48 ? phv_data_7 : _GEN_3811; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3813 = 14'h8 == parameter_2_48 ? phv_data_8 : _GEN_3812; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3814 = 14'h9 == parameter_2_48 ? phv_data_9 : _GEN_3813; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3815 = 14'ha == parameter_2_48 ? phv_data_10 : _GEN_3814; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3816 = 14'hb == parameter_2_48 ? phv_data_11 : _GEN_3815; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3817 = 14'hc == parameter_2_48 ? phv_data_12 : _GEN_3816; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3818 = 14'hd == parameter_2_48 ? phv_data_13 : _GEN_3817; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3819 = 14'he == parameter_2_48 ? phv_data_14 : _GEN_3818; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3820 = 14'hf == parameter_2_48 ? phv_data_15 : _GEN_3819; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3821 = 14'h10 == parameter_2_48 ? phv_data_16 : _GEN_3820; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3822 = 14'h11 == parameter_2_48 ? phv_data_17 : _GEN_3821; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3823 = 14'h12 == parameter_2_48 ? phv_data_18 : _GEN_3822; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3824 = 14'h13 == parameter_2_48 ? phv_data_19 : _GEN_3823; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3825 = 14'h14 == parameter_2_48 ? phv_data_20 : _GEN_3824; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3826 = 14'h15 == parameter_2_48 ? phv_data_21 : _GEN_3825; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3827 = 14'h16 == parameter_2_48 ? phv_data_22 : _GEN_3826; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3828 = 14'h17 == parameter_2_48 ? phv_data_23 : _GEN_3827; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3829 = 14'h18 == parameter_2_48 ? phv_data_24 : _GEN_3828; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3830 = 14'h19 == parameter_2_48 ? phv_data_25 : _GEN_3829; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3831 = 14'h1a == parameter_2_48 ? phv_data_26 : _GEN_3830; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3832 = 14'h1b == parameter_2_48 ? phv_data_27 : _GEN_3831; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3833 = 14'h1c == parameter_2_48 ? phv_data_28 : _GEN_3832; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3834 = 14'h1d == parameter_2_48 ? phv_data_29 : _GEN_3833; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3835 = 14'h1e == parameter_2_48 ? phv_data_30 : _GEN_3834; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3836 = 14'h1f == parameter_2_48 ? phv_data_31 : _GEN_3835; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3837 = 14'h20 == parameter_2_48 ? phv_data_32 : _GEN_3836; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3838 = 14'h21 == parameter_2_48 ? phv_data_33 : _GEN_3837; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3839 = 14'h22 == parameter_2_48 ? phv_data_34 : _GEN_3838; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3840 = 14'h23 == parameter_2_48 ? phv_data_35 : _GEN_3839; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3841 = 14'h24 == parameter_2_48 ? phv_data_36 : _GEN_3840; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3842 = 14'h25 == parameter_2_48 ? phv_data_37 : _GEN_3841; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3843 = 14'h26 == parameter_2_48 ? phv_data_38 : _GEN_3842; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3844 = 14'h27 == parameter_2_48 ? phv_data_39 : _GEN_3843; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3845 = 14'h28 == parameter_2_48 ? phv_data_40 : _GEN_3844; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3846 = 14'h29 == parameter_2_48 ? phv_data_41 : _GEN_3845; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3847 = 14'h2a == parameter_2_48 ? phv_data_42 : _GEN_3846; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3848 = 14'h2b == parameter_2_48 ? phv_data_43 : _GEN_3847; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3849 = 14'h2c == parameter_2_48 ? phv_data_44 : _GEN_3848; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3850 = 14'h2d == parameter_2_48 ? phv_data_45 : _GEN_3849; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3851 = 14'h2e == parameter_2_48 ? phv_data_46 : _GEN_3850; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3852 = 14'h2f == parameter_2_48 ? phv_data_47 : _GEN_3851; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3853 = 14'h30 == parameter_2_48 ? phv_data_48 : _GEN_3852; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3854 = 14'h31 == parameter_2_48 ? phv_data_49 : _GEN_3853; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3855 = 14'h32 == parameter_2_48 ? phv_data_50 : _GEN_3854; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3856 = 14'h33 == parameter_2_48 ? phv_data_51 : _GEN_3855; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3857 = 14'h34 == parameter_2_48 ? phv_data_52 : _GEN_3856; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3858 = 14'h35 == parameter_2_48 ? phv_data_53 : _GEN_3857; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3859 = 14'h36 == parameter_2_48 ? phv_data_54 : _GEN_3858; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3860 = 14'h37 == parameter_2_48 ? phv_data_55 : _GEN_3859; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3861 = 14'h38 == parameter_2_48 ? phv_data_56 : _GEN_3860; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3862 = 14'h39 == parameter_2_48 ? phv_data_57 : _GEN_3861; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3863 = 14'h3a == parameter_2_48 ? phv_data_58 : _GEN_3862; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3864 = 14'h3b == parameter_2_48 ? phv_data_59 : _GEN_3863; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3865 = 14'h3c == parameter_2_48 ? phv_data_60 : _GEN_3864; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3866 = 14'h3d == parameter_2_48 ? phv_data_61 : _GEN_3865; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3867 = 14'h3e == parameter_2_48 ? phv_data_62 : _GEN_3866; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3868 = 14'h3f == parameter_2_48 ? phv_data_63 : _GEN_3867; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_49 = vliw_49[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_49 = vliw_49[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_49 = parameter_2_49[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_49 = parameter_2_49[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_49 = {{1'd0}, args_offset_49}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_49 = _total_offset_T_49[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3872 = 3'h1 == total_offset_49 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3873 = 3'h2 == total_offset_49 ? args_2 : _GEN_3872; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3874 = 3'h3 == total_offset_49 ? args_3 : _GEN_3873; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3875 = 3'h4 == total_offset_49 ? args_4 : _GEN_3874; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3876 = 3'h5 == total_offset_49 ? args_5 : _GEN_3875; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3877 = 3'h6 == total_offset_49 ? args_6 : _GEN_3876; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3878 = total_offset_49 < 3'h7 ? _GEN_3877 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_49_0 = 3'h0 < args_length_49 ? _GEN_3878 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_3880 = opcode_49 == 4'ha ? field_bytes_49_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3881 = opcode_49 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_3482 = opcode_49 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_99 = _T_3482 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_3882 = opcode_49 == 4'h8 | opcode_49 == 4'hb ? parameter_2_49[7:0] : _GEN_3880; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_3883 = opcode_49 == 4'h8 | opcode_49 == 4'hb ? _field_tag_T_99 : _GEN_3881; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_3884 = 14'h0 == parameter_2_49 ? phv_data_0 : _GEN_3882; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3885 = 14'h1 == parameter_2_49 ? phv_data_1 : _GEN_3884; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3886 = 14'h2 == parameter_2_49 ? phv_data_2 : _GEN_3885; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3887 = 14'h3 == parameter_2_49 ? phv_data_3 : _GEN_3886; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3888 = 14'h4 == parameter_2_49 ? phv_data_4 : _GEN_3887; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3889 = 14'h5 == parameter_2_49 ? phv_data_5 : _GEN_3888; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3890 = 14'h6 == parameter_2_49 ? phv_data_6 : _GEN_3889; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3891 = 14'h7 == parameter_2_49 ? phv_data_7 : _GEN_3890; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3892 = 14'h8 == parameter_2_49 ? phv_data_8 : _GEN_3891; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3893 = 14'h9 == parameter_2_49 ? phv_data_9 : _GEN_3892; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3894 = 14'ha == parameter_2_49 ? phv_data_10 : _GEN_3893; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3895 = 14'hb == parameter_2_49 ? phv_data_11 : _GEN_3894; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3896 = 14'hc == parameter_2_49 ? phv_data_12 : _GEN_3895; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3897 = 14'hd == parameter_2_49 ? phv_data_13 : _GEN_3896; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3898 = 14'he == parameter_2_49 ? phv_data_14 : _GEN_3897; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3899 = 14'hf == parameter_2_49 ? phv_data_15 : _GEN_3898; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3900 = 14'h10 == parameter_2_49 ? phv_data_16 : _GEN_3899; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3901 = 14'h11 == parameter_2_49 ? phv_data_17 : _GEN_3900; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3902 = 14'h12 == parameter_2_49 ? phv_data_18 : _GEN_3901; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3903 = 14'h13 == parameter_2_49 ? phv_data_19 : _GEN_3902; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3904 = 14'h14 == parameter_2_49 ? phv_data_20 : _GEN_3903; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3905 = 14'h15 == parameter_2_49 ? phv_data_21 : _GEN_3904; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3906 = 14'h16 == parameter_2_49 ? phv_data_22 : _GEN_3905; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3907 = 14'h17 == parameter_2_49 ? phv_data_23 : _GEN_3906; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3908 = 14'h18 == parameter_2_49 ? phv_data_24 : _GEN_3907; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3909 = 14'h19 == parameter_2_49 ? phv_data_25 : _GEN_3908; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3910 = 14'h1a == parameter_2_49 ? phv_data_26 : _GEN_3909; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3911 = 14'h1b == parameter_2_49 ? phv_data_27 : _GEN_3910; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3912 = 14'h1c == parameter_2_49 ? phv_data_28 : _GEN_3911; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3913 = 14'h1d == parameter_2_49 ? phv_data_29 : _GEN_3912; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3914 = 14'h1e == parameter_2_49 ? phv_data_30 : _GEN_3913; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3915 = 14'h1f == parameter_2_49 ? phv_data_31 : _GEN_3914; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3916 = 14'h20 == parameter_2_49 ? phv_data_32 : _GEN_3915; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3917 = 14'h21 == parameter_2_49 ? phv_data_33 : _GEN_3916; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3918 = 14'h22 == parameter_2_49 ? phv_data_34 : _GEN_3917; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3919 = 14'h23 == parameter_2_49 ? phv_data_35 : _GEN_3918; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3920 = 14'h24 == parameter_2_49 ? phv_data_36 : _GEN_3919; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3921 = 14'h25 == parameter_2_49 ? phv_data_37 : _GEN_3920; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3922 = 14'h26 == parameter_2_49 ? phv_data_38 : _GEN_3921; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3923 = 14'h27 == parameter_2_49 ? phv_data_39 : _GEN_3922; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3924 = 14'h28 == parameter_2_49 ? phv_data_40 : _GEN_3923; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3925 = 14'h29 == parameter_2_49 ? phv_data_41 : _GEN_3924; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3926 = 14'h2a == parameter_2_49 ? phv_data_42 : _GEN_3925; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3927 = 14'h2b == parameter_2_49 ? phv_data_43 : _GEN_3926; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3928 = 14'h2c == parameter_2_49 ? phv_data_44 : _GEN_3927; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3929 = 14'h2d == parameter_2_49 ? phv_data_45 : _GEN_3928; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3930 = 14'h2e == parameter_2_49 ? phv_data_46 : _GEN_3929; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3931 = 14'h2f == parameter_2_49 ? phv_data_47 : _GEN_3930; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3932 = 14'h30 == parameter_2_49 ? phv_data_48 : _GEN_3931; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3933 = 14'h31 == parameter_2_49 ? phv_data_49 : _GEN_3932; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3934 = 14'h32 == parameter_2_49 ? phv_data_50 : _GEN_3933; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3935 = 14'h33 == parameter_2_49 ? phv_data_51 : _GEN_3934; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3936 = 14'h34 == parameter_2_49 ? phv_data_52 : _GEN_3935; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3937 = 14'h35 == parameter_2_49 ? phv_data_53 : _GEN_3936; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3938 = 14'h36 == parameter_2_49 ? phv_data_54 : _GEN_3937; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3939 = 14'h37 == parameter_2_49 ? phv_data_55 : _GEN_3938; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3940 = 14'h38 == parameter_2_49 ? phv_data_56 : _GEN_3939; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3941 = 14'h39 == parameter_2_49 ? phv_data_57 : _GEN_3940; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3942 = 14'h3a == parameter_2_49 ? phv_data_58 : _GEN_3941; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3943 = 14'h3b == parameter_2_49 ? phv_data_59 : _GEN_3942; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3944 = 14'h3c == parameter_2_49 ? phv_data_60 : _GEN_3943; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3945 = 14'h3d == parameter_2_49 ? phv_data_61 : _GEN_3944; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3946 = 14'h3e == parameter_2_49 ? phv_data_62 : _GEN_3945; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3947 = 14'h3f == parameter_2_49 ? phv_data_63 : _GEN_3946; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_50 = vliw_50[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_50 = vliw_50[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_50 = parameter_2_50[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_50 = parameter_2_50[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_50 = {{1'd0}, args_offset_50}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_50 = _total_offset_T_50[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3951 = 3'h1 == total_offset_50 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3952 = 3'h2 == total_offset_50 ? args_2 : _GEN_3951; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3953 = 3'h3 == total_offset_50 ? args_3 : _GEN_3952; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3954 = 3'h4 == total_offset_50 ? args_4 : _GEN_3953; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3955 = 3'h5 == total_offset_50 ? args_5 : _GEN_3954; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3956 = 3'h6 == total_offset_50 ? args_6 : _GEN_3955; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3957 = total_offset_50 < 3'h7 ? _GEN_3956 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_50_0 = 3'h0 < args_length_50 ? _GEN_3957 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_3959 = opcode_50 == 4'ha ? field_bytes_50_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3960 = opcode_50 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_3553 = opcode_50 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_101 = _T_3553 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_3961 = opcode_50 == 4'h8 | opcode_50 == 4'hb ? parameter_2_50[7:0] : _GEN_3959; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_3962 = opcode_50 == 4'h8 | opcode_50 == 4'hb ? _field_tag_T_101 : _GEN_3960; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_3963 = 14'h0 == parameter_2_50 ? phv_data_0 : _GEN_3961; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3964 = 14'h1 == parameter_2_50 ? phv_data_1 : _GEN_3963; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3965 = 14'h2 == parameter_2_50 ? phv_data_2 : _GEN_3964; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3966 = 14'h3 == parameter_2_50 ? phv_data_3 : _GEN_3965; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3967 = 14'h4 == parameter_2_50 ? phv_data_4 : _GEN_3966; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3968 = 14'h5 == parameter_2_50 ? phv_data_5 : _GEN_3967; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3969 = 14'h6 == parameter_2_50 ? phv_data_6 : _GEN_3968; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3970 = 14'h7 == parameter_2_50 ? phv_data_7 : _GEN_3969; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3971 = 14'h8 == parameter_2_50 ? phv_data_8 : _GEN_3970; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3972 = 14'h9 == parameter_2_50 ? phv_data_9 : _GEN_3971; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3973 = 14'ha == parameter_2_50 ? phv_data_10 : _GEN_3972; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3974 = 14'hb == parameter_2_50 ? phv_data_11 : _GEN_3973; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3975 = 14'hc == parameter_2_50 ? phv_data_12 : _GEN_3974; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3976 = 14'hd == parameter_2_50 ? phv_data_13 : _GEN_3975; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3977 = 14'he == parameter_2_50 ? phv_data_14 : _GEN_3976; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3978 = 14'hf == parameter_2_50 ? phv_data_15 : _GEN_3977; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3979 = 14'h10 == parameter_2_50 ? phv_data_16 : _GEN_3978; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3980 = 14'h11 == parameter_2_50 ? phv_data_17 : _GEN_3979; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3981 = 14'h12 == parameter_2_50 ? phv_data_18 : _GEN_3980; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3982 = 14'h13 == parameter_2_50 ? phv_data_19 : _GEN_3981; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3983 = 14'h14 == parameter_2_50 ? phv_data_20 : _GEN_3982; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3984 = 14'h15 == parameter_2_50 ? phv_data_21 : _GEN_3983; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3985 = 14'h16 == parameter_2_50 ? phv_data_22 : _GEN_3984; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3986 = 14'h17 == parameter_2_50 ? phv_data_23 : _GEN_3985; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3987 = 14'h18 == parameter_2_50 ? phv_data_24 : _GEN_3986; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3988 = 14'h19 == parameter_2_50 ? phv_data_25 : _GEN_3987; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3989 = 14'h1a == parameter_2_50 ? phv_data_26 : _GEN_3988; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3990 = 14'h1b == parameter_2_50 ? phv_data_27 : _GEN_3989; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3991 = 14'h1c == parameter_2_50 ? phv_data_28 : _GEN_3990; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3992 = 14'h1d == parameter_2_50 ? phv_data_29 : _GEN_3991; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3993 = 14'h1e == parameter_2_50 ? phv_data_30 : _GEN_3992; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3994 = 14'h1f == parameter_2_50 ? phv_data_31 : _GEN_3993; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3995 = 14'h20 == parameter_2_50 ? phv_data_32 : _GEN_3994; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3996 = 14'h21 == parameter_2_50 ? phv_data_33 : _GEN_3995; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3997 = 14'h22 == parameter_2_50 ? phv_data_34 : _GEN_3996; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3998 = 14'h23 == parameter_2_50 ? phv_data_35 : _GEN_3997; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_3999 = 14'h24 == parameter_2_50 ? phv_data_36 : _GEN_3998; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4000 = 14'h25 == parameter_2_50 ? phv_data_37 : _GEN_3999; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4001 = 14'h26 == parameter_2_50 ? phv_data_38 : _GEN_4000; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4002 = 14'h27 == parameter_2_50 ? phv_data_39 : _GEN_4001; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4003 = 14'h28 == parameter_2_50 ? phv_data_40 : _GEN_4002; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4004 = 14'h29 == parameter_2_50 ? phv_data_41 : _GEN_4003; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4005 = 14'h2a == parameter_2_50 ? phv_data_42 : _GEN_4004; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4006 = 14'h2b == parameter_2_50 ? phv_data_43 : _GEN_4005; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4007 = 14'h2c == parameter_2_50 ? phv_data_44 : _GEN_4006; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4008 = 14'h2d == parameter_2_50 ? phv_data_45 : _GEN_4007; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4009 = 14'h2e == parameter_2_50 ? phv_data_46 : _GEN_4008; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4010 = 14'h2f == parameter_2_50 ? phv_data_47 : _GEN_4009; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4011 = 14'h30 == parameter_2_50 ? phv_data_48 : _GEN_4010; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4012 = 14'h31 == parameter_2_50 ? phv_data_49 : _GEN_4011; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4013 = 14'h32 == parameter_2_50 ? phv_data_50 : _GEN_4012; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4014 = 14'h33 == parameter_2_50 ? phv_data_51 : _GEN_4013; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4015 = 14'h34 == parameter_2_50 ? phv_data_52 : _GEN_4014; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4016 = 14'h35 == parameter_2_50 ? phv_data_53 : _GEN_4015; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4017 = 14'h36 == parameter_2_50 ? phv_data_54 : _GEN_4016; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4018 = 14'h37 == parameter_2_50 ? phv_data_55 : _GEN_4017; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4019 = 14'h38 == parameter_2_50 ? phv_data_56 : _GEN_4018; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4020 = 14'h39 == parameter_2_50 ? phv_data_57 : _GEN_4019; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4021 = 14'h3a == parameter_2_50 ? phv_data_58 : _GEN_4020; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4022 = 14'h3b == parameter_2_50 ? phv_data_59 : _GEN_4021; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4023 = 14'h3c == parameter_2_50 ? phv_data_60 : _GEN_4022; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4024 = 14'h3d == parameter_2_50 ? phv_data_61 : _GEN_4023; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4025 = 14'h3e == parameter_2_50 ? phv_data_62 : _GEN_4024; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4026 = 14'h3f == parameter_2_50 ? phv_data_63 : _GEN_4025; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_51 = vliw_51[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_51 = vliw_51[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_51 = parameter_2_51[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_51 = parameter_2_51[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_51 = {{1'd0}, args_offset_51}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_51 = _total_offset_T_51[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_4030 = 3'h1 == total_offset_51 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4031 = 3'h2 == total_offset_51 ? args_2 : _GEN_4030; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4032 = 3'h3 == total_offset_51 ? args_3 : _GEN_4031; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4033 = 3'h4 == total_offset_51 ? args_4 : _GEN_4032; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4034 = 3'h5 == total_offset_51 ? args_5 : _GEN_4033; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4035 = 3'h6 == total_offset_51 ? args_6 : _GEN_4034; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4036 = total_offset_51 < 3'h7 ? _GEN_4035 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_51_0 = 3'h0 < args_length_51 ? _GEN_4036 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_4038 = opcode_51 == 4'ha ? field_bytes_51_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_4039 = opcode_51 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_3624 = opcode_51 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_103 = _T_3624 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_4040 = opcode_51 == 4'h8 | opcode_51 == 4'hb ? parameter_2_51[7:0] : _GEN_4038; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_4041 = opcode_51 == 4'h8 | opcode_51 == 4'hb ? _field_tag_T_103 : _GEN_4039; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_4042 = 14'h0 == parameter_2_51 ? phv_data_0 : _GEN_4040; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4043 = 14'h1 == parameter_2_51 ? phv_data_1 : _GEN_4042; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4044 = 14'h2 == parameter_2_51 ? phv_data_2 : _GEN_4043; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4045 = 14'h3 == parameter_2_51 ? phv_data_3 : _GEN_4044; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4046 = 14'h4 == parameter_2_51 ? phv_data_4 : _GEN_4045; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4047 = 14'h5 == parameter_2_51 ? phv_data_5 : _GEN_4046; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4048 = 14'h6 == parameter_2_51 ? phv_data_6 : _GEN_4047; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4049 = 14'h7 == parameter_2_51 ? phv_data_7 : _GEN_4048; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4050 = 14'h8 == parameter_2_51 ? phv_data_8 : _GEN_4049; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4051 = 14'h9 == parameter_2_51 ? phv_data_9 : _GEN_4050; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4052 = 14'ha == parameter_2_51 ? phv_data_10 : _GEN_4051; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4053 = 14'hb == parameter_2_51 ? phv_data_11 : _GEN_4052; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4054 = 14'hc == parameter_2_51 ? phv_data_12 : _GEN_4053; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4055 = 14'hd == parameter_2_51 ? phv_data_13 : _GEN_4054; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4056 = 14'he == parameter_2_51 ? phv_data_14 : _GEN_4055; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4057 = 14'hf == parameter_2_51 ? phv_data_15 : _GEN_4056; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4058 = 14'h10 == parameter_2_51 ? phv_data_16 : _GEN_4057; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4059 = 14'h11 == parameter_2_51 ? phv_data_17 : _GEN_4058; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4060 = 14'h12 == parameter_2_51 ? phv_data_18 : _GEN_4059; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4061 = 14'h13 == parameter_2_51 ? phv_data_19 : _GEN_4060; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4062 = 14'h14 == parameter_2_51 ? phv_data_20 : _GEN_4061; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4063 = 14'h15 == parameter_2_51 ? phv_data_21 : _GEN_4062; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4064 = 14'h16 == parameter_2_51 ? phv_data_22 : _GEN_4063; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4065 = 14'h17 == parameter_2_51 ? phv_data_23 : _GEN_4064; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4066 = 14'h18 == parameter_2_51 ? phv_data_24 : _GEN_4065; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4067 = 14'h19 == parameter_2_51 ? phv_data_25 : _GEN_4066; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4068 = 14'h1a == parameter_2_51 ? phv_data_26 : _GEN_4067; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4069 = 14'h1b == parameter_2_51 ? phv_data_27 : _GEN_4068; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4070 = 14'h1c == parameter_2_51 ? phv_data_28 : _GEN_4069; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4071 = 14'h1d == parameter_2_51 ? phv_data_29 : _GEN_4070; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4072 = 14'h1e == parameter_2_51 ? phv_data_30 : _GEN_4071; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4073 = 14'h1f == parameter_2_51 ? phv_data_31 : _GEN_4072; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4074 = 14'h20 == parameter_2_51 ? phv_data_32 : _GEN_4073; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4075 = 14'h21 == parameter_2_51 ? phv_data_33 : _GEN_4074; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4076 = 14'h22 == parameter_2_51 ? phv_data_34 : _GEN_4075; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4077 = 14'h23 == parameter_2_51 ? phv_data_35 : _GEN_4076; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4078 = 14'h24 == parameter_2_51 ? phv_data_36 : _GEN_4077; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4079 = 14'h25 == parameter_2_51 ? phv_data_37 : _GEN_4078; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4080 = 14'h26 == parameter_2_51 ? phv_data_38 : _GEN_4079; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4081 = 14'h27 == parameter_2_51 ? phv_data_39 : _GEN_4080; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4082 = 14'h28 == parameter_2_51 ? phv_data_40 : _GEN_4081; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4083 = 14'h29 == parameter_2_51 ? phv_data_41 : _GEN_4082; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4084 = 14'h2a == parameter_2_51 ? phv_data_42 : _GEN_4083; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4085 = 14'h2b == parameter_2_51 ? phv_data_43 : _GEN_4084; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4086 = 14'h2c == parameter_2_51 ? phv_data_44 : _GEN_4085; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4087 = 14'h2d == parameter_2_51 ? phv_data_45 : _GEN_4086; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4088 = 14'h2e == parameter_2_51 ? phv_data_46 : _GEN_4087; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4089 = 14'h2f == parameter_2_51 ? phv_data_47 : _GEN_4088; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4090 = 14'h30 == parameter_2_51 ? phv_data_48 : _GEN_4089; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4091 = 14'h31 == parameter_2_51 ? phv_data_49 : _GEN_4090; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4092 = 14'h32 == parameter_2_51 ? phv_data_50 : _GEN_4091; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4093 = 14'h33 == parameter_2_51 ? phv_data_51 : _GEN_4092; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4094 = 14'h34 == parameter_2_51 ? phv_data_52 : _GEN_4093; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4095 = 14'h35 == parameter_2_51 ? phv_data_53 : _GEN_4094; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4096 = 14'h36 == parameter_2_51 ? phv_data_54 : _GEN_4095; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4097 = 14'h37 == parameter_2_51 ? phv_data_55 : _GEN_4096; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4098 = 14'h38 == parameter_2_51 ? phv_data_56 : _GEN_4097; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4099 = 14'h39 == parameter_2_51 ? phv_data_57 : _GEN_4098; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4100 = 14'h3a == parameter_2_51 ? phv_data_58 : _GEN_4099; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4101 = 14'h3b == parameter_2_51 ? phv_data_59 : _GEN_4100; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4102 = 14'h3c == parameter_2_51 ? phv_data_60 : _GEN_4101; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4103 = 14'h3d == parameter_2_51 ? phv_data_61 : _GEN_4102; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4104 = 14'h3e == parameter_2_51 ? phv_data_62 : _GEN_4103; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4105 = 14'h3f == parameter_2_51 ? phv_data_63 : _GEN_4104; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_52 = vliw_52[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_52 = vliw_52[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_52 = parameter_2_52[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_52 = parameter_2_52[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_52 = {{1'd0}, args_offset_52}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_52 = _total_offset_T_52[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_4109 = 3'h1 == total_offset_52 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4110 = 3'h2 == total_offset_52 ? args_2 : _GEN_4109; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4111 = 3'h3 == total_offset_52 ? args_3 : _GEN_4110; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4112 = 3'h4 == total_offset_52 ? args_4 : _GEN_4111; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4113 = 3'h5 == total_offset_52 ? args_5 : _GEN_4112; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4114 = 3'h6 == total_offset_52 ? args_6 : _GEN_4113; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4115 = total_offset_52 < 3'h7 ? _GEN_4114 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_52_0 = 3'h0 < args_length_52 ? _GEN_4115 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_4117 = opcode_52 == 4'ha ? field_bytes_52_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_4118 = opcode_52 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_3695 = opcode_52 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_105 = _T_3695 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_4119 = opcode_52 == 4'h8 | opcode_52 == 4'hb ? parameter_2_52[7:0] : _GEN_4117; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_4120 = opcode_52 == 4'h8 | opcode_52 == 4'hb ? _field_tag_T_105 : _GEN_4118; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_4121 = 14'h0 == parameter_2_52 ? phv_data_0 : _GEN_4119; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4122 = 14'h1 == parameter_2_52 ? phv_data_1 : _GEN_4121; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4123 = 14'h2 == parameter_2_52 ? phv_data_2 : _GEN_4122; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4124 = 14'h3 == parameter_2_52 ? phv_data_3 : _GEN_4123; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4125 = 14'h4 == parameter_2_52 ? phv_data_4 : _GEN_4124; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4126 = 14'h5 == parameter_2_52 ? phv_data_5 : _GEN_4125; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4127 = 14'h6 == parameter_2_52 ? phv_data_6 : _GEN_4126; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4128 = 14'h7 == parameter_2_52 ? phv_data_7 : _GEN_4127; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4129 = 14'h8 == parameter_2_52 ? phv_data_8 : _GEN_4128; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4130 = 14'h9 == parameter_2_52 ? phv_data_9 : _GEN_4129; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4131 = 14'ha == parameter_2_52 ? phv_data_10 : _GEN_4130; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4132 = 14'hb == parameter_2_52 ? phv_data_11 : _GEN_4131; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4133 = 14'hc == parameter_2_52 ? phv_data_12 : _GEN_4132; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4134 = 14'hd == parameter_2_52 ? phv_data_13 : _GEN_4133; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4135 = 14'he == parameter_2_52 ? phv_data_14 : _GEN_4134; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4136 = 14'hf == parameter_2_52 ? phv_data_15 : _GEN_4135; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4137 = 14'h10 == parameter_2_52 ? phv_data_16 : _GEN_4136; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4138 = 14'h11 == parameter_2_52 ? phv_data_17 : _GEN_4137; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4139 = 14'h12 == parameter_2_52 ? phv_data_18 : _GEN_4138; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4140 = 14'h13 == parameter_2_52 ? phv_data_19 : _GEN_4139; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4141 = 14'h14 == parameter_2_52 ? phv_data_20 : _GEN_4140; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4142 = 14'h15 == parameter_2_52 ? phv_data_21 : _GEN_4141; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4143 = 14'h16 == parameter_2_52 ? phv_data_22 : _GEN_4142; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4144 = 14'h17 == parameter_2_52 ? phv_data_23 : _GEN_4143; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4145 = 14'h18 == parameter_2_52 ? phv_data_24 : _GEN_4144; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4146 = 14'h19 == parameter_2_52 ? phv_data_25 : _GEN_4145; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4147 = 14'h1a == parameter_2_52 ? phv_data_26 : _GEN_4146; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4148 = 14'h1b == parameter_2_52 ? phv_data_27 : _GEN_4147; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4149 = 14'h1c == parameter_2_52 ? phv_data_28 : _GEN_4148; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4150 = 14'h1d == parameter_2_52 ? phv_data_29 : _GEN_4149; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4151 = 14'h1e == parameter_2_52 ? phv_data_30 : _GEN_4150; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4152 = 14'h1f == parameter_2_52 ? phv_data_31 : _GEN_4151; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4153 = 14'h20 == parameter_2_52 ? phv_data_32 : _GEN_4152; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4154 = 14'h21 == parameter_2_52 ? phv_data_33 : _GEN_4153; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4155 = 14'h22 == parameter_2_52 ? phv_data_34 : _GEN_4154; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4156 = 14'h23 == parameter_2_52 ? phv_data_35 : _GEN_4155; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4157 = 14'h24 == parameter_2_52 ? phv_data_36 : _GEN_4156; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4158 = 14'h25 == parameter_2_52 ? phv_data_37 : _GEN_4157; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4159 = 14'h26 == parameter_2_52 ? phv_data_38 : _GEN_4158; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4160 = 14'h27 == parameter_2_52 ? phv_data_39 : _GEN_4159; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4161 = 14'h28 == parameter_2_52 ? phv_data_40 : _GEN_4160; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4162 = 14'h29 == parameter_2_52 ? phv_data_41 : _GEN_4161; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4163 = 14'h2a == parameter_2_52 ? phv_data_42 : _GEN_4162; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4164 = 14'h2b == parameter_2_52 ? phv_data_43 : _GEN_4163; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4165 = 14'h2c == parameter_2_52 ? phv_data_44 : _GEN_4164; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4166 = 14'h2d == parameter_2_52 ? phv_data_45 : _GEN_4165; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4167 = 14'h2e == parameter_2_52 ? phv_data_46 : _GEN_4166; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4168 = 14'h2f == parameter_2_52 ? phv_data_47 : _GEN_4167; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4169 = 14'h30 == parameter_2_52 ? phv_data_48 : _GEN_4168; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4170 = 14'h31 == parameter_2_52 ? phv_data_49 : _GEN_4169; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4171 = 14'h32 == parameter_2_52 ? phv_data_50 : _GEN_4170; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4172 = 14'h33 == parameter_2_52 ? phv_data_51 : _GEN_4171; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4173 = 14'h34 == parameter_2_52 ? phv_data_52 : _GEN_4172; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4174 = 14'h35 == parameter_2_52 ? phv_data_53 : _GEN_4173; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4175 = 14'h36 == parameter_2_52 ? phv_data_54 : _GEN_4174; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4176 = 14'h37 == parameter_2_52 ? phv_data_55 : _GEN_4175; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4177 = 14'h38 == parameter_2_52 ? phv_data_56 : _GEN_4176; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4178 = 14'h39 == parameter_2_52 ? phv_data_57 : _GEN_4177; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4179 = 14'h3a == parameter_2_52 ? phv_data_58 : _GEN_4178; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4180 = 14'h3b == parameter_2_52 ? phv_data_59 : _GEN_4179; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4181 = 14'h3c == parameter_2_52 ? phv_data_60 : _GEN_4180; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4182 = 14'h3d == parameter_2_52 ? phv_data_61 : _GEN_4181; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4183 = 14'h3e == parameter_2_52 ? phv_data_62 : _GEN_4182; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4184 = 14'h3f == parameter_2_52 ? phv_data_63 : _GEN_4183; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_53 = vliw_53[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_53 = vliw_53[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_53 = parameter_2_53[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_53 = parameter_2_53[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_53 = {{1'd0}, args_offset_53}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_53 = _total_offset_T_53[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_4188 = 3'h1 == total_offset_53 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4189 = 3'h2 == total_offset_53 ? args_2 : _GEN_4188; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4190 = 3'h3 == total_offset_53 ? args_3 : _GEN_4189; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4191 = 3'h4 == total_offset_53 ? args_4 : _GEN_4190; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4192 = 3'h5 == total_offset_53 ? args_5 : _GEN_4191; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4193 = 3'h6 == total_offset_53 ? args_6 : _GEN_4192; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4194 = total_offset_53 < 3'h7 ? _GEN_4193 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_53_0 = 3'h0 < args_length_53 ? _GEN_4194 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_4196 = opcode_53 == 4'ha ? field_bytes_53_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_4197 = opcode_53 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_3766 = opcode_53 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_107 = _T_3766 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_4198 = opcode_53 == 4'h8 | opcode_53 == 4'hb ? parameter_2_53[7:0] : _GEN_4196; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_4199 = opcode_53 == 4'h8 | opcode_53 == 4'hb ? _field_tag_T_107 : _GEN_4197; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_4200 = 14'h0 == parameter_2_53 ? phv_data_0 : _GEN_4198; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4201 = 14'h1 == parameter_2_53 ? phv_data_1 : _GEN_4200; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4202 = 14'h2 == parameter_2_53 ? phv_data_2 : _GEN_4201; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4203 = 14'h3 == parameter_2_53 ? phv_data_3 : _GEN_4202; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4204 = 14'h4 == parameter_2_53 ? phv_data_4 : _GEN_4203; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4205 = 14'h5 == parameter_2_53 ? phv_data_5 : _GEN_4204; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4206 = 14'h6 == parameter_2_53 ? phv_data_6 : _GEN_4205; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4207 = 14'h7 == parameter_2_53 ? phv_data_7 : _GEN_4206; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4208 = 14'h8 == parameter_2_53 ? phv_data_8 : _GEN_4207; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4209 = 14'h9 == parameter_2_53 ? phv_data_9 : _GEN_4208; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4210 = 14'ha == parameter_2_53 ? phv_data_10 : _GEN_4209; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4211 = 14'hb == parameter_2_53 ? phv_data_11 : _GEN_4210; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4212 = 14'hc == parameter_2_53 ? phv_data_12 : _GEN_4211; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4213 = 14'hd == parameter_2_53 ? phv_data_13 : _GEN_4212; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4214 = 14'he == parameter_2_53 ? phv_data_14 : _GEN_4213; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4215 = 14'hf == parameter_2_53 ? phv_data_15 : _GEN_4214; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4216 = 14'h10 == parameter_2_53 ? phv_data_16 : _GEN_4215; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4217 = 14'h11 == parameter_2_53 ? phv_data_17 : _GEN_4216; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4218 = 14'h12 == parameter_2_53 ? phv_data_18 : _GEN_4217; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4219 = 14'h13 == parameter_2_53 ? phv_data_19 : _GEN_4218; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4220 = 14'h14 == parameter_2_53 ? phv_data_20 : _GEN_4219; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4221 = 14'h15 == parameter_2_53 ? phv_data_21 : _GEN_4220; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4222 = 14'h16 == parameter_2_53 ? phv_data_22 : _GEN_4221; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4223 = 14'h17 == parameter_2_53 ? phv_data_23 : _GEN_4222; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4224 = 14'h18 == parameter_2_53 ? phv_data_24 : _GEN_4223; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4225 = 14'h19 == parameter_2_53 ? phv_data_25 : _GEN_4224; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4226 = 14'h1a == parameter_2_53 ? phv_data_26 : _GEN_4225; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4227 = 14'h1b == parameter_2_53 ? phv_data_27 : _GEN_4226; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4228 = 14'h1c == parameter_2_53 ? phv_data_28 : _GEN_4227; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4229 = 14'h1d == parameter_2_53 ? phv_data_29 : _GEN_4228; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4230 = 14'h1e == parameter_2_53 ? phv_data_30 : _GEN_4229; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4231 = 14'h1f == parameter_2_53 ? phv_data_31 : _GEN_4230; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4232 = 14'h20 == parameter_2_53 ? phv_data_32 : _GEN_4231; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4233 = 14'h21 == parameter_2_53 ? phv_data_33 : _GEN_4232; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4234 = 14'h22 == parameter_2_53 ? phv_data_34 : _GEN_4233; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4235 = 14'h23 == parameter_2_53 ? phv_data_35 : _GEN_4234; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4236 = 14'h24 == parameter_2_53 ? phv_data_36 : _GEN_4235; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4237 = 14'h25 == parameter_2_53 ? phv_data_37 : _GEN_4236; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4238 = 14'h26 == parameter_2_53 ? phv_data_38 : _GEN_4237; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4239 = 14'h27 == parameter_2_53 ? phv_data_39 : _GEN_4238; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4240 = 14'h28 == parameter_2_53 ? phv_data_40 : _GEN_4239; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4241 = 14'h29 == parameter_2_53 ? phv_data_41 : _GEN_4240; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4242 = 14'h2a == parameter_2_53 ? phv_data_42 : _GEN_4241; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4243 = 14'h2b == parameter_2_53 ? phv_data_43 : _GEN_4242; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4244 = 14'h2c == parameter_2_53 ? phv_data_44 : _GEN_4243; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4245 = 14'h2d == parameter_2_53 ? phv_data_45 : _GEN_4244; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4246 = 14'h2e == parameter_2_53 ? phv_data_46 : _GEN_4245; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4247 = 14'h2f == parameter_2_53 ? phv_data_47 : _GEN_4246; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4248 = 14'h30 == parameter_2_53 ? phv_data_48 : _GEN_4247; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4249 = 14'h31 == parameter_2_53 ? phv_data_49 : _GEN_4248; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4250 = 14'h32 == parameter_2_53 ? phv_data_50 : _GEN_4249; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4251 = 14'h33 == parameter_2_53 ? phv_data_51 : _GEN_4250; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4252 = 14'h34 == parameter_2_53 ? phv_data_52 : _GEN_4251; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4253 = 14'h35 == parameter_2_53 ? phv_data_53 : _GEN_4252; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4254 = 14'h36 == parameter_2_53 ? phv_data_54 : _GEN_4253; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4255 = 14'h37 == parameter_2_53 ? phv_data_55 : _GEN_4254; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4256 = 14'h38 == parameter_2_53 ? phv_data_56 : _GEN_4255; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4257 = 14'h39 == parameter_2_53 ? phv_data_57 : _GEN_4256; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4258 = 14'h3a == parameter_2_53 ? phv_data_58 : _GEN_4257; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4259 = 14'h3b == parameter_2_53 ? phv_data_59 : _GEN_4258; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4260 = 14'h3c == parameter_2_53 ? phv_data_60 : _GEN_4259; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4261 = 14'h3d == parameter_2_53 ? phv_data_61 : _GEN_4260; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4262 = 14'h3e == parameter_2_53 ? phv_data_62 : _GEN_4261; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4263 = 14'h3f == parameter_2_53 ? phv_data_63 : _GEN_4262; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_54 = vliw_54[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_54 = vliw_54[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_54 = parameter_2_54[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_54 = parameter_2_54[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_54 = {{1'd0}, args_offset_54}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_54 = _total_offset_T_54[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_4267 = 3'h1 == total_offset_54 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4268 = 3'h2 == total_offset_54 ? args_2 : _GEN_4267; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4269 = 3'h3 == total_offset_54 ? args_3 : _GEN_4268; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4270 = 3'h4 == total_offset_54 ? args_4 : _GEN_4269; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4271 = 3'h5 == total_offset_54 ? args_5 : _GEN_4270; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4272 = 3'h6 == total_offset_54 ? args_6 : _GEN_4271; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4273 = total_offset_54 < 3'h7 ? _GEN_4272 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_54_0 = 3'h0 < args_length_54 ? _GEN_4273 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_4275 = opcode_54 == 4'ha ? field_bytes_54_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_4276 = opcode_54 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_3837 = opcode_54 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_109 = _T_3837 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_4277 = opcode_54 == 4'h8 | opcode_54 == 4'hb ? parameter_2_54[7:0] : _GEN_4275; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_4278 = opcode_54 == 4'h8 | opcode_54 == 4'hb ? _field_tag_T_109 : _GEN_4276; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_4279 = 14'h0 == parameter_2_54 ? phv_data_0 : _GEN_4277; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4280 = 14'h1 == parameter_2_54 ? phv_data_1 : _GEN_4279; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4281 = 14'h2 == parameter_2_54 ? phv_data_2 : _GEN_4280; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4282 = 14'h3 == parameter_2_54 ? phv_data_3 : _GEN_4281; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4283 = 14'h4 == parameter_2_54 ? phv_data_4 : _GEN_4282; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4284 = 14'h5 == parameter_2_54 ? phv_data_5 : _GEN_4283; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4285 = 14'h6 == parameter_2_54 ? phv_data_6 : _GEN_4284; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4286 = 14'h7 == parameter_2_54 ? phv_data_7 : _GEN_4285; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4287 = 14'h8 == parameter_2_54 ? phv_data_8 : _GEN_4286; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4288 = 14'h9 == parameter_2_54 ? phv_data_9 : _GEN_4287; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4289 = 14'ha == parameter_2_54 ? phv_data_10 : _GEN_4288; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4290 = 14'hb == parameter_2_54 ? phv_data_11 : _GEN_4289; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4291 = 14'hc == parameter_2_54 ? phv_data_12 : _GEN_4290; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4292 = 14'hd == parameter_2_54 ? phv_data_13 : _GEN_4291; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4293 = 14'he == parameter_2_54 ? phv_data_14 : _GEN_4292; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4294 = 14'hf == parameter_2_54 ? phv_data_15 : _GEN_4293; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4295 = 14'h10 == parameter_2_54 ? phv_data_16 : _GEN_4294; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4296 = 14'h11 == parameter_2_54 ? phv_data_17 : _GEN_4295; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4297 = 14'h12 == parameter_2_54 ? phv_data_18 : _GEN_4296; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4298 = 14'h13 == parameter_2_54 ? phv_data_19 : _GEN_4297; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4299 = 14'h14 == parameter_2_54 ? phv_data_20 : _GEN_4298; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4300 = 14'h15 == parameter_2_54 ? phv_data_21 : _GEN_4299; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4301 = 14'h16 == parameter_2_54 ? phv_data_22 : _GEN_4300; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4302 = 14'h17 == parameter_2_54 ? phv_data_23 : _GEN_4301; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4303 = 14'h18 == parameter_2_54 ? phv_data_24 : _GEN_4302; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4304 = 14'h19 == parameter_2_54 ? phv_data_25 : _GEN_4303; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4305 = 14'h1a == parameter_2_54 ? phv_data_26 : _GEN_4304; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4306 = 14'h1b == parameter_2_54 ? phv_data_27 : _GEN_4305; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4307 = 14'h1c == parameter_2_54 ? phv_data_28 : _GEN_4306; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4308 = 14'h1d == parameter_2_54 ? phv_data_29 : _GEN_4307; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4309 = 14'h1e == parameter_2_54 ? phv_data_30 : _GEN_4308; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4310 = 14'h1f == parameter_2_54 ? phv_data_31 : _GEN_4309; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4311 = 14'h20 == parameter_2_54 ? phv_data_32 : _GEN_4310; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4312 = 14'h21 == parameter_2_54 ? phv_data_33 : _GEN_4311; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4313 = 14'h22 == parameter_2_54 ? phv_data_34 : _GEN_4312; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4314 = 14'h23 == parameter_2_54 ? phv_data_35 : _GEN_4313; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4315 = 14'h24 == parameter_2_54 ? phv_data_36 : _GEN_4314; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4316 = 14'h25 == parameter_2_54 ? phv_data_37 : _GEN_4315; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4317 = 14'h26 == parameter_2_54 ? phv_data_38 : _GEN_4316; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4318 = 14'h27 == parameter_2_54 ? phv_data_39 : _GEN_4317; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4319 = 14'h28 == parameter_2_54 ? phv_data_40 : _GEN_4318; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4320 = 14'h29 == parameter_2_54 ? phv_data_41 : _GEN_4319; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4321 = 14'h2a == parameter_2_54 ? phv_data_42 : _GEN_4320; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4322 = 14'h2b == parameter_2_54 ? phv_data_43 : _GEN_4321; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4323 = 14'h2c == parameter_2_54 ? phv_data_44 : _GEN_4322; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4324 = 14'h2d == parameter_2_54 ? phv_data_45 : _GEN_4323; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4325 = 14'h2e == parameter_2_54 ? phv_data_46 : _GEN_4324; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4326 = 14'h2f == parameter_2_54 ? phv_data_47 : _GEN_4325; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4327 = 14'h30 == parameter_2_54 ? phv_data_48 : _GEN_4326; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4328 = 14'h31 == parameter_2_54 ? phv_data_49 : _GEN_4327; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4329 = 14'h32 == parameter_2_54 ? phv_data_50 : _GEN_4328; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4330 = 14'h33 == parameter_2_54 ? phv_data_51 : _GEN_4329; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4331 = 14'h34 == parameter_2_54 ? phv_data_52 : _GEN_4330; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4332 = 14'h35 == parameter_2_54 ? phv_data_53 : _GEN_4331; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4333 = 14'h36 == parameter_2_54 ? phv_data_54 : _GEN_4332; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4334 = 14'h37 == parameter_2_54 ? phv_data_55 : _GEN_4333; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4335 = 14'h38 == parameter_2_54 ? phv_data_56 : _GEN_4334; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4336 = 14'h39 == parameter_2_54 ? phv_data_57 : _GEN_4335; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4337 = 14'h3a == parameter_2_54 ? phv_data_58 : _GEN_4336; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4338 = 14'h3b == parameter_2_54 ? phv_data_59 : _GEN_4337; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4339 = 14'h3c == parameter_2_54 ? phv_data_60 : _GEN_4338; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4340 = 14'h3d == parameter_2_54 ? phv_data_61 : _GEN_4339; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4341 = 14'h3e == parameter_2_54 ? phv_data_62 : _GEN_4340; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4342 = 14'h3f == parameter_2_54 ? phv_data_63 : _GEN_4341; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_55 = vliw_55[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_55 = vliw_55[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_55 = parameter_2_55[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_55 = parameter_2_55[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_55 = {{1'd0}, args_offset_55}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_55 = _total_offset_T_55[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_4346 = 3'h1 == total_offset_55 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4347 = 3'h2 == total_offset_55 ? args_2 : _GEN_4346; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4348 = 3'h3 == total_offset_55 ? args_3 : _GEN_4347; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4349 = 3'h4 == total_offset_55 ? args_4 : _GEN_4348; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4350 = 3'h5 == total_offset_55 ? args_5 : _GEN_4349; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4351 = 3'h6 == total_offset_55 ? args_6 : _GEN_4350; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4352 = total_offset_55 < 3'h7 ? _GEN_4351 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_55_0 = 3'h0 < args_length_55 ? _GEN_4352 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_4354 = opcode_55 == 4'ha ? field_bytes_55_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_4355 = opcode_55 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_3908 = opcode_55 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_111 = _T_3908 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_4356 = opcode_55 == 4'h8 | opcode_55 == 4'hb ? parameter_2_55[7:0] : _GEN_4354; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_4357 = opcode_55 == 4'h8 | opcode_55 == 4'hb ? _field_tag_T_111 : _GEN_4355; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_4358 = 14'h0 == parameter_2_55 ? phv_data_0 : _GEN_4356; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4359 = 14'h1 == parameter_2_55 ? phv_data_1 : _GEN_4358; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4360 = 14'h2 == parameter_2_55 ? phv_data_2 : _GEN_4359; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4361 = 14'h3 == parameter_2_55 ? phv_data_3 : _GEN_4360; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4362 = 14'h4 == parameter_2_55 ? phv_data_4 : _GEN_4361; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4363 = 14'h5 == parameter_2_55 ? phv_data_5 : _GEN_4362; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4364 = 14'h6 == parameter_2_55 ? phv_data_6 : _GEN_4363; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4365 = 14'h7 == parameter_2_55 ? phv_data_7 : _GEN_4364; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4366 = 14'h8 == parameter_2_55 ? phv_data_8 : _GEN_4365; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4367 = 14'h9 == parameter_2_55 ? phv_data_9 : _GEN_4366; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4368 = 14'ha == parameter_2_55 ? phv_data_10 : _GEN_4367; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4369 = 14'hb == parameter_2_55 ? phv_data_11 : _GEN_4368; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4370 = 14'hc == parameter_2_55 ? phv_data_12 : _GEN_4369; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4371 = 14'hd == parameter_2_55 ? phv_data_13 : _GEN_4370; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4372 = 14'he == parameter_2_55 ? phv_data_14 : _GEN_4371; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4373 = 14'hf == parameter_2_55 ? phv_data_15 : _GEN_4372; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4374 = 14'h10 == parameter_2_55 ? phv_data_16 : _GEN_4373; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4375 = 14'h11 == parameter_2_55 ? phv_data_17 : _GEN_4374; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4376 = 14'h12 == parameter_2_55 ? phv_data_18 : _GEN_4375; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4377 = 14'h13 == parameter_2_55 ? phv_data_19 : _GEN_4376; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4378 = 14'h14 == parameter_2_55 ? phv_data_20 : _GEN_4377; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4379 = 14'h15 == parameter_2_55 ? phv_data_21 : _GEN_4378; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4380 = 14'h16 == parameter_2_55 ? phv_data_22 : _GEN_4379; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4381 = 14'h17 == parameter_2_55 ? phv_data_23 : _GEN_4380; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4382 = 14'h18 == parameter_2_55 ? phv_data_24 : _GEN_4381; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4383 = 14'h19 == parameter_2_55 ? phv_data_25 : _GEN_4382; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4384 = 14'h1a == parameter_2_55 ? phv_data_26 : _GEN_4383; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4385 = 14'h1b == parameter_2_55 ? phv_data_27 : _GEN_4384; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4386 = 14'h1c == parameter_2_55 ? phv_data_28 : _GEN_4385; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4387 = 14'h1d == parameter_2_55 ? phv_data_29 : _GEN_4386; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4388 = 14'h1e == parameter_2_55 ? phv_data_30 : _GEN_4387; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4389 = 14'h1f == parameter_2_55 ? phv_data_31 : _GEN_4388; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4390 = 14'h20 == parameter_2_55 ? phv_data_32 : _GEN_4389; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4391 = 14'h21 == parameter_2_55 ? phv_data_33 : _GEN_4390; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4392 = 14'h22 == parameter_2_55 ? phv_data_34 : _GEN_4391; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4393 = 14'h23 == parameter_2_55 ? phv_data_35 : _GEN_4392; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4394 = 14'h24 == parameter_2_55 ? phv_data_36 : _GEN_4393; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4395 = 14'h25 == parameter_2_55 ? phv_data_37 : _GEN_4394; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4396 = 14'h26 == parameter_2_55 ? phv_data_38 : _GEN_4395; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4397 = 14'h27 == parameter_2_55 ? phv_data_39 : _GEN_4396; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4398 = 14'h28 == parameter_2_55 ? phv_data_40 : _GEN_4397; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4399 = 14'h29 == parameter_2_55 ? phv_data_41 : _GEN_4398; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4400 = 14'h2a == parameter_2_55 ? phv_data_42 : _GEN_4399; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4401 = 14'h2b == parameter_2_55 ? phv_data_43 : _GEN_4400; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4402 = 14'h2c == parameter_2_55 ? phv_data_44 : _GEN_4401; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4403 = 14'h2d == parameter_2_55 ? phv_data_45 : _GEN_4402; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4404 = 14'h2e == parameter_2_55 ? phv_data_46 : _GEN_4403; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4405 = 14'h2f == parameter_2_55 ? phv_data_47 : _GEN_4404; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4406 = 14'h30 == parameter_2_55 ? phv_data_48 : _GEN_4405; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4407 = 14'h31 == parameter_2_55 ? phv_data_49 : _GEN_4406; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4408 = 14'h32 == parameter_2_55 ? phv_data_50 : _GEN_4407; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4409 = 14'h33 == parameter_2_55 ? phv_data_51 : _GEN_4408; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4410 = 14'h34 == parameter_2_55 ? phv_data_52 : _GEN_4409; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4411 = 14'h35 == parameter_2_55 ? phv_data_53 : _GEN_4410; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4412 = 14'h36 == parameter_2_55 ? phv_data_54 : _GEN_4411; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4413 = 14'h37 == parameter_2_55 ? phv_data_55 : _GEN_4412; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4414 = 14'h38 == parameter_2_55 ? phv_data_56 : _GEN_4413; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4415 = 14'h39 == parameter_2_55 ? phv_data_57 : _GEN_4414; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4416 = 14'h3a == parameter_2_55 ? phv_data_58 : _GEN_4415; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4417 = 14'h3b == parameter_2_55 ? phv_data_59 : _GEN_4416; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4418 = 14'h3c == parameter_2_55 ? phv_data_60 : _GEN_4417; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4419 = 14'h3d == parameter_2_55 ? phv_data_61 : _GEN_4418; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4420 = 14'h3e == parameter_2_55 ? phv_data_62 : _GEN_4419; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4421 = 14'h3f == parameter_2_55 ? phv_data_63 : _GEN_4420; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_56 = vliw_56[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_56 = vliw_56[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_56 = parameter_2_56[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_56 = parameter_2_56[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_56 = {{1'd0}, args_offset_56}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_56 = _total_offset_T_56[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_4425 = 3'h1 == total_offset_56 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4426 = 3'h2 == total_offset_56 ? args_2 : _GEN_4425; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4427 = 3'h3 == total_offset_56 ? args_3 : _GEN_4426; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4428 = 3'h4 == total_offset_56 ? args_4 : _GEN_4427; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4429 = 3'h5 == total_offset_56 ? args_5 : _GEN_4428; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4430 = 3'h6 == total_offset_56 ? args_6 : _GEN_4429; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4431 = total_offset_56 < 3'h7 ? _GEN_4430 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_56_0 = 3'h0 < args_length_56 ? _GEN_4431 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_4433 = opcode_56 == 4'ha ? field_bytes_56_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_4434 = opcode_56 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_3979 = opcode_56 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_113 = _T_3979 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_4435 = opcode_56 == 4'h8 | opcode_56 == 4'hb ? parameter_2_56[7:0] : _GEN_4433; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_4436 = opcode_56 == 4'h8 | opcode_56 == 4'hb ? _field_tag_T_113 : _GEN_4434; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_4437 = 14'h0 == parameter_2_56 ? phv_data_0 : _GEN_4435; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4438 = 14'h1 == parameter_2_56 ? phv_data_1 : _GEN_4437; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4439 = 14'h2 == parameter_2_56 ? phv_data_2 : _GEN_4438; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4440 = 14'h3 == parameter_2_56 ? phv_data_3 : _GEN_4439; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4441 = 14'h4 == parameter_2_56 ? phv_data_4 : _GEN_4440; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4442 = 14'h5 == parameter_2_56 ? phv_data_5 : _GEN_4441; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4443 = 14'h6 == parameter_2_56 ? phv_data_6 : _GEN_4442; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4444 = 14'h7 == parameter_2_56 ? phv_data_7 : _GEN_4443; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4445 = 14'h8 == parameter_2_56 ? phv_data_8 : _GEN_4444; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4446 = 14'h9 == parameter_2_56 ? phv_data_9 : _GEN_4445; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4447 = 14'ha == parameter_2_56 ? phv_data_10 : _GEN_4446; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4448 = 14'hb == parameter_2_56 ? phv_data_11 : _GEN_4447; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4449 = 14'hc == parameter_2_56 ? phv_data_12 : _GEN_4448; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4450 = 14'hd == parameter_2_56 ? phv_data_13 : _GEN_4449; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4451 = 14'he == parameter_2_56 ? phv_data_14 : _GEN_4450; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4452 = 14'hf == parameter_2_56 ? phv_data_15 : _GEN_4451; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4453 = 14'h10 == parameter_2_56 ? phv_data_16 : _GEN_4452; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4454 = 14'h11 == parameter_2_56 ? phv_data_17 : _GEN_4453; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4455 = 14'h12 == parameter_2_56 ? phv_data_18 : _GEN_4454; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4456 = 14'h13 == parameter_2_56 ? phv_data_19 : _GEN_4455; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4457 = 14'h14 == parameter_2_56 ? phv_data_20 : _GEN_4456; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4458 = 14'h15 == parameter_2_56 ? phv_data_21 : _GEN_4457; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4459 = 14'h16 == parameter_2_56 ? phv_data_22 : _GEN_4458; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4460 = 14'h17 == parameter_2_56 ? phv_data_23 : _GEN_4459; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4461 = 14'h18 == parameter_2_56 ? phv_data_24 : _GEN_4460; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4462 = 14'h19 == parameter_2_56 ? phv_data_25 : _GEN_4461; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4463 = 14'h1a == parameter_2_56 ? phv_data_26 : _GEN_4462; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4464 = 14'h1b == parameter_2_56 ? phv_data_27 : _GEN_4463; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4465 = 14'h1c == parameter_2_56 ? phv_data_28 : _GEN_4464; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4466 = 14'h1d == parameter_2_56 ? phv_data_29 : _GEN_4465; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4467 = 14'h1e == parameter_2_56 ? phv_data_30 : _GEN_4466; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4468 = 14'h1f == parameter_2_56 ? phv_data_31 : _GEN_4467; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4469 = 14'h20 == parameter_2_56 ? phv_data_32 : _GEN_4468; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4470 = 14'h21 == parameter_2_56 ? phv_data_33 : _GEN_4469; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4471 = 14'h22 == parameter_2_56 ? phv_data_34 : _GEN_4470; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4472 = 14'h23 == parameter_2_56 ? phv_data_35 : _GEN_4471; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4473 = 14'h24 == parameter_2_56 ? phv_data_36 : _GEN_4472; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4474 = 14'h25 == parameter_2_56 ? phv_data_37 : _GEN_4473; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4475 = 14'h26 == parameter_2_56 ? phv_data_38 : _GEN_4474; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4476 = 14'h27 == parameter_2_56 ? phv_data_39 : _GEN_4475; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4477 = 14'h28 == parameter_2_56 ? phv_data_40 : _GEN_4476; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4478 = 14'h29 == parameter_2_56 ? phv_data_41 : _GEN_4477; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4479 = 14'h2a == parameter_2_56 ? phv_data_42 : _GEN_4478; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4480 = 14'h2b == parameter_2_56 ? phv_data_43 : _GEN_4479; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4481 = 14'h2c == parameter_2_56 ? phv_data_44 : _GEN_4480; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4482 = 14'h2d == parameter_2_56 ? phv_data_45 : _GEN_4481; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4483 = 14'h2e == parameter_2_56 ? phv_data_46 : _GEN_4482; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4484 = 14'h2f == parameter_2_56 ? phv_data_47 : _GEN_4483; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4485 = 14'h30 == parameter_2_56 ? phv_data_48 : _GEN_4484; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4486 = 14'h31 == parameter_2_56 ? phv_data_49 : _GEN_4485; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4487 = 14'h32 == parameter_2_56 ? phv_data_50 : _GEN_4486; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4488 = 14'h33 == parameter_2_56 ? phv_data_51 : _GEN_4487; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4489 = 14'h34 == parameter_2_56 ? phv_data_52 : _GEN_4488; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4490 = 14'h35 == parameter_2_56 ? phv_data_53 : _GEN_4489; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4491 = 14'h36 == parameter_2_56 ? phv_data_54 : _GEN_4490; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4492 = 14'h37 == parameter_2_56 ? phv_data_55 : _GEN_4491; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4493 = 14'h38 == parameter_2_56 ? phv_data_56 : _GEN_4492; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4494 = 14'h39 == parameter_2_56 ? phv_data_57 : _GEN_4493; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4495 = 14'h3a == parameter_2_56 ? phv_data_58 : _GEN_4494; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4496 = 14'h3b == parameter_2_56 ? phv_data_59 : _GEN_4495; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4497 = 14'h3c == parameter_2_56 ? phv_data_60 : _GEN_4496; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4498 = 14'h3d == parameter_2_56 ? phv_data_61 : _GEN_4497; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4499 = 14'h3e == parameter_2_56 ? phv_data_62 : _GEN_4498; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4500 = 14'h3f == parameter_2_56 ? phv_data_63 : _GEN_4499; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_57 = vliw_57[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_57 = vliw_57[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_57 = parameter_2_57[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_57 = parameter_2_57[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_57 = {{1'd0}, args_offset_57}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_57 = _total_offset_T_57[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_4504 = 3'h1 == total_offset_57 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4505 = 3'h2 == total_offset_57 ? args_2 : _GEN_4504; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4506 = 3'h3 == total_offset_57 ? args_3 : _GEN_4505; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4507 = 3'h4 == total_offset_57 ? args_4 : _GEN_4506; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4508 = 3'h5 == total_offset_57 ? args_5 : _GEN_4507; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4509 = 3'h6 == total_offset_57 ? args_6 : _GEN_4508; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4510 = total_offset_57 < 3'h7 ? _GEN_4509 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_57_0 = 3'h0 < args_length_57 ? _GEN_4510 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_4512 = opcode_57 == 4'ha ? field_bytes_57_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_4513 = opcode_57 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_4050 = opcode_57 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_115 = _T_4050 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_4514 = opcode_57 == 4'h8 | opcode_57 == 4'hb ? parameter_2_57[7:0] : _GEN_4512; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_4515 = opcode_57 == 4'h8 | opcode_57 == 4'hb ? _field_tag_T_115 : _GEN_4513; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_4516 = 14'h0 == parameter_2_57 ? phv_data_0 : _GEN_4514; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4517 = 14'h1 == parameter_2_57 ? phv_data_1 : _GEN_4516; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4518 = 14'h2 == parameter_2_57 ? phv_data_2 : _GEN_4517; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4519 = 14'h3 == parameter_2_57 ? phv_data_3 : _GEN_4518; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4520 = 14'h4 == parameter_2_57 ? phv_data_4 : _GEN_4519; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4521 = 14'h5 == parameter_2_57 ? phv_data_5 : _GEN_4520; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4522 = 14'h6 == parameter_2_57 ? phv_data_6 : _GEN_4521; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4523 = 14'h7 == parameter_2_57 ? phv_data_7 : _GEN_4522; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4524 = 14'h8 == parameter_2_57 ? phv_data_8 : _GEN_4523; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4525 = 14'h9 == parameter_2_57 ? phv_data_9 : _GEN_4524; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4526 = 14'ha == parameter_2_57 ? phv_data_10 : _GEN_4525; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4527 = 14'hb == parameter_2_57 ? phv_data_11 : _GEN_4526; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4528 = 14'hc == parameter_2_57 ? phv_data_12 : _GEN_4527; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4529 = 14'hd == parameter_2_57 ? phv_data_13 : _GEN_4528; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4530 = 14'he == parameter_2_57 ? phv_data_14 : _GEN_4529; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4531 = 14'hf == parameter_2_57 ? phv_data_15 : _GEN_4530; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4532 = 14'h10 == parameter_2_57 ? phv_data_16 : _GEN_4531; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4533 = 14'h11 == parameter_2_57 ? phv_data_17 : _GEN_4532; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4534 = 14'h12 == parameter_2_57 ? phv_data_18 : _GEN_4533; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4535 = 14'h13 == parameter_2_57 ? phv_data_19 : _GEN_4534; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4536 = 14'h14 == parameter_2_57 ? phv_data_20 : _GEN_4535; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4537 = 14'h15 == parameter_2_57 ? phv_data_21 : _GEN_4536; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4538 = 14'h16 == parameter_2_57 ? phv_data_22 : _GEN_4537; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4539 = 14'h17 == parameter_2_57 ? phv_data_23 : _GEN_4538; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4540 = 14'h18 == parameter_2_57 ? phv_data_24 : _GEN_4539; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4541 = 14'h19 == parameter_2_57 ? phv_data_25 : _GEN_4540; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4542 = 14'h1a == parameter_2_57 ? phv_data_26 : _GEN_4541; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4543 = 14'h1b == parameter_2_57 ? phv_data_27 : _GEN_4542; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4544 = 14'h1c == parameter_2_57 ? phv_data_28 : _GEN_4543; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4545 = 14'h1d == parameter_2_57 ? phv_data_29 : _GEN_4544; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4546 = 14'h1e == parameter_2_57 ? phv_data_30 : _GEN_4545; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4547 = 14'h1f == parameter_2_57 ? phv_data_31 : _GEN_4546; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4548 = 14'h20 == parameter_2_57 ? phv_data_32 : _GEN_4547; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4549 = 14'h21 == parameter_2_57 ? phv_data_33 : _GEN_4548; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4550 = 14'h22 == parameter_2_57 ? phv_data_34 : _GEN_4549; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4551 = 14'h23 == parameter_2_57 ? phv_data_35 : _GEN_4550; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4552 = 14'h24 == parameter_2_57 ? phv_data_36 : _GEN_4551; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4553 = 14'h25 == parameter_2_57 ? phv_data_37 : _GEN_4552; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4554 = 14'h26 == parameter_2_57 ? phv_data_38 : _GEN_4553; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4555 = 14'h27 == parameter_2_57 ? phv_data_39 : _GEN_4554; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4556 = 14'h28 == parameter_2_57 ? phv_data_40 : _GEN_4555; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4557 = 14'h29 == parameter_2_57 ? phv_data_41 : _GEN_4556; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4558 = 14'h2a == parameter_2_57 ? phv_data_42 : _GEN_4557; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4559 = 14'h2b == parameter_2_57 ? phv_data_43 : _GEN_4558; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4560 = 14'h2c == parameter_2_57 ? phv_data_44 : _GEN_4559; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4561 = 14'h2d == parameter_2_57 ? phv_data_45 : _GEN_4560; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4562 = 14'h2e == parameter_2_57 ? phv_data_46 : _GEN_4561; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4563 = 14'h2f == parameter_2_57 ? phv_data_47 : _GEN_4562; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4564 = 14'h30 == parameter_2_57 ? phv_data_48 : _GEN_4563; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4565 = 14'h31 == parameter_2_57 ? phv_data_49 : _GEN_4564; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4566 = 14'h32 == parameter_2_57 ? phv_data_50 : _GEN_4565; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4567 = 14'h33 == parameter_2_57 ? phv_data_51 : _GEN_4566; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4568 = 14'h34 == parameter_2_57 ? phv_data_52 : _GEN_4567; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4569 = 14'h35 == parameter_2_57 ? phv_data_53 : _GEN_4568; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4570 = 14'h36 == parameter_2_57 ? phv_data_54 : _GEN_4569; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4571 = 14'h37 == parameter_2_57 ? phv_data_55 : _GEN_4570; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4572 = 14'h38 == parameter_2_57 ? phv_data_56 : _GEN_4571; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4573 = 14'h39 == parameter_2_57 ? phv_data_57 : _GEN_4572; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4574 = 14'h3a == parameter_2_57 ? phv_data_58 : _GEN_4573; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4575 = 14'h3b == parameter_2_57 ? phv_data_59 : _GEN_4574; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4576 = 14'h3c == parameter_2_57 ? phv_data_60 : _GEN_4575; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4577 = 14'h3d == parameter_2_57 ? phv_data_61 : _GEN_4576; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4578 = 14'h3e == parameter_2_57 ? phv_data_62 : _GEN_4577; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4579 = 14'h3f == parameter_2_57 ? phv_data_63 : _GEN_4578; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_58 = vliw_58[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_58 = vliw_58[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_58 = parameter_2_58[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_58 = parameter_2_58[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_58 = {{1'd0}, args_offset_58}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_58 = _total_offset_T_58[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_4583 = 3'h1 == total_offset_58 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4584 = 3'h2 == total_offset_58 ? args_2 : _GEN_4583; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4585 = 3'h3 == total_offset_58 ? args_3 : _GEN_4584; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4586 = 3'h4 == total_offset_58 ? args_4 : _GEN_4585; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4587 = 3'h5 == total_offset_58 ? args_5 : _GEN_4586; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4588 = 3'h6 == total_offset_58 ? args_6 : _GEN_4587; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4589 = total_offset_58 < 3'h7 ? _GEN_4588 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_58_0 = 3'h0 < args_length_58 ? _GEN_4589 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_4591 = opcode_58 == 4'ha ? field_bytes_58_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_4592 = opcode_58 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_4121 = opcode_58 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_117 = _T_4121 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_4593 = opcode_58 == 4'h8 | opcode_58 == 4'hb ? parameter_2_58[7:0] : _GEN_4591; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_4594 = opcode_58 == 4'h8 | opcode_58 == 4'hb ? _field_tag_T_117 : _GEN_4592; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_4595 = 14'h0 == parameter_2_58 ? phv_data_0 : _GEN_4593; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4596 = 14'h1 == parameter_2_58 ? phv_data_1 : _GEN_4595; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4597 = 14'h2 == parameter_2_58 ? phv_data_2 : _GEN_4596; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4598 = 14'h3 == parameter_2_58 ? phv_data_3 : _GEN_4597; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4599 = 14'h4 == parameter_2_58 ? phv_data_4 : _GEN_4598; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4600 = 14'h5 == parameter_2_58 ? phv_data_5 : _GEN_4599; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4601 = 14'h6 == parameter_2_58 ? phv_data_6 : _GEN_4600; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4602 = 14'h7 == parameter_2_58 ? phv_data_7 : _GEN_4601; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4603 = 14'h8 == parameter_2_58 ? phv_data_8 : _GEN_4602; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4604 = 14'h9 == parameter_2_58 ? phv_data_9 : _GEN_4603; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4605 = 14'ha == parameter_2_58 ? phv_data_10 : _GEN_4604; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4606 = 14'hb == parameter_2_58 ? phv_data_11 : _GEN_4605; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4607 = 14'hc == parameter_2_58 ? phv_data_12 : _GEN_4606; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4608 = 14'hd == parameter_2_58 ? phv_data_13 : _GEN_4607; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4609 = 14'he == parameter_2_58 ? phv_data_14 : _GEN_4608; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4610 = 14'hf == parameter_2_58 ? phv_data_15 : _GEN_4609; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4611 = 14'h10 == parameter_2_58 ? phv_data_16 : _GEN_4610; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4612 = 14'h11 == parameter_2_58 ? phv_data_17 : _GEN_4611; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4613 = 14'h12 == parameter_2_58 ? phv_data_18 : _GEN_4612; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4614 = 14'h13 == parameter_2_58 ? phv_data_19 : _GEN_4613; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4615 = 14'h14 == parameter_2_58 ? phv_data_20 : _GEN_4614; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4616 = 14'h15 == parameter_2_58 ? phv_data_21 : _GEN_4615; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4617 = 14'h16 == parameter_2_58 ? phv_data_22 : _GEN_4616; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4618 = 14'h17 == parameter_2_58 ? phv_data_23 : _GEN_4617; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4619 = 14'h18 == parameter_2_58 ? phv_data_24 : _GEN_4618; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4620 = 14'h19 == parameter_2_58 ? phv_data_25 : _GEN_4619; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4621 = 14'h1a == parameter_2_58 ? phv_data_26 : _GEN_4620; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4622 = 14'h1b == parameter_2_58 ? phv_data_27 : _GEN_4621; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4623 = 14'h1c == parameter_2_58 ? phv_data_28 : _GEN_4622; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4624 = 14'h1d == parameter_2_58 ? phv_data_29 : _GEN_4623; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4625 = 14'h1e == parameter_2_58 ? phv_data_30 : _GEN_4624; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4626 = 14'h1f == parameter_2_58 ? phv_data_31 : _GEN_4625; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4627 = 14'h20 == parameter_2_58 ? phv_data_32 : _GEN_4626; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4628 = 14'h21 == parameter_2_58 ? phv_data_33 : _GEN_4627; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4629 = 14'h22 == parameter_2_58 ? phv_data_34 : _GEN_4628; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4630 = 14'h23 == parameter_2_58 ? phv_data_35 : _GEN_4629; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4631 = 14'h24 == parameter_2_58 ? phv_data_36 : _GEN_4630; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4632 = 14'h25 == parameter_2_58 ? phv_data_37 : _GEN_4631; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4633 = 14'h26 == parameter_2_58 ? phv_data_38 : _GEN_4632; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4634 = 14'h27 == parameter_2_58 ? phv_data_39 : _GEN_4633; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4635 = 14'h28 == parameter_2_58 ? phv_data_40 : _GEN_4634; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4636 = 14'h29 == parameter_2_58 ? phv_data_41 : _GEN_4635; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4637 = 14'h2a == parameter_2_58 ? phv_data_42 : _GEN_4636; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4638 = 14'h2b == parameter_2_58 ? phv_data_43 : _GEN_4637; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4639 = 14'h2c == parameter_2_58 ? phv_data_44 : _GEN_4638; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4640 = 14'h2d == parameter_2_58 ? phv_data_45 : _GEN_4639; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4641 = 14'h2e == parameter_2_58 ? phv_data_46 : _GEN_4640; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4642 = 14'h2f == parameter_2_58 ? phv_data_47 : _GEN_4641; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4643 = 14'h30 == parameter_2_58 ? phv_data_48 : _GEN_4642; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4644 = 14'h31 == parameter_2_58 ? phv_data_49 : _GEN_4643; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4645 = 14'h32 == parameter_2_58 ? phv_data_50 : _GEN_4644; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4646 = 14'h33 == parameter_2_58 ? phv_data_51 : _GEN_4645; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4647 = 14'h34 == parameter_2_58 ? phv_data_52 : _GEN_4646; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4648 = 14'h35 == parameter_2_58 ? phv_data_53 : _GEN_4647; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4649 = 14'h36 == parameter_2_58 ? phv_data_54 : _GEN_4648; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4650 = 14'h37 == parameter_2_58 ? phv_data_55 : _GEN_4649; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4651 = 14'h38 == parameter_2_58 ? phv_data_56 : _GEN_4650; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4652 = 14'h39 == parameter_2_58 ? phv_data_57 : _GEN_4651; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4653 = 14'h3a == parameter_2_58 ? phv_data_58 : _GEN_4652; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4654 = 14'h3b == parameter_2_58 ? phv_data_59 : _GEN_4653; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4655 = 14'h3c == parameter_2_58 ? phv_data_60 : _GEN_4654; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4656 = 14'h3d == parameter_2_58 ? phv_data_61 : _GEN_4655; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4657 = 14'h3e == parameter_2_58 ? phv_data_62 : _GEN_4656; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4658 = 14'h3f == parameter_2_58 ? phv_data_63 : _GEN_4657; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_59 = vliw_59[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_59 = vliw_59[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_59 = parameter_2_59[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_59 = parameter_2_59[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_59 = {{1'd0}, args_offset_59}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_59 = _total_offset_T_59[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_4662 = 3'h1 == total_offset_59 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4663 = 3'h2 == total_offset_59 ? args_2 : _GEN_4662; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4664 = 3'h3 == total_offset_59 ? args_3 : _GEN_4663; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4665 = 3'h4 == total_offset_59 ? args_4 : _GEN_4664; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4666 = 3'h5 == total_offset_59 ? args_5 : _GEN_4665; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4667 = 3'h6 == total_offset_59 ? args_6 : _GEN_4666; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4668 = total_offset_59 < 3'h7 ? _GEN_4667 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_59_0 = 3'h0 < args_length_59 ? _GEN_4668 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_4670 = opcode_59 == 4'ha ? field_bytes_59_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_4671 = opcode_59 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_4192 = opcode_59 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_119 = _T_4192 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_4672 = opcode_59 == 4'h8 | opcode_59 == 4'hb ? parameter_2_59[7:0] : _GEN_4670; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_4673 = opcode_59 == 4'h8 | opcode_59 == 4'hb ? _field_tag_T_119 : _GEN_4671; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_4674 = 14'h0 == parameter_2_59 ? phv_data_0 : _GEN_4672; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4675 = 14'h1 == parameter_2_59 ? phv_data_1 : _GEN_4674; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4676 = 14'h2 == parameter_2_59 ? phv_data_2 : _GEN_4675; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4677 = 14'h3 == parameter_2_59 ? phv_data_3 : _GEN_4676; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4678 = 14'h4 == parameter_2_59 ? phv_data_4 : _GEN_4677; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4679 = 14'h5 == parameter_2_59 ? phv_data_5 : _GEN_4678; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4680 = 14'h6 == parameter_2_59 ? phv_data_6 : _GEN_4679; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4681 = 14'h7 == parameter_2_59 ? phv_data_7 : _GEN_4680; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4682 = 14'h8 == parameter_2_59 ? phv_data_8 : _GEN_4681; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4683 = 14'h9 == parameter_2_59 ? phv_data_9 : _GEN_4682; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4684 = 14'ha == parameter_2_59 ? phv_data_10 : _GEN_4683; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4685 = 14'hb == parameter_2_59 ? phv_data_11 : _GEN_4684; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4686 = 14'hc == parameter_2_59 ? phv_data_12 : _GEN_4685; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4687 = 14'hd == parameter_2_59 ? phv_data_13 : _GEN_4686; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4688 = 14'he == parameter_2_59 ? phv_data_14 : _GEN_4687; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4689 = 14'hf == parameter_2_59 ? phv_data_15 : _GEN_4688; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4690 = 14'h10 == parameter_2_59 ? phv_data_16 : _GEN_4689; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4691 = 14'h11 == parameter_2_59 ? phv_data_17 : _GEN_4690; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4692 = 14'h12 == parameter_2_59 ? phv_data_18 : _GEN_4691; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4693 = 14'h13 == parameter_2_59 ? phv_data_19 : _GEN_4692; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4694 = 14'h14 == parameter_2_59 ? phv_data_20 : _GEN_4693; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4695 = 14'h15 == parameter_2_59 ? phv_data_21 : _GEN_4694; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4696 = 14'h16 == parameter_2_59 ? phv_data_22 : _GEN_4695; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4697 = 14'h17 == parameter_2_59 ? phv_data_23 : _GEN_4696; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4698 = 14'h18 == parameter_2_59 ? phv_data_24 : _GEN_4697; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4699 = 14'h19 == parameter_2_59 ? phv_data_25 : _GEN_4698; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4700 = 14'h1a == parameter_2_59 ? phv_data_26 : _GEN_4699; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4701 = 14'h1b == parameter_2_59 ? phv_data_27 : _GEN_4700; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4702 = 14'h1c == parameter_2_59 ? phv_data_28 : _GEN_4701; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4703 = 14'h1d == parameter_2_59 ? phv_data_29 : _GEN_4702; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4704 = 14'h1e == parameter_2_59 ? phv_data_30 : _GEN_4703; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4705 = 14'h1f == parameter_2_59 ? phv_data_31 : _GEN_4704; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4706 = 14'h20 == parameter_2_59 ? phv_data_32 : _GEN_4705; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4707 = 14'h21 == parameter_2_59 ? phv_data_33 : _GEN_4706; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4708 = 14'h22 == parameter_2_59 ? phv_data_34 : _GEN_4707; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4709 = 14'h23 == parameter_2_59 ? phv_data_35 : _GEN_4708; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4710 = 14'h24 == parameter_2_59 ? phv_data_36 : _GEN_4709; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4711 = 14'h25 == parameter_2_59 ? phv_data_37 : _GEN_4710; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4712 = 14'h26 == parameter_2_59 ? phv_data_38 : _GEN_4711; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4713 = 14'h27 == parameter_2_59 ? phv_data_39 : _GEN_4712; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4714 = 14'h28 == parameter_2_59 ? phv_data_40 : _GEN_4713; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4715 = 14'h29 == parameter_2_59 ? phv_data_41 : _GEN_4714; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4716 = 14'h2a == parameter_2_59 ? phv_data_42 : _GEN_4715; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4717 = 14'h2b == parameter_2_59 ? phv_data_43 : _GEN_4716; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4718 = 14'h2c == parameter_2_59 ? phv_data_44 : _GEN_4717; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4719 = 14'h2d == parameter_2_59 ? phv_data_45 : _GEN_4718; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4720 = 14'h2e == parameter_2_59 ? phv_data_46 : _GEN_4719; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4721 = 14'h2f == parameter_2_59 ? phv_data_47 : _GEN_4720; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4722 = 14'h30 == parameter_2_59 ? phv_data_48 : _GEN_4721; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4723 = 14'h31 == parameter_2_59 ? phv_data_49 : _GEN_4722; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4724 = 14'h32 == parameter_2_59 ? phv_data_50 : _GEN_4723; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4725 = 14'h33 == parameter_2_59 ? phv_data_51 : _GEN_4724; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4726 = 14'h34 == parameter_2_59 ? phv_data_52 : _GEN_4725; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4727 = 14'h35 == parameter_2_59 ? phv_data_53 : _GEN_4726; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4728 = 14'h36 == parameter_2_59 ? phv_data_54 : _GEN_4727; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4729 = 14'h37 == parameter_2_59 ? phv_data_55 : _GEN_4728; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4730 = 14'h38 == parameter_2_59 ? phv_data_56 : _GEN_4729; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4731 = 14'h39 == parameter_2_59 ? phv_data_57 : _GEN_4730; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4732 = 14'h3a == parameter_2_59 ? phv_data_58 : _GEN_4731; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4733 = 14'h3b == parameter_2_59 ? phv_data_59 : _GEN_4732; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4734 = 14'h3c == parameter_2_59 ? phv_data_60 : _GEN_4733; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4735 = 14'h3d == parameter_2_59 ? phv_data_61 : _GEN_4734; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4736 = 14'h3e == parameter_2_59 ? phv_data_62 : _GEN_4735; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4737 = 14'h3f == parameter_2_59 ? phv_data_63 : _GEN_4736; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_60 = vliw_60[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_60 = vliw_60[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_60 = parameter_2_60[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_60 = parameter_2_60[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_60 = {{1'd0}, args_offset_60}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_60 = _total_offset_T_60[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_4741 = 3'h1 == total_offset_60 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4742 = 3'h2 == total_offset_60 ? args_2 : _GEN_4741; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4743 = 3'h3 == total_offset_60 ? args_3 : _GEN_4742; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4744 = 3'h4 == total_offset_60 ? args_4 : _GEN_4743; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4745 = 3'h5 == total_offset_60 ? args_5 : _GEN_4744; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4746 = 3'h6 == total_offset_60 ? args_6 : _GEN_4745; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4747 = total_offset_60 < 3'h7 ? _GEN_4746 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_60_0 = 3'h0 < args_length_60 ? _GEN_4747 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_4749 = opcode_60 == 4'ha ? field_bytes_60_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_4750 = opcode_60 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_4263 = opcode_60 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_121 = _T_4263 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_4751 = opcode_60 == 4'h8 | opcode_60 == 4'hb ? parameter_2_60[7:0] : _GEN_4749; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_4752 = opcode_60 == 4'h8 | opcode_60 == 4'hb ? _field_tag_T_121 : _GEN_4750; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_4753 = 14'h0 == parameter_2_60 ? phv_data_0 : _GEN_4751; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4754 = 14'h1 == parameter_2_60 ? phv_data_1 : _GEN_4753; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4755 = 14'h2 == parameter_2_60 ? phv_data_2 : _GEN_4754; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4756 = 14'h3 == parameter_2_60 ? phv_data_3 : _GEN_4755; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4757 = 14'h4 == parameter_2_60 ? phv_data_4 : _GEN_4756; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4758 = 14'h5 == parameter_2_60 ? phv_data_5 : _GEN_4757; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4759 = 14'h6 == parameter_2_60 ? phv_data_6 : _GEN_4758; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4760 = 14'h7 == parameter_2_60 ? phv_data_7 : _GEN_4759; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4761 = 14'h8 == parameter_2_60 ? phv_data_8 : _GEN_4760; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4762 = 14'h9 == parameter_2_60 ? phv_data_9 : _GEN_4761; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4763 = 14'ha == parameter_2_60 ? phv_data_10 : _GEN_4762; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4764 = 14'hb == parameter_2_60 ? phv_data_11 : _GEN_4763; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4765 = 14'hc == parameter_2_60 ? phv_data_12 : _GEN_4764; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4766 = 14'hd == parameter_2_60 ? phv_data_13 : _GEN_4765; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4767 = 14'he == parameter_2_60 ? phv_data_14 : _GEN_4766; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4768 = 14'hf == parameter_2_60 ? phv_data_15 : _GEN_4767; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4769 = 14'h10 == parameter_2_60 ? phv_data_16 : _GEN_4768; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4770 = 14'h11 == parameter_2_60 ? phv_data_17 : _GEN_4769; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4771 = 14'h12 == parameter_2_60 ? phv_data_18 : _GEN_4770; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4772 = 14'h13 == parameter_2_60 ? phv_data_19 : _GEN_4771; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4773 = 14'h14 == parameter_2_60 ? phv_data_20 : _GEN_4772; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4774 = 14'h15 == parameter_2_60 ? phv_data_21 : _GEN_4773; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4775 = 14'h16 == parameter_2_60 ? phv_data_22 : _GEN_4774; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4776 = 14'h17 == parameter_2_60 ? phv_data_23 : _GEN_4775; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4777 = 14'h18 == parameter_2_60 ? phv_data_24 : _GEN_4776; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4778 = 14'h19 == parameter_2_60 ? phv_data_25 : _GEN_4777; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4779 = 14'h1a == parameter_2_60 ? phv_data_26 : _GEN_4778; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4780 = 14'h1b == parameter_2_60 ? phv_data_27 : _GEN_4779; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4781 = 14'h1c == parameter_2_60 ? phv_data_28 : _GEN_4780; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4782 = 14'h1d == parameter_2_60 ? phv_data_29 : _GEN_4781; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4783 = 14'h1e == parameter_2_60 ? phv_data_30 : _GEN_4782; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4784 = 14'h1f == parameter_2_60 ? phv_data_31 : _GEN_4783; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4785 = 14'h20 == parameter_2_60 ? phv_data_32 : _GEN_4784; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4786 = 14'h21 == parameter_2_60 ? phv_data_33 : _GEN_4785; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4787 = 14'h22 == parameter_2_60 ? phv_data_34 : _GEN_4786; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4788 = 14'h23 == parameter_2_60 ? phv_data_35 : _GEN_4787; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4789 = 14'h24 == parameter_2_60 ? phv_data_36 : _GEN_4788; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4790 = 14'h25 == parameter_2_60 ? phv_data_37 : _GEN_4789; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4791 = 14'h26 == parameter_2_60 ? phv_data_38 : _GEN_4790; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4792 = 14'h27 == parameter_2_60 ? phv_data_39 : _GEN_4791; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4793 = 14'h28 == parameter_2_60 ? phv_data_40 : _GEN_4792; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4794 = 14'h29 == parameter_2_60 ? phv_data_41 : _GEN_4793; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4795 = 14'h2a == parameter_2_60 ? phv_data_42 : _GEN_4794; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4796 = 14'h2b == parameter_2_60 ? phv_data_43 : _GEN_4795; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4797 = 14'h2c == parameter_2_60 ? phv_data_44 : _GEN_4796; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4798 = 14'h2d == parameter_2_60 ? phv_data_45 : _GEN_4797; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4799 = 14'h2e == parameter_2_60 ? phv_data_46 : _GEN_4798; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4800 = 14'h2f == parameter_2_60 ? phv_data_47 : _GEN_4799; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4801 = 14'h30 == parameter_2_60 ? phv_data_48 : _GEN_4800; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4802 = 14'h31 == parameter_2_60 ? phv_data_49 : _GEN_4801; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4803 = 14'h32 == parameter_2_60 ? phv_data_50 : _GEN_4802; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4804 = 14'h33 == parameter_2_60 ? phv_data_51 : _GEN_4803; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4805 = 14'h34 == parameter_2_60 ? phv_data_52 : _GEN_4804; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4806 = 14'h35 == parameter_2_60 ? phv_data_53 : _GEN_4805; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4807 = 14'h36 == parameter_2_60 ? phv_data_54 : _GEN_4806; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4808 = 14'h37 == parameter_2_60 ? phv_data_55 : _GEN_4807; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4809 = 14'h38 == parameter_2_60 ? phv_data_56 : _GEN_4808; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4810 = 14'h39 == parameter_2_60 ? phv_data_57 : _GEN_4809; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4811 = 14'h3a == parameter_2_60 ? phv_data_58 : _GEN_4810; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4812 = 14'h3b == parameter_2_60 ? phv_data_59 : _GEN_4811; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4813 = 14'h3c == parameter_2_60 ? phv_data_60 : _GEN_4812; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4814 = 14'h3d == parameter_2_60 ? phv_data_61 : _GEN_4813; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4815 = 14'h3e == parameter_2_60 ? phv_data_62 : _GEN_4814; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4816 = 14'h3f == parameter_2_60 ? phv_data_63 : _GEN_4815; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_61 = vliw_61[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_61 = vliw_61[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_61 = parameter_2_61[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_61 = parameter_2_61[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_61 = {{1'd0}, args_offset_61}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_61 = _total_offset_T_61[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_4820 = 3'h1 == total_offset_61 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4821 = 3'h2 == total_offset_61 ? args_2 : _GEN_4820; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4822 = 3'h3 == total_offset_61 ? args_3 : _GEN_4821; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4823 = 3'h4 == total_offset_61 ? args_4 : _GEN_4822; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4824 = 3'h5 == total_offset_61 ? args_5 : _GEN_4823; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4825 = 3'h6 == total_offset_61 ? args_6 : _GEN_4824; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4826 = total_offset_61 < 3'h7 ? _GEN_4825 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_61_0 = 3'h0 < args_length_61 ? _GEN_4826 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_4828 = opcode_61 == 4'ha ? field_bytes_61_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_4829 = opcode_61 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_4334 = opcode_61 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_123 = _T_4334 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_4830 = opcode_61 == 4'h8 | opcode_61 == 4'hb ? parameter_2_61[7:0] : _GEN_4828; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_4831 = opcode_61 == 4'h8 | opcode_61 == 4'hb ? _field_tag_T_123 : _GEN_4829; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_4832 = 14'h0 == parameter_2_61 ? phv_data_0 : _GEN_4830; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4833 = 14'h1 == parameter_2_61 ? phv_data_1 : _GEN_4832; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4834 = 14'h2 == parameter_2_61 ? phv_data_2 : _GEN_4833; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4835 = 14'h3 == parameter_2_61 ? phv_data_3 : _GEN_4834; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4836 = 14'h4 == parameter_2_61 ? phv_data_4 : _GEN_4835; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4837 = 14'h5 == parameter_2_61 ? phv_data_5 : _GEN_4836; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4838 = 14'h6 == parameter_2_61 ? phv_data_6 : _GEN_4837; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4839 = 14'h7 == parameter_2_61 ? phv_data_7 : _GEN_4838; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4840 = 14'h8 == parameter_2_61 ? phv_data_8 : _GEN_4839; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4841 = 14'h9 == parameter_2_61 ? phv_data_9 : _GEN_4840; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4842 = 14'ha == parameter_2_61 ? phv_data_10 : _GEN_4841; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4843 = 14'hb == parameter_2_61 ? phv_data_11 : _GEN_4842; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4844 = 14'hc == parameter_2_61 ? phv_data_12 : _GEN_4843; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4845 = 14'hd == parameter_2_61 ? phv_data_13 : _GEN_4844; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4846 = 14'he == parameter_2_61 ? phv_data_14 : _GEN_4845; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4847 = 14'hf == parameter_2_61 ? phv_data_15 : _GEN_4846; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4848 = 14'h10 == parameter_2_61 ? phv_data_16 : _GEN_4847; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4849 = 14'h11 == parameter_2_61 ? phv_data_17 : _GEN_4848; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4850 = 14'h12 == parameter_2_61 ? phv_data_18 : _GEN_4849; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4851 = 14'h13 == parameter_2_61 ? phv_data_19 : _GEN_4850; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4852 = 14'h14 == parameter_2_61 ? phv_data_20 : _GEN_4851; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4853 = 14'h15 == parameter_2_61 ? phv_data_21 : _GEN_4852; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4854 = 14'h16 == parameter_2_61 ? phv_data_22 : _GEN_4853; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4855 = 14'h17 == parameter_2_61 ? phv_data_23 : _GEN_4854; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4856 = 14'h18 == parameter_2_61 ? phv_data_24 : _GEN_4855; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4857 = 14'h19 == parameter_2_61 ? phv_data_25 : _GEN_4856; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4858 = 14'h1a == parameter_2_61 ? phv_data_26 : _GEN_4857; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4859 = 14'h1b == parameter_2_61 ? phv_data_27 : _GEN_4858; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4860 = 14'h1c == parameter_2_61 ? phv_data_28 : _GEN_4859; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4861 = 14'h1d == parameter_2_61 ? phv_data_29 : _GEN_4860; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4862 = 14'h1e == parameter_2_61 ? phv_data_30 : _GEN_4861; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4863 = 14'h1f == parameter_2_61 ? phv_data_31 : _GEN_4862; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4864 = 14'h20 == parameter_2_61 ? phv_data_32 : _GEN_4863; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4865 = 14'h21 == parameter_2_61 ? phv_data_33 : _GEN_4864; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4866 = 14'h22 == parameter_2_61 ? phv_data_34 : _GEN_4865; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4867 = 14'h23 == parameter_2_61 ? phv_data_35 : _GEN_4866; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4868 = 14'h24 == parameter_2_61 ? phv_data_36 : _GEN_4867; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4869 = 14'h25 == parameter_2_61 ? phv_data_37 : _GEN_4868; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4870 = 14'h26 == parameter_2_61 ? phv_data_38 : _GEN_4869; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4871 = 14'h27 == parameter_2_61 ? phv_data_39 : _GEN_4870; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4872 = 14'h28 == parameter_2_61 ? phv_data_40 : _GEN_4871; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4873 = 14'h29 == parameter_2_61 ? phv_data_41 : _GEN_4872; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4874 = 14'h2a == parameter_2_61 ? phv_data_42 : _GEN_4873; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4875 = 14'h2b == parameter_2_61 ? phv_data_43 : _GEN_4874; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4876 = 14'h2c == parameter_2_61 ? phv_data_44 : _GEN_4875; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4877 = 14'h2d == parameter_2_61 ? phv_data_45 : _GEN_4876; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4878 = 14'h2e == parameter_2_61 ? phv_data_46 : _GEN_4877; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4879 = 14'h2f == parameter_2_61 ? phv_data_47 : _GEN_4878; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4880 = 14'h30 == parameter_2_61 ? phv_data_48 : _GEN_4879; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4881 = 14'h31 == parameter_2_61 ? phv_data_49 : _GEN_4880; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4882 = 14'h32 == parameter_2_61 ? phv_data_50 : _GEN_4881; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4883 = 14'h33 == parameter_2_61 ? phv_data_51 : _GEN_4882; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4884 = 14'h34 == parameter_2_61 ? phv_data_52 : _GEN_4883; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4885 = 14'h35 == parameter_2_61 ? phv_data_53 : _GEN_4884; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4886 = 14'h36 == parameter_2_61 ? phv_data_54 : _GEN_4885; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4887 = 14'h37 == parameter_2_61 ? phv_data_55 : _GEN_4886; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4888 = 14'h38 == parameter_2_61 ? phv_data_56 : _GEN_4887; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4889 = 14'h39 == parameter_2_61 ? phv_data_57 : _GEN_4888; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4890 = 14'h3a == parameter_2_61 ? phv_data_58 : _GEN_4889; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4891 = 14'h3b == parameter_2_61 ? phv_data_59 : _GEN_4890; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4892 = 14'h3c == parameter_2_61 ? phv_data_60 : _GEN_4891; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4893 = 14'h3d == parameter_2_61 ? phv_data_61 : _GEN_4892; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4894 = 14'h3e == parameter_2_61 ? phv_data_62 : _GEN_4893; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4895 = 14'h3f == parameter_2_61 ? phv_data_63 : _GEN_4894; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_62 = vliw_62[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_62 = vliw_62[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_62 = parameter_2_62[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_62 = parameter_2_62[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_62 = {{1'd0}, args_offset_62}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_62 = _total_offset_T_62[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_4899 = 3'h1 == total_offset_62 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4900 = 3'h2 == total_offset_62 ? args_2 : _GEN_4899; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4901 = 3'h3 == total_offset_62 ? args_3 : _GEN_4900; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4902 = 3'h4 == total_offset_62 ? args_4 : _GEN_4901; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4903 = 3'h5 == total_offset_62 ? args_5 : _GEN_4902; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4904 = 3'h6 == total_offset_62 ? args_6 : _GEN_4903; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4905 = total_offset_62 < 3'h7 ? _GEN_4904 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_62_0 = 3'h0 < args_length_62 ? _GEN_4905 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_4907 = opcode_62 == 4'ha ? field_bytes_62_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_4908 = opcode_62 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_4405 = opcode_62 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_125 = _T_4405 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_4909 = opcode_62 == 4'h8 | opcode_62 == 4'hb ? parameter_2_62[7:0] : _GEN_4907; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_4910 = opcode_62 == 4'h8 | opcode_62 == 4'hb ? _field_tag_T_125 : _GEN_4908; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_4911 = 14'h0 == parameter_2_62 ? phv_data_0 : _GEN_4909; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4912 = 14'h1 == parameter_2_62 ? phv_data_1 : _GEN_4911; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4913 = 14'h2 == parameter_2_62 ? phv_data_2 : _GEN_4912; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4914 = 14'h3 == parameter_2_62 ? phv_data_3 : _GEN_4913; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4915 = 14'h4 == parameter_2_62 ? phv_data_4 : _GEN_4914; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4916 = 14'h5 == parameter_2_62 ? phv_data_5 : _GEN_4915; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4917 = 14'h6 == parameter_2_62 ? phv_data_6 : _GEN_4916; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4918 = 14'h7 == parameter_2_62 ? phv_data_7 : _GEN_4917; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4919 = 14'h8 == parameter_2_62 ? phv_data_8 : _GEN_4918; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4920 = 14'h9 == parameter_2_62 ? phv_data_9 : _GEN_4919; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4921 = 14'ha == parameter_2_62 ? phv_data_10 : _GEN_4920; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4922 = 14'hb == parameter_2_62 ? phv_data_11 : _GEN_4921; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4923 = 14'hc == parameter_2_62 ? phv_data_12 : _GEN_4922; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4924 = 14'hd == parameter_2_62 ? phv_data_13 : _GEN_4923; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4925 = 14'he == parameter_2_62 ? phv_data_14 : _GEN_4924; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4926 = 14'hf == parameter_2_62 ? phv_data_15 : _GEN_4925; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4927 = 14'h10 == parameter_2_62 ? phv_data_16 : _GEN_4926; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4928 = 14'h11 == parameter_2_62 ? phv_data_17 : _GEN_4927; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4929 = 14'h12 == parameter_2_62 ? phv_data_18 : _GEN_4928; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4930 = 14'h13 == parameter_2_62 ? phv_data_19 : _GEN_4929; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4931 = 14'h14 == parameter_2_62 ? phv_data_20 : _GEN_4930; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4932 = 14'h15 == parameter_2_62 ? phv_data_21 : _GEN_4931; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4933 = 14'h16 == parameter_2_62 ? phv_data_22 : _GEN_4932; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4934 = 14'h17 == parameter_2_62 ? phv_data_23 : _GEN_4933; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4935 = 14'h18 == parameter_2_62 ? phv_data_24 : _GEN_4934; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4936 = 14'h19 == parameter_2_62 ? phv_data_25 : _GEN_4935; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4937 = 14'h1a == parameter_2_62 ? phv_data_26 : _GEN_4936; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4938 = 14'h1b == parameter_2_62 ? phv_data_27 : _GEN_4937; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4939 = 14'h1c == parameter_2_62 ? phv_data_28 : _GEN_4938; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4940 = 14'h1d == parameter_2_62 ? phv_data_29 : _GEN_4939; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4941 = 14'h1e == parameter_2_62 ? phv_data_30 : _GEN_4940; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4942 = 14'h1f == parameter_2_62 ? phv_data_31 : _GEN_4941; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4943 = 14'h20 == parameter_2_62 ? phv_data_32 : _GEN_4942; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4944 = 14'h21 == parameter_2_62 ? phv_data_33 : _GEN_4943; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4945 = 14'h22 == parameter_2_62 ? phv_data_34 : _GEN_4944; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4946 = 14'h23 == parameter_2_62 ? phv_data_35 : _GEN_4945; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4947 = 14'h24 == parameter_2_62 ? phv_data_36 : _GEN_4946; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4948 = 14'h25 == parameter_2_62 ? phv_data_37 : _GEN_4947; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4949 = 14'h26 == parameter_2_62 ? phv_data_38 : _GEN_4948; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4950 = 14'h27 == parameter_2_62 ? phv_data_39 : _GEN_4949; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4951 = 14'h28 == parameter_2_62 ? phv_data_40 : _GEN_4950; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4952 = 14'h29 == parameter_2_62 ? phv_data_41 : _GEN_4951; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4953 = 14'h2a == parameter_2_62 ? phv_data_42 : _GEN_4952; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4954 = 14'h2b == parameter_2_62 ? phv_data_43 : _GEN_4953; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4955 = 14'h2c == parameter_2_62 ? phv_data_44 : _GEN_4954; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4956 = 14'h2d == parameter_2_62 ? phv_data_45 : _GEN_4955; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4957 = 14'h2e == parameter_2_62 ? phv_data_46 : _GEN_4956; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4958 = 14'h2f == parameter_2_62 ? phv_data_47 : _GEN_4957; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4959 = 14'h30 == parameter_2_62 ? phv_data_48 : _GEN_4958; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4960 = 14'h31 == parameter_2_62 ? phv_data_49 : _GEN_4959; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4961 = 14'h32 == parameter_2_62 ? phv_data_50 : _GEN_4960; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4962 = 14'h33 == parameter_2_62 ? phv_data_51 : _GEN_4961; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4963 = 14'h34 == parameter_2_62 ? phv_data_52 : _GEN_4962; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4964 = 14'h35 == parameter_2_62 ? phv_data_53 : _GEN_4963; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4965 = 14'h36 == parameter_2_62 ? phv_data_54 : _GEN_4964; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4966 = 14'h37 == parameter_2_62 ? phv_data_55 : _GEN_4965; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4967 = 14'h38 == parameter_2_62 ? phv_data_56 : _GEN_4966; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4968 = 14'h39 == parameter_2_62 ? phv_data_57 : _GEN_4967; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4969 = 14'h3a == parameter_2_62 ? phv_data_58 : _GEN_4968; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4970 = 14'h3b == parameter_2_62 ? phv_data_59 : _GEN_4969; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4971 = 14'h3c == parameter_2_62 ? phv_data_60 : _GEN_4970; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4972 = 14'h3d == parameter_2_62 ? phv_data_61 : _GEN_4971; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4973 = 14'h3e == parameter_2_62 ? phv_data_62 : _GEN_4972; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4974 = 14'h3f == parameter_2_62 ? phv_data_63 : _GEN_4973; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_63 = vliw_63[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_63 = vliw_63[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_63 = parameter_2_63[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_63 = parameter_2_63[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_63 = {{1'd0}, args_offset_63}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_63 = _total_offset_T_63[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_4978 = 3'h1 == total_offset_63 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4979 = 3'h2 == total_offset_63 ? args_2 : _GEN_4978; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4980 = 3'h3 == total_offset_63 ? args_3 : _GEN_4979; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4981 = 3'h4 == total_offset_63 ? args_4 : _GEN_4980; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4982 = 3'h5 == total_offset_63 ? args_5 : _GEN_4981; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4983 = 3'h6 == total_offset_63 ? args_6 : _GEN_4982; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4984 = total_offset_63 < 3'h7 ? _GEN_4983 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_63_0 = 3'h0 < args_length_63 ? _GEN_4984 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_4986 = opcode_63 == 4'ha ? field_bytes_63_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_4987 = opcode_63 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_4476 = opcode_63 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_127 = _T_4476 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_4988 = opcode_63 == 4'h8 | opcode_63 == 4'hb ? parameter_2_63[7:0] : _GEN_4986; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_4989 = opcode_63 == 4'h8 | opcode_63 == 4'hb ? _field_tag_T_127 : _GEN_4987; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_4990 = 14'h0 == parameter_2_63 ? phv_data_0 : _GEN_4988; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4991 = 14'h1 == parameter_2_63 ? phv_data_1 : _GEN_4990; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4992 = 14'h2 == parameter_2_63 ? phv_data_2 : _GEN_4991; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4993 = 14'h3 == parameter_2_63 ? phv_data_3 : _GEN_4992; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4994 = 14'h4 == parameter_2_63 ? phv_data_4 : _GEN_4993; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4995 = 14'h5 == parameter_2_63 ? phv_data_5 : _GEN_4994; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4996 = 14'h6 == parameter_2_63 ? phv_data_6 : _GEN_4995; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4997 = 14'h7 == parameter_2_63 ? phv_data_7 : _GEN_4996; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4998 = 14'h8 == parameter_2_63 ? phv_data_8 : _GEN_4997; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_4999 = 14'h9 == parameter_2_63 ? phv_data_9 : _GEN_4998; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5000 = 14'ha == parameter_2_63 ? phv_data_10 : _GEN_4999; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5001 = 14'hb == parameter_2_63 ? phv_data_11 : _GEN_5000; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5002 = 14'hc == parameter_2_63 ? phv_data_12 : _GEN_5001; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5003 = 14'hd == parameter_2_63 ? phv_data_13 : _GEN_5002; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5004 = 14'he == parameter_2_63 ? phv_data_14 : _GEN_5003; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5005 = 14'hf == parameter_2_63 ? phv_data_15 : _GEN_5004; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5006 = 14'h10 == parameter_2_63 ? phv_data_16 : _GEN_5005; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5007 = 14'h11 == parameter_2_63 ? phv_data_17 : _GEN_5006; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5008 = 14'h12 == parameter_2_63 ? phv_data_18 : _GEN_5007; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5009 = 14'h13 == parameter_2_63 ? phv_data_19 : _GEN_5008; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5010 = 14'h14 == parameter_2_63 ? phv_data_20 : _GEN_5009; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5011 = 14'h15 == parameter_2_63 ? phv_data_21 : _GEN_5010; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5012 = 14'h16 == parameter_2_63 ? phv_data_22 : _GEN_5011; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5013 = 14'h17 == parameter_2_63 ? phv_data_23 : _GEN_5012; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5014 = 14'h18 == parameter_2_63 ? phv_data_24 : _GEN_5013; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5015 = 14'h19 == parameter_2_63 ? phv_data_25 : _GEN_5014; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5016 = 14'h1a == parameter_2_63 ? phv_data_26 : _GEN_5015; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5017 = 14'h1b == parameter_2_63 ? phv_data_27 : _GEN_5016; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5018 = 14'h1c == parameter_2_63 ? phv_data_28 : _GEN_5017; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5019 = 14'h1d == parameter_2_63 ? phv_data_29 : _GEN_5018; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5020 = 14'h1e == parameter_2_63 ? phv_data_30 : _GEN_5019; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5021 = 14'h1f == parameter_2_63 ? phv_data_31 : _GEN_5020; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5022 = 14'h20 == parameter_2_63 ? phv_data_32 : _GEN_5021; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5023 = 14'h21 == parameter_2_63 ? phv_data_33 : _GEN_5022; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5024 = 14'h22 == parameter_2_63 ? phv_data_34 : _GEN_5023; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5025 = 14'h23 == parameter_2_63 ? phv_data_35 : _GEN_5024; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5026 = 14'h24 == parameter_2_63 ? phv_data_36 : _GEN_5025; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5027 = 14'h25 == parameter_2_63 ? phv_data_37 : _GEN_5026; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5028 = 14'h26 == parameter_2_63 ? phv_data_38 : _GEN_5027; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5029 = 14'h27 == parameter_2_63 ? phv_data_39 : _GEN_5028; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5030 = 14'h28 == parameter_2_63 ? phv_data_40 : _GEN_5029; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5031 = 14'h29 == parameter_2_63 ? phv_data_41 : _GEN_5030; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5032 = 14'h2a == parameter_2_63 ? phv_data_42 : _GEN_5031; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5033 = 14'h2b == parameter_2_63 ? phv_data_43 : _GEN_5032; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5034 = 14'h2c == parameter_2_63 ? phv_data_44 : _GEN_5033; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5035 = 14'h2d == parameter_2_63 ? phv_data_45 : _GEN_5034; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5036 = 14'h2e == parameter_2_63 ? phv_data_46 : _GEN_5035; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5037 = 14'h2f == parameter_2_63 ? phv_data_47 : _GEN_5036; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5038 = 14'h30 == parameter_2_63 ? phv_data_48 : _GEN_5037; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5039 = 14'h31 == parameter_2_63 ? phv_data_49 : _GEN_5038; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5040 = 14'h32 == parameter_2_63 ? phv_data_50 : _GEN_5039; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5041 = 14'h33 == parameter_2_63 ? phv_data_51 : _GEN_5040; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5042 = 14'h34 == parameter_2_63 ? phv_data_52 : _GEN_5041; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5043 = 14'h35 == parameter_2_63 ? phv_data_53 : _GEN_5042; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5044 = 14'h36 == parameter_2_63 ? phv_data_54 : _GEN_5043; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5045 = 14'h37 == parameter_2_63 ? phv_data_55 : _GEN_5044; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5046 = 14'h38 == parameter_2_63 ? phv_data_56 : _GEN_5045; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5047 = 14'h39 == parameter_2_63 ? phv_data_57 : _GEN_5046; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5048 = 14'h3a == parameter_2_63 ? phv_data_58 : _GEN_5047; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5049 = 14'h3b == parameter_2_63 ? phv_data_59 : _GEN_5048; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5050 = 14'h3c == parameter_2_63 ? phv_data_60 : _GEN_5049; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5051 = 14'h3d == parameter_2_63 ? phv_data_61 : _GEN_5050; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5052 = 14'h3e == parameter_2_63 ? phv_data_62 : _GEN_5051; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_5053 = 14'h3f == parameter_2_63 ? phv_data_63 : _GEN_5052; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_64 = vliw_64[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo = vliw_64[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_64 = field_data_lo[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_64 = field_data_lo[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_64 = {{1'd0}, args_offset_64}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_64 = _total_offset_T_64[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_5057 = 3'h1 == total_offset_64 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5058 = 3'h2 == total_offset_64 ? args_2 : _GEN_5057; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5059 = 3'h3 == total_offset_64 ? args_3 : _GEN_5058; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5060 = 3'h4 == total_offset_64 ? args_4 : _GEN_5059; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5061 = 3'h5 == total_offset_64 ? args_5 : _GEN_5060; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5062 = 3'h6 == total_offset_64 ? args_6 : _GEN_5061; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5063 = total_offset_64 < 3'h7 ? _GEN_5062 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_64_1 = 3'h0 < args_length_64 ? _GEN_5063 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_65 = args_offset_64 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_5066 = 3'h1 == total_offset_65 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5067 = 3'h2 == total_offset_65 ? args_2 : _GEN_5066; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5068 = 3'h3 == total_offset_65 ? args_3 : _GEN_5067; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5069 = 3'h4 == total_offset_65 ? args_4 : _GEN_5068; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5070 = 3'h5 == total_offset_65 ? args_5 : _GEN_5069; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5071 = 3'h6 == total_offset_65 ? args_6 : _GEN_5070; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5072 = total_offset_65 < 3'h7 ? _GEN_5071 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_64_0 = 3'h1 < args_length_64 ? _GEN_5072 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_64 = {field_bytes_64_0,field_bytes_64_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5074 = opcode_64 == 4'ha ? _field_data_T_64 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_5075 = opcode_64 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_4549 = opcode_64 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi = field_data_lo[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_67 = {field_data_hi,field_data_lo}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_129 = _T_4549 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_5076 = opcode_64 == 4'h8 | opcode_64 == 4'hb ? _field_data_T_67 : _GEN_5074; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_5077 = opcode_64 == 4'h8 | opcode_64 == 4'hb ? _field_tag_T_129 : _GEN_5075; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _field_data_T_68 = {phv_data_64,phv_data_65}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5078 = 14'h40 == field_data_lo ? _field_data_T_68 : _GEN_5076; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_69 = {phv_data_66,phv_data_67}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5079 = 14'h41 == field_data_lo ? _field_data_T_69 : _GEN_5078; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_70 = {phv_data_68,phv_data_69}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5080 = 14'h42 == field_data_lo ? _field_data_T_70 : _GEN_5079; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_71 = {phv_data_70,phv_data_71}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5081 = 14'h43 == field_data_lo ? _field_data_T_71 : _GEN_5080; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_72 = {phv_data_72,phv_data_73}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5082 = 14'h44 == field_data_lo ? _field_data_T_72 : _GEN_5081; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_73 = {phv_data_74,phv_data_75}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5083 = 14'h45 == field_data_lo ? _field_data_T_73 : _GEN_5082; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_74 = {phv_data_76,phv_data_77}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5084 = 14'h46 == field_data_lo ? _field_data_T_74 : _GEN_5083; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_75 = {phv_data_78,phv_data_79}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5085 = 14'h47 == field_data_lo ? _field_data_T_75 : _GEN_5084; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_76 = {phv_data_80,phv_data_81}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5086 = 14'h48 == field_data_lo ? _field_data_T_76 : _GEN_5085; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_77 = {phv_data_82,phv_data_83}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5087 = 14'h49 == field_data_lo ? _field_data_T_77 : _GEN_5086; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_78 = {phv_data_84,phv_data_85}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5088 = 14'h4a == field_data_lo ? _field_data_T_78 : _GEN_5087; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_79 = {phv_data_86,phv_data_87}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5089 = 14'h4b == field_data_lo ? _field_data_T_79 : _GEN_5088; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_80 = {phv_data_88,phv_data_89}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5090 = 14'h4c == field_data_lo ? _field_data_T_80 : _GEN_5089; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_81 = {phv_data_90,phv_data_91}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5091 = 14'h4d == field_data_lo ? _field_data_T_81 : _GEN_5090; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_82 = {phv_data_92,phv_data_93}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5092 = 14'h4e == field_data_lo ? _field_data_T_82 : _GEN_5091; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_83 = {phv_data_94,phv_data_95}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5093 = 14'h4f == field_data_lo ? _field_data_T_83 : _GEN_5092; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_84 = {phv_data_96,phv_data_97}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5094 = 14'h50 == field_data_lo ? _field_data_T_84 : _GEN_5093; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_85 = {phv_data_98,phv_data_99}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5095 = 14'h51 == field_data_lo ? _field_data_T_85 : _GEN_5094; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_86 = {phv_data_100,phv_data_101}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5096 = 14'h52 == field_data_lo ? _field_data_T_86 : _GEN_5095; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_87 = {phv_data_102,phv_data_103}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5097 = 14'h53 == field_data_lo ? _field_data_T_87 : _GEN_5096; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_88 = {phv_data_104,phv_data_105}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5098 = 14'h54 == field_data_lo ? _field_data_T_88 : _GEN_5097; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_89 = {phv_data_106,phv_data_107}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5099 = 14'h55 == field_data_lo ? _field_data_T_89 : _GEN_5098; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_90 = {phv_data_108,phv_data_109}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5100 = 14'h56 == field_data_lo ? _field_data_T_90 : _GEN_5099; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_91 = {phv_data_110,phv_data_111}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5101 = 14'h57 == field_data_lo ? _field_data_T_91 : _GEN_5100; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_92 = {phv_data_112,phv_data_113}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5102 = 14'h58 == field_data_lo ? _field_data_T_92 : _GEN_5101; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_93 = {phv_data_114,phv_data_115}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5103 = 14'h59 == field_data_lo ? _field_data_T_93 : _GEN_5102; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_94 = {phv_data_116,phv_data_117}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5104 = 14'h5a == field_data_lo ? _field_data_T_94 : _GEN_5103; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_95 = {phv_data_118,phv_data_119}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5105 = 14'h5b == field_data_lo ? _field_data_T_95 : _GEN_5104; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_96 = {phv_data_120,phv_data_121}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5106 = 14'h5c == field_data_lo ? _field_data_T_96 : _GEN_5105; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_97 = {phv_data_122,phv_data_123}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5107 = 14'h5d == field_data_lo ? _field_data_T_97 : _GEN_5106; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_98 = {phv_data_124,phv_data_125}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5108 = 14'h5e == field_data_lo ? _field_data_T_98 : _GEN_5107; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_99 = {phv_data_126,phv_data_127}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5109 = 14'h5f == field_data_lo ? _field_data_T_99 : _GEN_5108; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_100 = {phv_data_128,phv_data_129}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5110 = 14'h60 == field_data_lo ? _field_data_T_100 : _GEN_5109; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_101 = {phv_data_130,phv_data_131}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5111 = 14'h61 == field_data_lo ? _field_data_T_101 : _GEN_5110; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_102 = {phv_data_132,phv_data_133}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5112 = 14'h62 == field_data_lo ? _field_data_T_102 : _GEN_5111; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_103 = {phv_data_134,phv_data_135}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5113 = 14'h63 == field_data_lo ? _field_data_T_103 : _GEN_5112; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_104 = {phv_data_136,phv_data_137}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5114 = 14'h64 == field_data_lo ? _field_data_T_104 : _GEN_5113; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_105 = {phv_data_138,phv_data_139}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5115 = 14'h65 == field_data_lo ? _field_data_T_105 : _GEN_5114; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_106 = {phv_data_140,phv_data_141}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5116 = 14'h66 == field_data_lo ? _field_data_T_106 : _GEN_5115; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_107 = {phv_data_142,phv_data_143}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5117 = 14'h67 == field_data_lo ? _field_data_T_107 : _GEN_5116; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_108 = {phv_data_144,phv_data_145}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5118 = 14'h68 == field_data_lo ? _field_data_T_108 : _GEN_5117; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_109 = {phv_data_146,phv_data_147}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5119 = 14'h69 == field_data_lo ? _field_data_T_109 : _GEN_5118; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_110 = {phv_data_148,phv_data_149}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5120 = 14'h6a == field_data_lo ? _field_data_T_110 : _GEN_5119; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_111 = {phv_data_150,phv_data_151}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5121 = 14'h6b == field_data_lo ? _field_data_T_111 : _GEN_5120; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_112 = {phv_data_152,phv_data_153}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5122 = 14'h6c == field_data_lo ? _field_data_T_112 : _GEN_5121; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_113 = {phv_data_154,phv_data_155}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5123 = 14'h6d == field_data_lo ? _field_data_T_113 : _GEN_5122; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_114 = {phv_data_156,phv_data_157}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5124 = 14'h6e == field_data_lo ? _field_data_T_114 : _GEN_5123; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_115 = {phv_data_158,phv_data_159}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5125 = 14'h6f == field_data_lo ? _field_data_T_115 : _GEN_5124; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_116 = {phv_data_160,phv_data_161}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5126 = 14'h70 == field_data_lo ? _field_data_T_116 : _GEN_5125; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_117 = {phv_data_162,phv_data_163}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5127 = 14'h71 == field_data_lo ? _field_data_T_117 : _GEN_5126; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_118 = {phv_data_164,phv_data_165}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5128 = 14'h72 == field_data_lo ? _field_data_T_118 : _GEN_5127; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_119 = {phv_data_166,phv_data_167}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5129 = 14'h73 == field_data_lo ? _field_data_T_119 : _GEN_5128; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_120 = {phv_data_168,phv_data_169}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5130 = 14'h74 == field_data_lo ? _field_data_T_120 : _GEN_5129; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_121 = {phv_data_170,phv_data_171}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5131 = 14'h75 == field_data_lo ? _field_data_T_121 : _GEN_5130; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_122 = {phv_data_172,phv_data_173}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5132 = 14'h76 == field_data_lo ? _field_data_T_122 : _GEN_5131; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_123 = {phv_data_174,phv_data_175}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5133 = 14'h77 == field_data_lo ? _field_data_T_123 : _GEN_5132; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_124 = {phv_data_176,phv_data_177}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5134 = 14'h78 == field_data_lo ? _field_data_T_124 : _GEN_5133; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_125 = {phv_data_178,phv_data_179}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5135 = 14'h79 == field_data_lo ? _field_data_T_125 : _GEN_5134; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_126 = {phv_data_180,phv_data_181}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5136 = 14'h7a == field_data_lo ? _field_data_T_126 : _GEN_5135; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_127 = {phv_data_182,phv_data_183}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5137 = 14'h7b == field_data_lo ? _field_data_T_127 : _GEN_5136; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_128 = {phv_data_184,phv_data_185}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5138 = 14'h7c == field_data_lo ? _field_data_T_128 : _GEN_5137; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_129 = {phv_data_186,phv_data_187}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5139 = 14'h7d == field_data_lo ? _field_data_T_129 : _GEN_5138; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_130 = {phv_data_188,phv_data_189}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5140 = 14'h7e == field_data_lo ? _field_data_T_130 : _GEN_5139; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_131 = {phv_data_190,phv_data_191}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5141 = 14'h7f == field_data_lo ? _field_data_T_131 : _GEN_5140; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_132 = {phv_data_192,phv_data_193}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5142 = 14'h80 == field_data_lo ? _field_data_T_132 : _GEN_5141; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_133 = {phv_data_194,phv_data_195}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5143 = 14'h81 == field_data_lo ? _field_data_T_133 : _GEN_5142; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_134 = {phv_data_196,phv_data_197}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5144 = 14'h82 == field_data_lo ? _field_data_T_134 : _GEN_5143; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_135 = {phv_data_198,phv_data_199}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5145 = 14'h83 == field_data_lo ? _field_data_T_135 : _GEN_5144; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_136 = {phv_data_200,phv_data_201}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5146 = 14'h84 == field_data_lo ? _field_data_T_136 : _GEN_5145; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_137 = {phv_data_202,phv_data_203}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5147 = 14'h85 == field_data_lo ? _field_data_T_137 : _GEN_5146; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_138 = {phv_data_204,phv_data_205}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5148 = 14'h86 == field_data_lo ? _field_data_T_138 : _GEN_5147; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_139 = {phv_data_206,phv_data_207}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5149 = 14'h87 == field_data_lo ? _field_data_T_139 : _GEN_5148; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_140 = {phv_data_208,phv_data_209}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5150 = 14'h88 == field_data_lo ? _field_data_T_140 : _GEN_5149; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_141 = {phv_data_210,phv_data_211}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5151 = 14'h89 == field_data_lo ? _field_data_T_141 : _GEN_5150; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_142 = {phv_data_212,phv_data_213}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5152 = 14'h8a == field_data_lo ? _field_data_T_142 : _GEN_5151; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_143 = {phv_data_214,phv_data_215}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5153 = 14'h8b == field_data_lo ? _field_data_T_143 : _GEN_5152; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_144 = {phv_data_216,phv_data_217}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5154 = 14'h8c == field_data_lo ? _field_data_T_144 : _GEN_5153; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_145 = {phv_data_218,phv_data_219}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5155 = 14'h8d == field_data_lo ? _field_data_T_145 : _GEN_5154; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_146 = {phv_data_220,phv_data_221}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5156 = 14'h8e == field_data_lo ? _field_data_T_146 : _GEN_5155; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_147 = {phv_data_222,phv_data_223}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5157 = 14'h8f == field_data_lo ? _field_data_T_147 : _GEN_5156; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_148 = {phv_data_224,phv_data_225}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5158 = 14'h90 == field_data_lo ? _field_data_T_148 : _GEN_5157; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_149 = {phv_data_226,phv_data_227}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5159 = 14'h91 == field_data_lo ? _field_data_T_149 : _GEN_5158; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_150 = {phv_data_228,phv_data_229}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5160 = 14'h92 == field_data_lo ? _field_data_T_150 : _GEN_5159; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_151 = {phv_data_230,phv_data_231}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5161 = 14'h93 == field_data_lo ? _field_data_T_151 : _GEN_5160; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_152 = {phv_data_232,phv_data_233}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5162 = 14'h94 == field_data_lo ? _field_data_T_152 : _GEN_5161; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_153 = {phv_data_234,phv_data_235}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5163 = 14'h95 == field_data_lo ? _field_data_T_153 : _GEN_5162; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_154 = {phv_data_236,phv_data_237}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5164 = 14'h96 == field_data_lo ? _field_data_T_154 : _GEN_5163; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_155 = {phv_data_238,phv_data_239}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5165 = 14'h97 == field_data_lo ? _field_data_T_155 : _GEN_5164; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_156 = {phv_data_240,phv_data_241}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5166 = 14'h98 == field_data_lo ? _field_data_T_156 : _GEN_5165; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_157 = {phv_data_242,phv_data_243}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5167 = 14'h99 == field_data_lo ? _field_data_T_157 : _GEN_5166; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_158 = {phv_data_244,phv_data_245}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5168 = 14'h9a == field_data_lo ? _field_data_T_158 : _GEN_5167; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_159 = {phv_data_246,phv_data_247}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5169 = 14'h9b == field_data_lo ? _field_data_T_159 : _GEN_5168; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_160 = {phv_data_248,phv_data_249}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5170 = 14'h9c == field_data_lo ? _field_data_T_160 : _GEN_5169; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_161 = {phv_data_250,phv_data_251}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5171 = 14'h9d == field_data_lo ? _field_data_T_161 : _GEN_5170; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_162 = {phv_data_252,phv_data_253}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5172 = 14'h9e == field_data_lo ? _field_data_T_162 : _GEN_5171; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_163 = {phv_data_254,phv_data_255}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5173 = 14'h9f == field_data_lo ? _field_data_T_163 : _GEN_5172; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_65 = vliw_65[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_1 = vliw_65[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_65 = field_data_lo_1[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_65 = field_data_lo_1[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_66 = {{1'd0}, args_offset_65}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_66 = _total_offset_T_66[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_5177 = 3'h1 == total_offset_66 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5178 = 3'h2 == total_offset_66 ? args_2 : _GEN_5177; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5179 = 3'h3 == total_offset_66 ? args_3 : _GEN_5178; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5180 = 3'h4 == total_offset_66 ? args_4 : _GEN_5179; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5181 = 3'h5 == total_offset_66 ? args_5 : _GEN_5180; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5182 = 3'h6 == total_offset_66 ? args_6 : _GEN_5181; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5183 = total_offset_66 < 3'h7 ? _GEN_5182 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_65_1 = 3'h0 < args_length_65 ? _GEN_5183 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_67 = args_offset_65 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_5186 = 3'h1 == total_offset_67 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5187 = 3'h2 == total_offset_67 ? args_2 : _GEN_5186; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5188 = 3'h3 == total_offset_67 ? args_3 : _GEN_5187; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5189 = 3'h4 == total_offset_67 ? args_4 : _GEN_5188; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5190 = 3'h5 == total_offset_67 ? args_5 : _GEN_5189; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5191 = 3'h6 == total_offset_67 ? args_6 : _GEN_5190; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5192 = total_offset_67 < 3'h7 ? _GEN_5191 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_65_0 = 3'h1 < args_length_65 ? _GEN_5192 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_164 = {field_bytes_65_0,field_bytes_65_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5194 = opcode_65 == 4'ha ? _field_data_T_164 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_5195 = opcode_65 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_4654 = opcode_65 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_1 = field_data_lo_1[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_167 = {field_data_hi_1,field_data_lo_1}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_131 = _T_4654 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_5196 = opcode_65 == 4'h8 | opcode_65 == 4'hb ? _field_data_T_167 : _GEN_5194; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_5197 = opcode_65 == 4'h8 | opcode_65 == 4'hb ? _field_tag_T_131 : _GEN_5195; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_5198 = 14'h40 == field_data_lo_1 ? _field_data_T_68 : _GEN_5196; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5199 = 14'h41 == field_data_lo_1 ? _field_data_T_69 : _GEN_5198; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5200 = 14'h42 == field_data_lo_1 ? _field_data_T_70 : _GEN_5199; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5201 = 14'h43 == field_data_lo_1 ? _field_data_T_71 : _GEN_5200; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5202 = 14'h44 == field_data_lo_1 ? _field_data_T_72 : _GEN_5201; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5203 = 14'h45 == field_data_lo_1 ? _field_data_T_73 : _GEN_5202; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5204 = 14'h46 == field_data_lo_1 ? _field_data_T_74 : _GEN_5203; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5205 = 14'h47 == field_data_lo_1 ? _field_data_T_75 : _GEN_5204; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5206 = 14'h48 == field_data_lo_1 ? _field_data_T_76 : _GEN_5205; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5207 = 14'h49 == field_data_lo_1 ? _field_data_T_77 : _GEN_5206; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5208 = 14'h4a == field_data_lo_1 ? _field_data_T_78 : _GEN_5207; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5209 = 14'h4b == field_data_lo_1 ? _field_data_T_79 : _GEN_5208; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5210 = 14'h4c == field_data_lo_1 ? _field_data_T_80 : _GEN_5209; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5211 = 14'h4d == field_data_lo_1 ? _field_data_T_81 : _GEN_5210; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5212 = 14'h4e == field_data_lo_1 ? _field_data_T_82 : _GEN_5211; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5213 = 14'h4f == field_data_lo_1 ? _field_data_T_83 : _GEN_5212; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5214 = 14'h50 == field_data_lo_1 ? _field_data_T_84 : _GEN_5213; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5215 = 14'h51 == field_data_lo_1 ? _field_data_T_85 : _GEN_5214; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5216 = 14'h52 == field_data_lo_1 ? _field_data_T_86 : _GEN_5215; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5217 = 14'h53 == field_data_lo_1 ? _field_data_T_87 : _GEN_5216; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5218 = 14'h54 == field_data_lo_1 ? _field_data_T_88 : _GEN_5217; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5219 = 14'h55 == field_data_lo_1 ? _field_data_T_89 : _GEN_5218; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5220 = 14'h56 == field_data_lo_1 ? _field_data_T_90 : _GEN_5219; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5221 = 14'h57 == field_data_lo_1 ? _field_data_T_91 : _GEN_5220; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5222 = 14'h58 == field_data_lo_1 ? _field_data_T_92 : _GEN_5221; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5223 = 14'h59 == field_data_lo_1 ? _field_data_T_93 : _GEN_5222; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5224 = 14'h5a == field_data_lo_1 ? _field_data_T_94 : _GEN_5223; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5225 = 14'h5b == field_data_lo_1 ? _field_data_T_95 : _GEN_5224; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5226 = 14'h5c == field_data_lo_1 ? _field_data_T_96 : _GEN_5225; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5227 = 14'h5d == field_data_lo_1 ? _field_data_T_97 : _GEN_5226; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5228 = 14'h5e == field_data_lo_1 ? _field_data_T_98 : _GEN_5227; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5229 = 14'h5f == field_data_lo_1 ? _field_data_T_99 : _GEN_5228; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5230 = 14'h60 == field_data_lo_1 ? _field_data_T_100 : _GEN_5229; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5231 = 14'h61 == field_data_lo_1 ? _field_data_T_101 : _GEN_5230; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5232 = 14'h62 == field_data_lo_1 ? _field_data_T_102 : _GEN_5231; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5233 = 14'h63 == field_data_lo_1 ? _field_data_T_103 : _GEN_5232; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5234 = 14'h64 == field_data_lo_1 ? _field_data_T_104 : _GEN_5233; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5235 = 14'h65 == field_data_lo_1 ? _field_data_T_105 : _GEN_5234; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5236 = 14'h66 == field_data_lo_1 ? _field_data_T_106 : _GEN_5235; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5237 = 14'h67 == field_data_lo_1 ? _field_data_T_107 : _GEN_5236; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5238 = 14'h68 == field_data_lo_1 ? _field_data_T_108 : _GEN_5237; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5239 = 14'h69 == field_data_lo_1 ? _field_data_T_109 : _GEN_5238; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5240 = 14'h6a == field_data_lo_1 ? _field_data_T_110 : _GEN_5239; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5241 = 14'h6b == field_data_lo_1 ? _field_data_T_111 : _GEN_5240; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5242 = 14'h6c == field_data_lo_1 ? _field_data_T_112 : _GEN_5241; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5243 = 14'h6d == field_data_lo_1 ? _field_data_T_113 : _GEN_5242; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5244 = 14'h6e == field_data_lo_1 ? _field_data_T_114 : _GEN_5243; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5245 = 14'h6f == field_data_lo_1 ? _field_data_T_115 : _GEN_5244; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5246 = 14'h70 == field_data_lo_1 ? _field_data_T_116 : _GEN_5245; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5247 = 14'h71 == field_data_lo_1 ? _field_data_T_117 : _GEN_5246; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5248 = 14'h72 == field_data_lo_1 ? _field_data_T_118 : _GEN_5247; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5249 = 14'h73 == field_data_lo_1 ? _field_data_T_119 : _GEN_5248; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5250 = 14'h74 == field_data_lo_1 ? _field_data_T_120 : _GEN_5249; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5251 = 14'h75 == field_data_lo_1 ? _field_data_T_121 : _GEN_5250; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5252 = 14'h76 == field_data_lo_1 ? _field_data_T_122 : _GEN_5251; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5253 = 14'h77 == field_data_lo_1 ? _field_data_T_123 : _GEN_5252; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5254 = 14'h78 == field_data_lo_1 ? _field_data_T_124 : _GEN_5253; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5255 = 14'h79 == field_data_lo_1 ? _field_data_T_125 : _GEN_5254; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5256 = 14'h7a == field_data_lo_1 ? _field_data_T_126 : _GEN_5255; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5257 = 14'h7b == field_data_lo_1 ? _field_data_T_127 : _GEN_5256; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5258 = 14'h7c == field_data_lo_1 ? _field_data_T_128 : _GEN_5257; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5259 = 14'h7d == field_data_lo_1 ? _field_data_T_129 : _GEN_5258; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5260 = 14'h7e == field_data_lo_1 ? _field_data_T_130 : _GEN_5259; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5261 = 14'h7f == field_data_lo_1 ? _field_data_T_131 : _GEN_5260; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5262 = 14'h80 == field_data_lo_1 ? _field_data_T_132 : _GEN_5261; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5263 = 14'h81 == field_data_lo_1 ? _field_data_T_133 : _GEN_5262; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5264 = 14'h82 == field_data_lo_1 ? _field_data_T_134 : _GEN_5263; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5265 = 14'h83 == field_data_lo_1 ? _field_data_T_135 : _GEN_5264; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5266 = 14'h84 == field_data_lo_1 ? _field_data_T_136 : _GEN_5265; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5267 = 14'h85 == field_data_lo_1 ? _field_data_T_137 : _GEN_5266; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5268 = 14'h86 == field_data_lo_1 ? _field_data_T_138 : _GEN_5267; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5269 = 14'h87 == field_data_lo_1 ? _field_data_T_139 : _GEN_5268; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5270 = 14'h88 == field_data_lo_1 ? _field_data_T_140 : _GEN_5269; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5271 = 14'h89 == field_data_lo_1 ? _field_data_T_141 : _GEN_5270; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5272 = 14'h8a == field_data_lo_1 ? _field_data_T_142 : _GEN_5271; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5273 = 14'h8b == field_data_lo_1 ? _field_data_T_143 : _GEN_5272; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5274 = 14'h8c == field_data_lo_1 ? _field_data_T_144 : _GEN_5273; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5275 = 14'h8d == field_data_lo_1 ? _field_data_T_145 : _GEN_5274; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5276 = 14'h8e == field_data_lo_1 ? _field_data_T_146 : _GEN_5275; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5277 = 14'h8f == field_data_lo_1 ? _field_data_T_147 : _GEN_5276; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5278 = 14'h90 == field_data_lo_1 ? _field_data_T_148 : _GEN_5277; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5279 = 14'h91 == field_data_lo_1 ? _field_data_T_149 : _GEN_5278; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5280 = 14'h92 == field_data_lo_1 ? _field_data_T_150 : _GEN_5279; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5281 = 14'h93 == field_data_lo_1 ? _field_data_T_151 : _GEN_5280; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5282 = 14'h94 == field_data_lo_1 ? _field_data_T_152 : _GEN_5281; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5283 = 14'h95 == field_data_lo_1 ? _field_data_T_153 : _GEN_5282; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5284 = 14'h96 == field_data_lo_1 ? _field_data_T_154 : _GEN_5283; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5285 = 14'h97 == field_data_lo_1 ? _field_data_T_155 : _GEN_5284; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5286 = 14'h98 == field_data_lo_1 ? _field_data_T_156 : _GEN_5285; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5287 = 14'h99 == field_data_lo_1 ? _field_data_T_157 : _GEN_5286; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5288 = 14'h9a == field_data_lo_1 ? _field_data_T_158 : _GEN_5287; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5289 = 14'h9b == field_data_lo_1 ? _field_data_T_159 : _GEN_5288; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5290 = 14'h9c == field_data_lo_1 ? _field_data_T_160 : _GEN_5289; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5291 = 14'h9d == field_data_lo_1 ? _field_data_T_161 : _GEN_5290; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5292 = 14'h9e == field_data_lo_1 ? _field_data_T_162 : _GEN_5291; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5293 = 14'h9f == field_data_lo_1 ? _field_data_T_163 : _GEN_5292; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_66 = vliw_66[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_2 = vliw_66[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_66 = field_data_lo_2[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_66 = field_data_lo_2[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_68 = {{1'd0}, args_offset_66}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_68 = _total_offset_T_68[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_5297 = 3'h1 == total_offset_68 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5298 = 3'h2 == total_offset_68 ? args_2 : _GEN_5297; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5299 = 3'h3 == total_offset_68 ? args_3 : _GEN_5298; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5300 = 3'h4 == total_offset_68 ? args_4 : _GEN_5299; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5301 = 3'h5 == total_offset_68 ? args_5 : _GEN_5300; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5302 = 3'h6 == total_offset_68 ? args_6 : _GEN_5301; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5303 = total_offset_68 < 3'h7 ? _GEN_5302 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_66_1 = 3'h0 < args_length_66 ? _GEN_5303 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_69 = args_offset_66 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_5306 = 3'h1 == total_offset_69 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5307 = 3'h2 == total_offset_69 ? args_2 : _GEN_5306; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5308 = 3'h3 == total_offset_69 ? args_3 : _GEN_5307; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5309 = 3'h4 == total_offset_69 ? args_4 : _GEN_5308; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5310 = 3'h5 == total_offset_69 ? args_5 : _GEN_5309; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5311 = 3'h6 == total_offset_69 ? args_6 : _GEN_5310; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5312 = total_offset_69 < 3'h7 ? _GEN_5311 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_66_0 = 3'h1 < args_length_66 ? _GEN_5312 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_264 = {field_bytes_66_0,field_bytes_66_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5314 = opcode_66 == 4'ha ? _field_data_T_264 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_5315 = opcode_66 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_4759 = opcode_66 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_2 = field_data_lo_2[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_267 = {field_data_hi_2,field_data_lo_2}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_133 = _T_4759 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_5316 = opcode_66 == 4'h8 | opcode_66 == 4'hb ? _field_data_T_267 : _GEN_5314; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_5317 = opcode_66 == 4'h8 | opcode_66 == 4'hb ? _field_tag_T_133 : _GEN_5315; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_5318 = 14'h40 == field_data_lo_2 ? _field_data_T_68 : _GEN_5316; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5319 = 14'h41 == field_data_lo_2 ? _field_data_T_69 : _GEN_5318; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5320 = 14'h42 == field_data_lo_2 ? _field_data_T_70 : _GEN_5319; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5321 = 14'h43 == field_data_lo_2 ? _field_data_T_71 : _GEN_5320; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5322 = 14'h44 == field_data_lo_2 ? _field_data_T_72 : _GEN_5321; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5323 = 14'h45 == field_data_lo_2 ? _field_data_T_73 : _GEN_5322; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5324 = 14'h46 == field_data_lo_2 ? _field_data_T_74 : _GEN_5323; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5325 = 14'h47 == field_data_lo_2 ? _field_data_T_75 : _GEN_5324; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5326 = 14'h48 == field_data_lo_2 ? _field_data_T_76 : _GEN_5325; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5327 = 14'h49 == field_data_lo_2 ? _field_data_T_77 : _GEN_5326; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5328 = 14'h4a == field_data_lo_2 ? _field_data_T_78 : _GEN_5327; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5329 = 14'h4b == field_data_lo_2 ? _field_data_T_79 : _GEN_5328; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5330 = 14'h4c == field_data_lo_2 ? _field_data_T_80 : _GEN_5329; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5331 = 14'h4d == field_data_lo_2 ? _field_data_T_81 : _GEN_5330; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5332 = 14'h4e == field_data_lo_2 ? _field_data_T_82 : _GEN_5331; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5333 = 14'h4f == field_data_lo_2 ? _field_data_T_83 : _GEN_5332; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5334 = 14'h50 == field_data_lo_2 ? _field_data_T_84 : _GEN_5333; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5335 = 14'h51 == field_data_lo_2 ? _field_data_T_85 : _GEN_5334; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5336 = 14'h52 == field_data_lo_2 ? _field_data_T_86 : _GEN_5335; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5337 = 14'h53 == field_data_lo_2 ? _field_data_T_87 : _GEN_5336; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5338 = 14'h54 == field_data_lo_2 ? _field_data_T_88 : _GEN_5337; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5339 = 14'h55 == field_data_lo_2 ? _field_data_T_89 : _GEN_5338; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5340 = 14'h56 == field_data_lo_2 ? _field_data_T_90 : _GEN_5339; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5341 = 14'h57 == field_data_lo_2 ? _field_data_T_91 : _GEN_5340; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5342 = 14'h58 == field_data_lo_2 ? _field_data_T_92 : _GEN_5341; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5343 = 14'h59 == field_data_lo_2 ? _field_data_T_93 : _GEN_5342; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5344 = 14'h5a == field_data_lo_2 ? _field_data_T_94 : _GEN_5343; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5345 = 14'h5b == field_data_lo_2 ? _field_data_T_95 : _GEN_5344; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5346 = 14'h5c == field_data_lo_2 ? _field_data_T_96 : _GEN_5345; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5347 = 14'h5d == field_data_lo_2 ? _field_data_T_97 : _GEN_5346; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5348 = 14'h5e == field_data_lo_2 ? _field_data_T_98 : _GEN_5347; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5349 = 14'h5f == field_data_lo_2 ? _field_data_T_99 : _GEN_5348; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5350 = 14'h60 == field_data_lo_2 ? _field_data_T_100 : _GEN_5349; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5351 = 14'h61 == field_data_lo_2 ? _field_data_T_101 : _GEN_5350; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5352 = 14'h62 == field_data_lo_2 ? _field_data_T_102 : _GEN_5351; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5353 = 14'h63 == field_data_lo_2 ? _field_data_T_103 : _GEN_5352; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5354 = 14'h64 == field_data_lo_2 ? _field_data_T_104 : _GEN_5353; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5355 = 14'h65 == field_data_lo_2 ? _field_data_T_105 : _GEN_5354; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5356 = 14'h66 == field_data_lo_2 ? _field_data_T_106 : _GEN_5355; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5357 = 14'h67 == field_data_lo_2 ? _field_data_T_107 : _GEN_5356; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5358 = 14'h68 == field_data_lo_2 ? _field_data_T_108 : _GEN_5357; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5359 = 14'h69 == field_data_lo_2 ? _field_data_T_109 : _GEN_5358; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5360 = 14'h6a == field_data_lo_2 ? _field_data_T_110 : _GEN_5359; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5361 = 14'h6b == field_data_lo_2 ? _field_data_T_111 : _GEN_5360; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5362 = 14'h6c == field_data_lo_2 ? _field_data_T_112 : _GEN_5361; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5363 = 14'h6d == field_data_lo_2 ? _field_data_T_113 : _GEN_5362; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5364 = 14'h6e == field_data_lo_2 ? _field_data_T_114 : _GEN_5363; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5365 = 14'h6f == field_data_lo_2 ? _field_data_T_115 : _GEN_5364; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5366 = 14'h70 == field_data_lo_2 ? _field_data_T_116 : _GEN_5365; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5367 = 14'h71 == field_data_lo_2 ? _field_data_T_117 : _GEN_5366; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5368 = 14'h72 == field_data_lo_2 ? _field_data_T_118 : _GEN_5367; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5369 = 14'h73 == field_data_lo_2 ? _field_data_T_119 : _GEN_5368; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5370 = 14'h74 == field_data_lo_2 ? _field_data_T_120 : _GEN_5369; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5371 = 14'h75 == field_data_lo_2 ? _field_data_T_121 : _GEN_5370; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5372 = 14'h76 == field_data_lo_2 ? _field_data_T_122 : _GEN_5371; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5373 = 14'h77 == field_data_lo_2 ? _field_data_T_123 : _GEN_5372; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5374 = 14'h78 == field_data_lo_2 ? _field_data_T_124 : _GEN_5373; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5375 = 14'h79 == field_data_lo_2 ? _field_data_T_125 : _GEN_5374; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5376 = 14'h7a == field_data_lo_2 ? _field_data_T_126 : _GEN_5375; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5377 = 14'h7b == field_data_lo_2 ? _field_data_T_127 : _GEN_5376; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5378 = 14'h7c == field_data_lo_2 ? _field_data_T_128 : _GEN_5377; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5379 = 14'h7d == field_data_lo_2 ? _field_data_T_129 : _GEN_5378; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5380 = 14'h7e == field_data_lo_2 ? _field_data_T_130 : _GEN_5379; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5381 = 14'h7f == field_data_lo_2 ? _field_data_T_131 : _GEN_5380; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5382 = 14'h80 == field_data_lo_2 ? _field_data_T_132 : _GEN_5381; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5383 = 14'h81 == field_data_lo_2 ? _field_data_T_133 : _GEN_5382; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5384 = 14'h82 == field_data_lo_2 ? _field_data_T_134 : _GEN_5383; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5385 = 14'h83 == field_data_lo_2 ? _field_data_T_135 : _GEN_5384; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5386 = 14'h84 == field_data_lo_2 ? _field_data_T_136 : _GEN_5385; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5387 = 14'h85 == field_data_lo_2 ? _field_data_T_137 : _GEN_5386; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5388 = 14'h86 == field_data_lo_2 ? _field_data_T_138 : _GEN_5387; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5389 = 14'h87 == field_data_lo_2 ? _field_data_T_139 : _GEN_5388; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5390 = 14'h88 == field_data_lo_2 ? _field_data_T_140 : _GEN_5389; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5391 = 14'h89 == field_data_lo_2 ? _field_data_T_141 : _GEN_5390; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5392 = 14'h8a == field_data_lo_2 ? _field_data_T_142 : _GEN_5391; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5393 = 14'h8b == field_data_lo_2 ? _field_data_T_143 : _GEN_5392; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5394 = 14'h8c == field_data_lo_2 ? _field_data_T_144 : _GEN_5393; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5395 = 14'h8d == field_data_lo_2 ? _field_data_T_145 : _GEN_5394; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5396 = 14'h8e == field_data_lo_2 ? _field_data_T_146 : _GEN_5395; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5397 = 14'h8f == field_data_lo_2 ? _field_data_T_147 : _GEN_5396; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5398 = 14'h90 == field_data_lo_2 ? _field_data_T_148 : _GEN_5397; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5399 = 14'h91 == field_data_lo_2 ? _field_data_T_149 : _GEN_5398; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5400 = 14'h92 == field_data_lo_2 ? _field_data_T_150 : _GEN_5399; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5401 = 14'h93 == field_data_lo_2 ? _field_data_T_151 : _GEN_5400; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5402 = 14'h94 == field_data_lo_2 ? _field_data_T_152 : _GEN_5401; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5403 = 14'h95 == field_data_lo_2 ? _field_data_T_153 : _GEN_5402; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5404 = 14'h96 == field_data_lo_2 ? _field_data_T_154 : _GEN_5403; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5405 = 14'h97 == field_data_lo_2 ? _field_data_T_155 : _GEN_5404; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5406 = 14'h98 == field_data_lo_2 ? _field_data_T_156 : _GEN_5405; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5407 = 14'h99 == field_data_lo_2 ? _field_data_T_157 : _GEN_5406; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5408 = 14'h9a == field_data_lo_2 ? _field_data_T_158 : _GEN_5407; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5409 = 14'h9b == field_data_lo_2 ? _field_data_T_159 : _GEN_5408; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5410 = 14'h9c == field_data_lo_2 ? _field_data_T_160 : _GEN_5409; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5411 = 14'h9d == field_data_lo_2 ? _field_data_T_161 : _GEN_5410; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5412 = 14'h9e == field_data_lo_2 ? _field_data_T_162 : _GEN_5411; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5413 = 14'h9f == field_data_lo_2 ? _field_data_T_163 : _GEN_5412; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_67 = vliw_67[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_3 = vliw_67[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_67 = field_data_lo_3[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_67 = field_data_lo_3[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_70 = {{1'd0}, args_offset_67}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_70 = _total_offset_T_70[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_5417 = 3'h1 == total_offset_70 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5418 = 3'h2 == total_offset_70 ? args_2 : _GEN_5417; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5419 = 3'h3 == total_offset_70 ? args_3 : _GEN_5418; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5420 = 3'h4 == total_offset_70 ? args_4 : _GEN_5419; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5421 = 3'h5 == total_offset_70 ? args_5 : _GEN_5420; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5422 = 3'h6 == total_offset_70 ? args_6 : _GEN_5421; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5423 = total_offset_70 < 3'h7 ? _GEN_5422 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_67_1 = 3'h0 < args_length_67 ? _GEN_5423 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_71 = args_offset_67 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_5426 = 3'h1 == total_offset_71 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5427 = 3'h2 == total_offset_71 ? args_2 : _GEN_5426; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5428 = 3'h3 == total_offset_71 ? args_3 : _GEN_5427; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5429 = 3'h4 == total_offset_71 ? args_4 : _GEN_5428; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5430 = 3'h5 == total_offset_71 ? args_5 : _GEN_5429; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5431 = 3'h6 == total_offset_71 ? args_6 : _GEN_5430; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5432 = total_offset_71 < 3'h7 ? _GEN_5431 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_67_0 = 3'h1 < args_length_67 ? _GEN_5432 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_364 = {field_bytes_67_0,field_bytes_67_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5434 = opcode_67 == 4'ha ? _field_data_T_364 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_5435 = opcode_67 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_4864 = opcode_67 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_3 = field_data_lo_3[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_367 = {field_data_hi_3,field_data_lo_3}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_135 = _T_4864 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_5436 = opcode_67 == 4'h8 | opcode_67 == 4'hb ? _field_data_T_367 : _GEN_5434; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_5437 = opcode_67 == 4'h8 | opcode_67 == 4'hb ? _field_tag_T_135 : _GEN_5435; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_5438 = 14'h40 == field_data_lo_3 ? _field_data_T_68 : _GEN_5436; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5439 = 14'h41 == field_data_lo_3 ? _field_data_T_69 : _GEN_5438; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5440 = 14'h42 == field_data_lo_3 ? _field_data_T_70 : _GEN_5439; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5441 = 14'h43 == field_data_lo_3 ? _field_data_T_71 : _GEN_5440; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5442 = 14'h44 == field_data_lo_3 ? _field_data_T_72 : _GEN_5441; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5443 = 14'h45 == field_data_lo_3 ? _field_data_T_73 : _GEN_5442; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5444 = 14'h46 == field_data_lo_3 ? _field_data_T_74 : _GEN_5443; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5445 = 14'h47 == field_data_lo_3 ? _field_data_T_75 : _GEN_5444; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5446 = 14'h48 == field_data_lo_3 ? _field_data_T_76 : _GEN_5445; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5447 = 14'h49 == field_data_lo_3 ? _field_data_T_77 : _GEN_5446; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5448 = 14'h4a == field_data_lo_3 ? _field_data_T_78 : _GEN_5447; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5449 = 14'h4b == field_data_lo_3 ? _field_data_T_79 : _GEN_5448; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5450 = 14'h4c == field_data_lo_3 ? _field_data_T_80 : _GEN_5449; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5451 = 14'h4d == field_data_lo_3 ? _field_data_T_81 : _GEN_5450; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5452 = 14'h4e == field_data_lo_3 ? _field_data_T_82 : _GEN_5451; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5453 = 14'h4f == field_data_lo_3 ? _field_data_T_83 : _GEN_5452; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5454 = 14'h50 == field_data_lo_3 ? _field_data_T_84 : _GEN_5453; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5455 = 14'h51 == field_data_lo_3 ? _field_data_T_85 : _GEN_5454; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5456 = 14'h52 == field_data_lo_3 ? _field_data_T_86 : _GEN_5455; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5457 = 14'h53 == field_data_lo_3 ? _field_data_T_87 : _GEN_5456; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5458 = 14'h54 == field_data_lo_3 ? _field_data_T_88 : _GEN_5457; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5459 = 14'h55 == field_data_lo_3 ? _field_data_T_89 : _GEN_5458; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5460 = 14'h56 == field_data_lo_3 ? _field_data_T_90 : _GEN_5459; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5461 = 14'h57 == field_data_lo_3 ? _field_data_T_91 : _GEN_5460; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5462 = 14'h58 == field_data_lo_3 ? _field_data_T_92 : _GEN_5461; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5463 = 14'h59 == field_data_lo_3 ? _field_data_T_93 : _GEN_5462; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5464 = 14'h5a == field_data_lo_3 ? _field_data_T_94 : _GEN_5463; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5465 = 14'h5b == field_data_lo_3 ? _field_data_T_95 : _GEN_5464; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5466 = 14'h5c == field_data_lo_3 ? _field_data_T_96 : _GEN_5465; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5467 = 14'h5d == field_data_lo_3 ? _field_data_T_97 : _GEN_5466; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5468 = 14'h5e == field_data_lo_3 ? _field_data_T_98 : _GEN_5467; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5469 = 14'h5f == field_data_lo_3 ? _field_data_T_99 : _GEN_5468; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5470 = 14'h60 == field_data_lo_3 ? _field_data_T_100 : _GEN_5469; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5471 = 14'h61 == field_data_lo_3 ? _field_data_T_101 : _GEN_5470; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5472 = 14'h62 == field_data_lo_3 ? _field_data_T_102 : _GEN_5471; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5473 = 14'h63 == field_data_lo_3 ? _field_data_T_103 : _GEN_5472; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5474 = 14'h64 == field_data_lo_3 ? _field_data_T_104 : _GEN_5473; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5475 = 14'h65 == field_data_lo_3 ? _field_data_T_105 : _GEN_5474; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5476 = 14'h66 == field_data_lo_3 ? _field_data_T_106 : _GEN_5475; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5477 = 14'h67 == field_data_lo_3 ? _field_data_T_107 : _GEN_5476; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5478 = 14'h68 == field_data_lo_3 ? _field_data_T_108 : _GEN_5477; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5479 = 14'h69 == field_data_lo_3 ? _field_data_T_109 : _GEN_5478; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5480 = 14'h6a == field_data_lo_3 ? _field_data_T_110 : _GEN_5479; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5481 = 14'h6b == field_data_lo_3 ? _field_data_T_111 : _GEN_5480; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5482 = 14'h6c == field_data_lo_3 ? _field_data_T_112 : _GEN_5481; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5483 = 14'h6d == field_data_lo_3 ? _field_data_T_113 : _GEN_5482; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5484 = 14'h6e == field_data_lo_3 ? _field_data_T_114 : _GEN_5483; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5485 = 14'h6f == field_data_lo_3 ? _field_data_T_115 : _GEN_5484; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5486 = 14'h70 == field_data_lo_3 ? _field_data_T_116 : _GEN_5485; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5487 = 14'h71 == field_data_lo_3 ? _field_data_T_117 : _GEN_5486; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5488 = 14'h72 == field_data_lo_3 ? _field_data_T_118 : _GEN_5487; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5489 = 14'h73 == field_data_lo_3 ? _field_data_T_119 : _GEN_5488; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5490 = 14'h74 == field_data_lo_3 ? _field_data_T_120 : _GEN_5489; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5491 = 14'h75 == field_data_lo_3 ? _field_data_T_121 : _GEN_5490; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5492 = 14'h76 == field_data_lo_3 ? _field_data_T_122 : _GEN_5491; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5493 = 14'h77 == field_data_lo_3 ? _field_data_T_123 : _GEN_5492; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5494 = 14'h78 == field_data_lo_3 ? _field_data_T_124 : _GEN_5493; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5495 = 14'h79 == field_data_lo_3 ? _field_data_T_125 : _GEN_5494; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5496 = 14'h7a == field_data_lo_3 ? _field_data_T_126 : _GEN_5495; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5497 = 14'h7b == field_data_lo_3 ? _field_data_T_127 : _GEN_5496; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5498 = 14'h7c == field_data_lo_3 ? _field_data_T_128 : _GEN_5497; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5499 = 14'h7d == field_data_lo_3 ? _field_data_T_129 : _GEN_5498; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5500 = 14'h7e == field_data_lo_3 ? _field_data_T_130 : _GEN_5499; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5501 = 14'h7f == field_data_lo_3 ? _field_data_T_131 : _GEN_5500; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5502 = 14'h80 == field_data_lo_3 ? _field_data_T_132 : _GEN_5501; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5503 = 14'h81 == field_data_lo_3 ? _field_data_T_133 : _GEN_5502; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5504 = 14'h82 == field_data_lo_3 ? _field_data_T_134 : _GEN_5503; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5505 = 14'h83 == field_data_lo_3 ? _field_data_T_135 : _GEN_5504; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5506 = 14'h84 == field_data_lo_3 ? _field_data_T_136 : _GEN_5505; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5507 = 14'h85 == field_data_lo_3 ? _field_data_T_137 : _GEN_5506; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5508 = 14'h86 == field_data_lo_3 ? _field_data_T_138 : _GEN_5507; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5509 = 14'h87 == field_data_lo_3 ? _field_data_T_139 : _GEN_5508; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5510 = 14'h88 == field_data_lo_3 ? _field_data_T_140 : _GEN_5509; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5511 = 14'h89 == field_data_lo_3 ? _field_data_T_141 : _GEN_5510; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5512 = 14'h8a == field_data_lo_3 ? _field_data_T_142 : _GEN_5511; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5513 = 14'h8b == field_data_lo_3 ? _field_data_T_143 : _GEN_5512; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5514 = 14'h8c == field_data_lo_3 ? _field_data_T_144 : _GEN_5513; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5515 = 14'h8d == field_data_lo_3 ? _field_data_T_145 : _GEN_5514; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5516 = 14'h8e == field_data_lo_3 ? _field_data_T_146 : _GEN_5515; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5517 = 14'h8f == field_data_lo_3 ? _field_data_T_147 : _GEN_5516; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5518 = 14'h90 == field_data_lo_3 ? _field_data_T_148 : _GEN_5517; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5519 = 14'h91 == field_data_lo_3 ? _field_data_T_149 : _GEN_5518; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5520 = 14'h92 == field_data_lo_3 ? _field_data_T_150 : _GEN_5519; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5521 = 14'h93 == field_data_lo_3 ? _field_data_T_151 : _GEN_5520; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5522 = 14'h94 == field_data_lo_3 ? _field_data_T_152 : _GEN_5521; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5523 = 14'h95 == field_data_lo_3 ? _field_data_T_153 : _GEN_5522; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5524 = 14'h96 == field_data_lo_3 ? _field_data_T_154 : _GEN_5523; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5525 = 14'h97 == field_data_lo_3 ? _field_data_T_155 : _GEN_5524; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5526 = 14'h98 == field_data_lo_3 ? _field_data_T_156 : _GEN_5525; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5527 = 14'h99 == field_data_lo_3 ? _field_data_T_157 : _GEN_5526; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5528 = 14'h9a == field_data_lo_3 ? _field_data_T_158 : _GEN_5527; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5529 = 14'h9b == field_data_lo_3 ? _field_data_T_159 : _GEN_5528; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5530 = 14'h9c == field_data_lo_3 ? _field_data_T_160 : _GEN_5529; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5531 = 14'h9d == field_data_lo_3 ? _field_data_T_161 : _GEN_5530; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5532 = 14'h9e == field_data_lo_3 ? _field_data_T_162 : _GEN_5531; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5533 = 14'h9f == field_data_lo_3 ? _field_data_T_163 : _GEN_5532; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_68 = vliw_68[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_4 = vliw_68[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_68 = field_data_lo_4[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_68 = field_data_lo_4[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_72 = {{1'd0}, args_offset_68}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_72 = _total_offset_T_72[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_5537 = 3'h1 == total_offset_72 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5538 = 3'h2 == total_offset_72 ? args_2 : _GEN_5537; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5539 = 3'h3 == total_offset_72 ? args_3 : _GEN_5538; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5540 = 3'h4 == total_offset_72 ? args_4 : _GEN_5539; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5541 = 3'h5 == total_offset_72 ? args_5 : _GEN_5540; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5542 = 3'h6 == total_offset_72 ? args_6 : _GEN_5541; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5543 = total_offset_72 < 3'h7 ? _GEN_5542 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_68_1 = 3'h0 < args_length_68 ? _GEN_5543 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_73 = args_offset_68 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_5546 = 3'h1 == total_offset_73 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5547 = 3'h2 == total_offset_73 ? args_2 : _GEN_5546; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5548 = 3'h3 == total_offset_73 ? args_3 : _GEN_5547; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5549 = 3'h4 == total_offset_73 ? args_4 : _GEN_5548; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5550 = 3'h5 == total_offset_73 ? args_5 : _GEN_5549; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5551 = 3'h6 == total_offset_73 ? args_6 : _GEN_5550; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5552 = total_offset_73 < 3'h7 ? _GEN_5551 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_68_0 = 3'h1 < args_length_68 ? _GEN_5552 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_464 = {field_bytes_68_0,field_bytes_68_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5554 = opcode_68 == 4'ha ? _field_data_T_464 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_5555 = opcode_68 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_4969 = opcode_68 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_4 = field_data_lo_4[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_467 = {field_data_hi_4,field_data_lo_4}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_137 = _T_4969 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_5556 = opcode_68 == 4'h8 | opcode_68 == 4'hb ? _field_data_T_467 : _GEN_5554; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_5557 = opcode_68 == 4'h8 | opcode_68 == 4'hb ? _field_tag_T_137 : _GEN_5555; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_5558 = 14'h40 == field_data_lo_4 ? _field_data_T_68 : _GEN_5556; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5559 = 14'h41 == field_data_lo_4 ? _field_data_T_69 : _GEN_5558; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5560 = 14'h42 == field_data_lo_4 ? _field_data_T_70 : _GEN_5559; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5561 = 14'h43 == field_data_lo_4 ? _field_data_T_71 : _GEN_5560; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5562 = 14'h44 == field_data_lo_4 ? _field_data_T_72 : _GEN_5561; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5563 = 14'h45 == field_data_lo_4 ? _field_data_T_73 : _GEN_5562; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5564 = 14'h46 == field_data_lo_4 ? _field_data_T_74 : _GEN_5563; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5565 = 14'h47 == field_data_lo_4 ? _field_data_T_75 : _GEN_5564; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5566 = 14'h48 == field_data_lo_4 ? _field_data_T_76 : _GEN_5565; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5567 = 14'h49 == field_data_lo_4 ? _field_data_T_77 : _GEN_5566; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5568 = 14'h4a == field_data_lo_4 ? _field_data_T_78 : _GEN_5567; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5569 = 14'h4b == field_data_lo_4 ? _field_data_T_79 : _GEN_5568; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5570 = 14'h4c == field_data_lo_4 ? _field_data_T_80 : _GEN_5569; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5571 = 14'h4d == field_data_lo_4 ? _field_data_T_81 : _GEN_5570; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5572 = 14'h4e == field_data_lo_4 ? _field_data_T_82 : _GEN_5571; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5573 = 14'h4f == field_data_lo_4 ? _field_data_T_83 : _GEN_5572; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5574 = 14'h50 == field_data_lo_4 ? _field_data_T_84 : _GEN_5573; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5575 = 14'h51 == field_data_lo_4 ? _field_data_T_85 : _GEN_5574; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5576 = 14'h52 == field_data_lo_4 ? _field_data_T_86 : _GEN_5575; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5577 = 14'h53 == field_data_lo_4 ? _field_data_T_87 : _GEN_5576; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5578 = 14'h54 == field_data_lo_4 ? _field_data_T_88 : _GEN_5577; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5579 = 14'h55 == field_data_lo_4 ? _field_data_T_89 : _GEN_5578; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5580 = 14'h56 == field_data_lo_4 ? _field_data_T_90 : _GEN_5579; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5581 = 14'h57 == field_data_lo_4 ? _field_data_T_91 : _GEN_5580; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5582 = 14'h58 == field_data_lo_4 ? _field_data_T_92 : _GEN_5581; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5583 = 14'h59 == field_data_lo_4 ? _field_data_T_93 : _GEN_5582; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5584 = 14'h5a == field_data_lo_4 ? _field_data_T_94 : _GEN_5583; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5585 = 14'h5b == field_data_lo_4 ? _field_data_T_95 : _GEN_5584; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5586 = 14'h5c == field_data_lo_4 ? _field_data_T_96 : _GEN_5585; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5587 = 14'h5d == field_data_lo_4 ? _field_data_T_97 : _GEN_5586; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5588 = 14'h5e == field_data_lo_4 ? _field_data_T_98 : _GEN_5587; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5589 = 14'h5f == field_data_lo_4 ? _field_data_T_99 : _GEN_5588; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5590 = 14'h60 == field_data_lo_4 ? _field_data_T_100 : _GEN_5589; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5591 = 14'h61 == field_data_lo_4 ? _field_data_T_101 : _GEN_5590; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5592 = 14'h62 == field_data_lo_4 ? _field_data_T_102 : _GEN_5591; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5593 = 14'h63 == field_data_lo_4 ? _field_data_T_103 : _GEN_5592; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5594 = 14'h64 == field_data_lo_4 ? _field_data_T_104 : _GEN_5593; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5595 = 14'h65 == field_data_lo_4 ? _field_data_T_105 : _GEN_5594; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5596 = 14'h66 == field_data_lo_4 ? _field_data_T_106 : _GEN_5595; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5597 = 14'h67 == field_data_lo_4 ? _field_data_T_107 : _GEN_5596; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5598 = 14'h68 == field_data_lo_4 ? _field_data_T_108 : _GEN_5597; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5599 = 14'h69 == field_data_lo_4 ? _field_data_T_109 : _GEN_5598; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5600 = 14'h6a == field_data_lo_4 ? _field_data_T_110 : _GEN_5599; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5601 = 14'h6b == field_data_lo_4 ? _field_data_T_111 : _GEN_5600; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5602 = 14'h6c == field_data_lo_4 ? _field_data_T_112 : _GEN_5601; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5603 = 14'h6d == field_data_lo_4 ? _field_data_T_113 : _GEN_5602; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5604 = 14'h6e == field_data_lo_4 ? _field_data_T_114 : _GEN_5603; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5605 = 14'h6f == field_data_lo_4 ? _field_data_T_115 : _GEN_5604; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5606 = 14'h70 == field_data_lo_4 ? _field_data_T_116 : _GEN_5605; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5607 = 14'h71 == field_data_lo_4 ? _field_data_T_117 : _GEN_5606; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5608 = 14'h72 == field_data_lo_4 ? _field_data_T_118 : _GEN_5607; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5609 = 14'h73 == field_data_lo_4 ? _field_data_T_119 : _GEN_5608; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5610 = 14'h74 == field_data_lo_4 ? _field_data_T_120 : _GEN_5609; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5611 = 14'h75 == field_data_lo_4 ? _field_data_T_121 : _GEN_5610; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5612 = 14'h76 == field_data_lo_4 ? _field_data_T_122 : _GEN_5611; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5613 = 14'h77 == field_data_lo_4 ? _field_data_T_123 : _GEN_5612; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5614 = 14'h78 == field_data_lo_4 ? _field_data_T_124 : _GEN_5613; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5615 = 14'h79 == field_data_lo_4 ? _field_data_T_125 : _GEN_5614; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5616 = 14'h7a == field_data_lo_4 ? _field_data_T_126 : _GEN_5615; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5617 = 14'h7b == field_data_lo_4 ? _field_data_T_127 : _GEN_5616; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5618 = 14'h7c == field_data_lo_4 ? _field_data_T_128 : _GEN_5617; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5619 = 14'h7d == field_data_lo_4 ? _field_data_T_129 : _GEN_5618; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5620 = 14'h7e == field_data_lo_4 ? _field_data_T_130 : _GEN_5619; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5621 = 14'h7f == field_data_lo_4 ? _field_data_T_131 : _GEN_5620; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5622 = 14'h80 == field_data_lo_4 ? _field_data_T_132 : _GEN_5621; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5623 = 14'h81 == field_data_lo_4 ? _field_data_T_133 : _GEN_5622; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5624 = 14'h82 == field_data_lo_4 ? _field_data_T_134 : _GEN_5623; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5625 = 14'h83 == field_data_lo_4 ? _field_data_T_135 : _GEN_5624; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5626 = 14'h84 == field_data_lo_4 ? _field_data_T_136 : _GEN_5625; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5627 = 14'h85 == field_data_lo_4 ? _field_data_T_137 : _GEN_5626; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5628 = 14'h86 == field_data_lo_4 ? _field_data_T_138 : _GEN_5627; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5629 = 14'h87 == field_data_lo_4 ? _field_data_T_139 : _GEN_5628; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5630 = 14'h88 == field_data_lo_4 ? _field_data_T_140 : _GEN_5629; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5631 = 14'h89 == field_data_lo_4 ? _field_data_T_141 : _GEN_5630; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5632 = 14'h8a == field_data_lo_4 ? _field_data_T_142 : _GEN_5631; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5633 = 14'h8b == field_data_lo_4 ? _field_data_T_143 : _GEN_5632; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5634 = 14'h8c == field_data_lo_4 ? _field_data_T_144 : _GEN_5633; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5635 = 14'h8d == field_data_lo_4 ? _field_data_T_145 : _GEN_5634; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5636 = 14'h8e == field_data_lo_4 ? _field_data_T_146 : _GEN_5635; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5637 = 14'h8f == field_data_lo_4 ? _field_data_T_147 : _GEN_5636; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5638 = 14'h90 == field_data_lo_4 ? _field_data_T_148 : _GEN_5637; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5639 = 14'h91 == field_data_lo_4 ? _field_data_T_149 : _GEN_5638; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5640 = 14'h92 == field_data_lo_4 ? _field_data_T_150 : _GEN_5639; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5641 = 14'h93 == field_data_lo_4 ? _field_data_T_151 : _GEN_5640; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5642 = 14'h94 == field_data_lo_4 ? _field_data_T_152 : _GEN_5641; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5643 = 14'h95 == field_data_lo_4 ? _field_data_T_153 : _GEN_5642; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5644 = 14'h96 == field_data_lo_4 ? _field_data_T_154 : _GEN_5643; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5645 = 14'h97 == field_data_lo_4 ? _field_data_T_155 : _GEN_5644; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5646 = 14'h98 == field_data_lo_4 ? _field_data_T_156 : _GEN_5645; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5647 = 14'h99 == field_data_lo_4 ? _field_data_T_157 : _GEN_5646; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5648 = 14'h9a == field_data_lo_4 ? _field_data_T_158 : _GEN_5647; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5649 = 14'h9b == field_data_lo_4 ? _field_data_T_159 : _GEN_5648; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5650 = 14'h9c == field_data_lo_4 ? _field_data_T_160 : _GEN_5649; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5651 = 14'h9d == field_data_lo_4 ? _field_data_T_161 : _GEN_5650; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5652 = 14'h9e == field_data_lo_4 ? _field_data_T_162 : _GEN_5651; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5653 = 14'h9f == field_data_lo_4 ? _field_data_T_163 : _GEN_5652; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_69 = vliw_69[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_5 = vliw_69[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_69 = field_data_lo_5[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_69 = field_data_lo_5[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_74 = {{1'd0}, args_offset_69}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_74 = _total_offset_T_74[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_5657 = 3'h1 == total_offset_74 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5658 = 3'h2 == total_offset_74 ? args_2 : _GEN_5657; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5659 = 3'h3 == total_offset_74 ? args_3 : _GEN_5658; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5660 = 3'h4 == total_offset_74 ? args_4 : _GEN_5659; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5661 = 3'h5 == total_offset_74 ? args_5 : _GEN_5660; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5662 = 3'h6 == total_offset_74 ? args_6 : _GEN_5661; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5663 = total_offset_74 < 3'h7 ? _GEN_5662 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_69_1 = 3'h0 < args_length_69 ? _GEN_5663 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_75 = args_offset_69 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_5666 = 3'h1 == total_offset_75 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5667 = 3'h2 == total_offset_75 ? args_2 : _GEN_5666; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5668 = 3'h3 == total_offset_75 ? args_3 : _GEN_5667; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5669 = 3'h4 == total_offset_75 ? args_4 : _GEN_5668; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5670 = 3'h5 == total_offset_75 ? args_5 : _GEN_5669; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5671 = 3'h6 == total_offset_75 ? args_6 : _GEN_5670; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5672 = total_offset_75 < 3'h7 ? _GEN_5671 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_69_0 = 3'h1 < args_length_69 ? _GEN_5672 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_564 = {field_bytes_69_0,field_bytes_69_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_5674 = opcode_69 == 4'ha ? _field_data_T_564 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_5675 = opcode_69 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_5074 = opcode_69 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_5 = field_data_lo_5[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_567 = {field_data_hi_5,field_data_lo_5}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_139 = _T_5074 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_5676 = opcode_69 == 4'h8 | opcode_69 == 4'hb ? _field_data_T_567 : _GEN_5674; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_5677 = opcode_69 == 4'h8 | opcode_69 == 4'hb ? _field_tag_T_139 : _GEN_5675; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_5678 = 14'h40 == field_data_lo_5 ? _field_data_T_68 : _GEN_5676; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5679 = 14'h41 == field_data_lo_5 ? _field_data_T_69 : _GEN_5678; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5680 = 14'h42 == field_data_lo_5 ? _field_data_T_70 : _GEN_5679; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5681 = 14'h43 == field_data_lo_5 ? _field_data_T_71 : _GEN_5680; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5682 = 14'h44 == field_data_lo_5 ? _field_data_T_72 : _GEN_5681; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5683 = 14'h45 == field_data_lo_5 ? _field_data_T_73 : _GEN_5682; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5684 = 14'h46 == field_data_lo_5 ? _field_data_T_74 : _GEN_5683; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5685 = 14'h47 == field_data_lo_5 ? _field_data_T_75 : _GEN_5684; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5686 = 14'h48 == field_data_lo_5 ? _field_data_T_76 : _GEN_5685; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5687 = 14'h49 == field_data_lo_5 ? _field_data_T_77 : _GEN_5686; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5688 = 14'h4a == field_data_lo_5 ? _field_data_T_78 : _GEN_5687; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5689 = 14'h4b == field_data_lo_5 ? _field_data_T_79 : _GEN_5688; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5690 = 14'h4c == field_data_lo_5 ? _field_data_T_80 : _GEN_5689; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5691 = 14'h4d == field_data_lo_5 ? _field_data_T_81 : _GEN_5690; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5692 = 14'h4e == field_data_lo_5 ? _field_data_T_82 : _GEN_5691; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5693 = 14'h4f == field_data_lo_5 ? _field_data_T_83 : _GEN_5692; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5694 = 14'h50 == field_data_lo_5 ? _field_data_T_84 : _GEN_5693; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5695 = 14'h51 == field_data_lo_5 ? _field_data_T_85 : _GEN_5694; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5696 = 14'h52 == field_data_lo_5 ? _field_data_T_86 : _GEN_5695; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5697 = 14'h53 == field_data_lo_5 ? _field_data_T_87 : _GEN_5696; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5698 = 14'h54 == field_data_lo_5 ? _field_data_T_88 : _GEN_5697; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5699 = 14'h55 == field_data_lo_5 ? _field_data_T_89 : _GEN_5698; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5700 = 14'h56 == field_data_lo_5 ? _field_data_T_90 : _GEN_5699; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5701 = 14'h57 == field_data_lo_5 ? _field_data_T_91 : _GEN_5700; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5702 = 14'h58 == field_data_lo_5 ? _field_data_T_92 : _GEN_5701; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5703 = 14'h59 == field_data_lo_5 ? _field_data_T_93 : _GEN_5702; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5704 = 14'h5a == field_data_lo_5 ? _field_data_T_94 : _GEN_5703; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5705 = 14'h5b == field_data_lo_5 ? _field_data_T_95 : _GEN_5704; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5706 = 14'h5c == field_data_lo_5 ? _field_data_T_96 : _GEN_5705; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5707 = 14'h5d == field_data_lo_5 ? _field_data_T_97 : _GEN_5706; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5708 = 14'h5e == field_data_lo_5 ? _field_data_T_98 : _GEN_5707; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5709 = 14'h5f == field_data_lo_5 ? _field_data_T_99 : _GEN_5708; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5710 = 14'h60 == field_data_lo_5 ? _field_data_T_100 : _GEN_5709; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5711 = 14'h61 == field_data_lo_5 ? _field_data_T_101 : _GEN_5710; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5712 = 14'h62 == field_data_lo_5 ? _field_data_T_102 : _GEN_5711; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5713 = 14'h63 == field_data_lo_5 ? _field_data_T_103 : _GEN_5712; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5714 = 14'h64 == field_data_lo_5 ? _field_data_T_104 : _GEN_5713; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5715 = 14'h65 == field_data_lo_5 ? _field_data_T_105 : _GEN_5714; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5716 = 14'h66 == field_data_lo_5 ? _field_data_T_106 : _GEN_5715; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5717 = 14'h67 == field_data_lo_5 ? _field_data_T_107 : _GEN_5716; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5718 = 14'h68 == field_data_lo_5 ? _field_data_T_108 : _GEN_5717; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5719 = 14'h69 == field_data_lo_5 ? _field_data_T_109 : _GEN_5718; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5720 = 14'h6a == field_data_lo_5 ? _field_data_T_110 : _GEN_5719; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5721 = 14'h6b == field_data_lo_5 ? _field_data_T_111 : _GEN_5720; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5722 = 14'h6c == field_data_lo_5 ? _field_data_T_112 : _GEN_5721; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5723 = 14'h6d == field_data_lo_5 ? _field_data_T_113 : _GEN_5722; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5724 = 14'h6e == field_data_lo_5 ? _field_data_T_114 : _GEN_5723; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5725 = 14'h6f == field_data_lo_5 ? _field_data_T_115 : _GEN_5724; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5726 = 14'h70 == field_data_lo_5 ? _field_data_T_116 : _GEN_5725; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5727 = 14'h71 == field_data_lo_5 ? _field_data_T_117 : _GEN_5726; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5728 = 14'h72 == field_data_lo_5 ? _field_data_T_118 : _GEN_5727; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5729 = 14'h73 == field_data_lo_5 ? _field_data_T_119 : _GEN_5728; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5730 = 14'h74 == field_data_lo_5 ? _field_data_T_120 : _GEN_5729; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5731 = 14'h75 == field_data_lo_5 ? _field_data_T_121 : _GEN_5730; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5732 = 14'h76 == field_data_lo_5 ? _field_data_T_122 : _GEN_5731; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5733 = 14'h77 == field_data_lo_5 ? _field_data_T_123 : _GEN_5732; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5734 = 14'h78 == field_data_lo_5 ? _field_data_T_124 : _GEN_5733; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5735 = 14'h79 == field_data_lo_5 ? _field_data_T_125 : _GEN_5734; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5736 = 14'h7a == field_data_lo_5 ? _field_data_T_126 : _GEN_5735; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5737 = 14'h7b == field_data_lo_5 ? _field_data_T_127 : _GEN_5736; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5738 = 14'h7c == field_data_lo_5 ? _field_data_T_128 : _GEN_5737; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5739 = 14'h7d == field_data_lo_5 ? _field_data_T_129 : _GEN_5738; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5740 = 14'h7e == field_data_lo_5 ? _field_data_T_130 : _GEN_5739; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5741 = 14'h7f == field_data_lo_5 ? _field_data_T_131 : _GEN_5740; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5742 = 14'h80 == field_data_lo_5 ? _field_data_T_132 : _GEN_5741; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5743 = 14'h81 == field_data_lo_5 ? _field_data_T_133 : _GEN_5742; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5744 = 14'h82 == field_data_lo_5 ? _field_data_T_134 : _GEN_5743; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5745 = 14'h83 == field_data_lo_5 ? _field_data_T_135 : _GEN_5744; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5746 = 14'h84 == field_data_lo_5 ? _field_data_T_136 : _GEN_5745; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5747 = 14'h85 == field_data_lo_5 ? _field_data_T_137 : _GEN_5746; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5748 = 14'h86 == field_data_lo_5 ? _field_data_T_138 : _GEN_5747; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5749 = 14'h87 == field_data_lo_5 ? _field_data_T_139 : _GEN_5748; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5750 = 14'h88 == field_data_lo_5 ? _field_data_T_140 : _GEN_5749; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5751 = 14'h89 == field_data_lo_5 ? _field_data_T_141 : _GEN_5750; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5752 = 14'h8a == field_data_lo_5 ? _field_data_T_142 : _GEN_5751; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5753 = 14'h8b == field_data_lo_5 ? _field_data_T_143 : _GEN_5752; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5754 = 14'h8c == field_data_lo_5 ? _field_data_T_144 : _GEN_5753; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5755 = 14'h8d == field_data_lo_5 ? _field_data_T_145 : _GEN_5754; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5756 = 14'h8e == field_data_lo_5 ? _field_data_T_146 : _GEN_5755; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5757 = 14'h8f == field_data_lo_5 ? _field_data_T_147 : _GEN_5756; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5758 = 14'h90 == field_data_lo_5 ? _field_data_T_148 : _GEN_5757; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5759 = 14'h91 == field_data_lo_5 ? _field_data_T_149 : _GEN_5758; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5760 = 14'h92 == field_data_lo_5 ? _field_data_T_150 : _GEN_5759; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5761 = 14'h93 == field_data_lo_5 ? _field_data_T_151 : _GEN_5760; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5762 = 14'h94 == field_data_lo_5 ? _field_data_T_152 : _GEN_5761; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5763 = 14'h95 == field_data_lo_5 ? _field_data_T_153 : _GEN_5762; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5764 = 14'h96 == field_data_lo_5 ? _field_data_T_154 : _GEN_5763; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5765 = 14'h97 == field_data_lo_5 ? _field_data_T_155 : _GEN_5764; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5766 = 14'h98 == field_data_lo_5 ? _field_data_T_156 : _GEN_5765; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5767 = 14'h99 == field_data_lo_5 ? _field_data_T_157 : _GEN_5766; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5768 = 14'h9a == field_data_lo_5 ? _field_data_T_158 : _GEN_5767; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5769 = 14'h9b == field_data_lo_5 ? _field_data_T_159 : _GEN_5768; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5770 = 14'h9c == field_data_lo_5 ? _field_data_T_160 : _GEN_5769; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5771 = 14'h9d == field_data_lo_5 ? _field_data_T_161 : _GEN_5770; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5772 = 14'h9e == field_data_lo_5 ? _field_data_T_162 : _GEN_5771; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_5773 = 14'h9f == field_data_lo_5 ? _field_data_T_163 : _GEN_5772; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_96 = phv_data_96; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_97 = phv_data_97; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_98 = phv_data_98; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_99 = phv_data_99; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_100 = phv_data_100; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_101 = phv_data_101; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_102 = phv_data_102; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_103 = phv_data_103; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_104 = phv_data_104; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_105 = phv_data_105; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_106 = phv_data_106; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_107 = phv_data_107; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_108 = phv_data_108; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_109 = phv_data_109; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_110 = phv_data_110; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_111 = phv_data_111; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_112 = phv_data_112; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_113 = phv_data_113; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_114 = phv_data_114; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_115 = phv_data_115; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_116 = phv_data_116; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_117 = phv_data_117; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_118 = phv_data_118; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_119 = phv_data_119; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_120 = phv_data_120; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_121 = phv_data_121; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_122 = phv_data_122; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_123 = phv_data_123; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_124 = phv_data_124; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_125 = phv_data_125; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_126 = phv_data_126; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_127 = phv_data_127; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_128 = phv_data_128; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_129 = phv_data_129; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_130 = phv_data_130; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_131 = phv_data_131; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_132 = phv_data_132; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_133 = phv_data_133; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_134 = phv_data_134; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_135 = phv_data_135; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_136 = phv_data_136; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_137 = phv_data_137; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_138 = phv_data_138; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_139 = phv_data_139; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_140 = phv_data_140; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_141 = phv_data_141; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_142 = phv_data_142; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_143 = phv_data_143; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_144 = phv_data_144; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_145 = phv_data_145; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_146 = phv_data_146; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_147 = phv_data_147; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_148 = phv_data_148; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_149 = phv_data_149; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_150 = phv_data_150; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_151 = phv_data_151; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_152 = phv_data_152; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_153 = phv_data_153; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_154 = phv_data_154; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_155 = phv_data_155; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_156 = phv_data_156; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_157 = phv_data_157; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_158 = phv_data_158; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_159 = phv_data_159; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_160 = phv_data_160; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_161 = phv_data_161; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_162 = phv_data_162; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_163 = phv_data_163; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_164 = phv_data_164; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_165 = phv_data_165; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_166 = phv_data_166; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_167 = phv_data_167; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_168 = phv_data_168; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_169 = phv_data_169; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_170 = phv_data_170; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_171 = phv_data_171; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_172 = phv_data_172; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_173 = phv_data_173; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_174 = phv_data_174; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_175 = phv_data_175; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_176 = phv_data_176; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_177 = phv_data_177; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_178 = phv_data_178; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_179 = phv_data_179; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_180 = phv_data_180; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_181 = phv_data_181; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_182 = phv_data_182; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_183 = phv_data_183; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_184 = phv_data_184; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_185 = phv_data_185; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_186 = phv_data_186; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_187 = phv_data_187; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_188 = phv_data_188; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_189 = phv_data_189; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_190 = phv_data_190; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_191 = phv_data_191; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_192 = phv_data_192; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_193 = phv_data_193; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_194 = phv_data_194; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_195 = phv_data_195; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_196 = phv_data_196; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_197 = phv_data_197; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_198 = phv_data_198; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_199 = phv_data_199; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_200 = phv_data_200; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_201 = phv_data_201; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_202 = phv_data_202; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_203 = phv_data_203; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_204 = phv_data_204; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_205 = phv_data_205; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_206 = phv_data_206; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_207 = phv_data_207; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_208 = phv_data_208; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_209 = phv_data_209; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_210 = phv_data_210; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_211 = phv_data_211; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_212 = phv_data_212; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_213 = phv_data_213; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_214 = phv_data_214; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_215 = phv_data_215; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_216 = phv_data_216; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_217 = phv_data_217; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_218 = phv_data_218; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_219 = phv_data_219; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_220 = phv_data_220; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_221 = phv_data_221; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_222 = phv_data_222; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_223 = phv_data_223; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_224 = phv_data_224; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_225 = phv_data_225; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_226 = phv_data_226; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_227 = phv_data_227; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_228 = phv_data_228; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_229 = phv_data_229; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_230 = phv_data_230; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_231 = phv_data_231; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_232 = phv_data_232; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_233 = phv_data_233; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_234 = phv_data_234; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_235 = phv_data_235; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_236 = phv_data_236; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_237 = phv_data_237; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_238 = phv_data_238; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_239 = phv_data_239; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_240 = phv_data_240; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_241 = phv_data_241; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_242 = phv_data_242; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_243 = phv_data_243; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_244 = phv_data_244; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_245 = phv_data_245; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_246 = phv_data_246; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_247 = phv_data_247; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_248 = phv_data_248; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_249 = phv_data_249; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_250 = phv_data_250; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_251 = phv_data_251; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_252 = phv_data_252; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_253 = phv_data_253; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_254 = phv_data_254; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_255 = phv_data_255; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_256 = phv_data_256; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_257 = phv_data_257; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_258 = phv_data_258; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_259 = phv_data_259; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_260 = phv_data_260; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_261 = phv_data_261; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_262 = phv_data_262; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_263 = phv_data_263; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_264 = phv_data_264; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_265 = phv_data_265; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_266 = phv_data_266; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_267 = phv_data_267; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_268 = phv_data_268; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_269 = phv_data_269; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_270 = phv_data_270; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_271 = phv_data_271; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_272 = phv_data_272; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_273 = phv_data_273; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_274 = phv_data_274; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_275 = phv_data_275; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_276 = phv_data_276; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_277 = phv_data_277; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_278 = phv_data_278; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_279 = phv_data_279; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_280 = phv_data_280; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_281 = phv_data_281; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_282 = phv_data_282; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_283 = phv_data_283; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_284 = phv_data_284; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_285 = phv_data_285; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_286 = phv_data_286; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_287 = phv_data_287; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_288 = phv_data_288; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_289 = phv_data_289; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_290 = phv_data_290; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_291 = phv_data_291; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_292 = phv_data_292; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_293 = phv_data_293; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_294 = phv_data_294; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_295 = phv_data_295; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_296 = phv_data_296; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_297 = phv_data_297; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_298 = phv_data_298; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_299 = phv_data_299; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_300 = phv_data_300; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_301 = phv_data_301; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_302 = phv_data_302; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_303 = phv_data_303; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_304 = phv_data_304; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_305 = phv_data_305; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_306 = phv_data_306; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_307 = phv_data_307; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_308 = phv_data_308; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_309 = phv_data_309; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_310 = phv_data_310; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_311 = phv_data_311; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_312 = phv_data_312; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_313 = phv_data_313; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_314 = phv_data_314; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_315 = phv_data_315; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_316 = phv_data_316; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_317 = phv_data_317; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_318 = phv_data_318; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_319 = phv_data_319; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_320 = phv_data_320; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_321 = phv_data_321; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_322 = phv_data_322; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_323 = phv_data_323; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_324 = phv_data_324; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_325 = phv_data_325; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_326 = phv_data_326; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_327 = phv_data_327; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_328 = phv_data_328; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_329 = phv_data_329; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_330 = phv_data_330; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_331 = phv_data_331; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_332 = phv_data_332; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_333 = phv_data_333; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_334 = phv_data_334; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_335 = phv_data_335; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_336 = phv_data_336; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_337 = phv_data_337; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_338 = phv_data_338; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_339 = phv_data_339; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_340 = phv_data_340; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_341 = phv_data_341; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_342 = phv_data_342; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_343 = phv_data_343; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_344 = phv_data_344; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_345 = phv_data_345; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_346 = phv_data_346; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_347 = phv_data_347; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_348 = phv_data_348; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_349 = phv_data_349; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_350 = phv_data_350; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_351 = phv_data_351; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_352 = phv_data_352; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_353 = phv_data_353; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_354 = phv_data_354; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_355 = phv_data_355; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_356 = phv_data_356; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_357 = phv_data_357; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_358 = phv_data_358; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_359 = phv_data_359; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_360 = phv_data_360; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_361 = phv_data_361; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_362 = phv_data_362; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_363 = phv_data_363; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_364 = phv_data_364; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_365 = phv_data_365; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_366 = phv_data_366; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_367 = phv_data_367; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_368 = phv_data_368; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_369 = phv_data_369; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_370 = phv_data_370; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_371 = phv_data_371; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_372 = phv_data_372; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_373 = phv_data_373; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_374 = phv_data_374; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_375 = phv_data_375; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_376 = phv_data_376; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_377 = phv_data_377; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_378 = phv_data_378; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_379 = phv_data_379; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_380 = phv_data_380; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_381 = phv_data_381; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_382 = phv_data_382; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_383 = phv_data_383; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_384 = phv_data_384; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_385 = phv_data_385; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_386 = phv_data_386; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_387 = phv_data_387; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_388 = phv_data_388; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_389 = phv_data_389; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_390 = phv_data_390; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_391 = phv_data_391; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_392 = phv_data_392; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_393 = phv_data_393; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_394 = phv_data_394; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_395 = phv_data_395; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_396 = phv_data_396; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_397 = phv_data_397; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_398 = phv_data_398; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_399 = phv_data_399; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_400 = phv_data_400; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_401 = phv_data_401; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_402 = phv_data_402; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_403 = phv_data_403; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_404 = phv_data_404; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_405 = phv_data_405; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_406 = phv_data_406; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_407 = phv_data_407; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_408 = phv_data_408; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_409 = phv_data_409; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_410 = phv_data_410; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_411 = phv_data_411; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_412 = phv_data_412; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_413 = phv_data_413; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_414 = phv_data_414; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_415 = phv_data_415; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_416 = phv_data_416; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_417 = phv_data_417; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_418 = phv_data_418; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_419 = phv_data_419; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_420 = phv_data_420; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_421 = phv_data_421; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_422 = phv_data_422; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_423 = phv_data_423; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_424 = phv_data_424; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_425 = phv_data_425; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_426 = phv_data_426; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_427 = phv_data_427; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_428 = phv_data_428; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_429 = phv_data_429; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_430 = phv_data_430; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_431 = phv_data_431; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_432 = phv_data_432; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_433 = phv_data_433; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_434 = phv_data_434; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_435 = phv_data_435; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_436 = phv_data_436; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_437 = phv_data_437; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_438 = phv_data_438; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_439 = phv_data_439; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_440 = phv_data_440; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_441 = phv_data_441; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_442 = phv_data_442; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_443 = phv_data_443; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_444 = phv_data_444; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_445 = phv_data_445; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_446 = phv_data_446; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_447 = phv_data_447; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_448 = phv_data_448; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_449 = phv_data_449; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_450 = phv_data_450; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_451 = phv_data_451; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_452 = phv_data_452; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_453 = phv_data_453; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_454 = phv_data_454; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_455 = phv_data_455; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_456 = phv_data_456; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_457 = phv_data_457; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_458 = phv_data_458; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_459 = phv_data_459; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_460 = phv_data_460; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_461 = phv_data_461; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_462 = phv_data_462; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_463 = phv_data_463; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_464 = phv_data_464; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_465 = phv_data_465; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_466 = phv_data_466; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_467 = phv_data_467; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_468 = phv_data_468; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_469 = phv_data_469; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_470 = phv_data_470; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_471 = phv_data_471; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_472 = phv_data_472; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_473 = phv_data_473; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_474 = phv_data_474; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_475 = phv_data_475; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_476 = phv_data_476; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_477 = phv_data_477; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_478 = phv_data_478; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_479 = phv_data_479; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_480 = phv_data_480; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_481 = phv_data_481; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_482 = phv_data_482; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_483 = phv_data_483; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_484 = phv_data_484; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_485 = phv_data_485; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_486 = phv_data_486; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_487 = phv_data_487; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_488 = phv_data_488; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_489 = phv_data_489; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_490 = phv_data_490; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_491 = phv_data_491; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_492 = phv_data_492; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_493 = phv_data_493; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_494 = phv_data_494; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_495 = phv_data_495; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_496 = phv_data_496; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_497 = phv_data_497; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_498 = phv_data_498; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_499 = phv_data_499; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_500 = phv_data_500; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_501 = phv_data_501; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_502 = phv_data_502; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_503 = phv_data_503; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_504 = phv_data_504; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_505 = phv_data_505; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_506 = phv_data_506; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_507 = phv_data_507; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_508 = phv_data_508; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_509 = phv_data_509; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_510 = phv_data_510; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_511 = phv_data_511; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[executor_pisa.scala 163:25]
  assign io_nid_out = nid; // @[executor_pisa.scala 173:20]
  assign io_tag_out_0 = opcode == 4'h9 ? 2'h2 : _GEN_12; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_1 = opcode_1 == 4'h9 ? 2'h2 : _GEN_91; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_2 = opcode_2 == 4'h9 ? 2'h2 : _GEN_170; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_3 = opcode_3 == 4'h9 ? 2'h2 : _GEN_249; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_4 = opcode_4 == 4'h9 ? 2'h2 : _GEN_328; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_5 = opcode_5 == 4'h9 ? 2'h2 : _GEN_407; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_6 = opcode_6 == 4'h9 ? 2'h2 : _GEN_486; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_7 = opcode_7 == 4'h9 ? 2'h2 : _GEN_565; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_8 = opcode_8 == 4'h9 ? 2'h2 : _GEN_644; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_9 = opcode_9 == 4'h9 ? 2'h2 : _GEN_723; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_10 = opcode_10 == 4'h9 ? 2'h2 : _GEN_802; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_11 = opcode_11 == 4'h9 ? 2'h2 : _GEN_881; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_12 = opcode_12 == 4'h9 ? 2'h2 : _GEN_960; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_13 = opcode_13 == 4'h9 ? 2'h2 : _GEN_1039; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_14 = opcode_14 == 4'h9 ? 2'h2 : _GEN_1118; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_15 = opcode_15 == 4'h9 ? 2'h2 : _GEN_1197; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_16 = opcode_16 == 4'h9 ? 2'h2 : _GEN_1276; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_17 = opcode_17 == 4'h9 ? 2'h2 : _GEN_1355; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_18 = opcode_18 == 4'h9 ? 2'h2 : _GEN_1434; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_19 = opcode_19 == 4'h9 ? 2'h2 : _GEN_1513; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_20 = opcode_20 == 4'h9 ? 2'h2 : _GEN_1592; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_21 = opcode_21 == 4'h9 ? 2'h2 : _GEN_1671; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_22 = opcode_22 == 4'h9 ? 2'h2 : _GEN_1750; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_23 = opcode_23 == 4'h9 ? 2'h2 : _GEN_1829; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_24 = opcode_24 == 4'h9 ? 2'h2 : _GEN_1908; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_25 = opcode_25 == 4'h9 ? 2'h2 : _GEN_1987; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_26 = opcode_26 == 4'h9 ? 2'h2 : _GEN_2066; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_27 = opcode_27 == 4'h9 ? 2'h2 : _GEN_2145; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_28 = opcode_28 == 4'h9 ? 2'h2 : _GEN_2224; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_29 = opcode_29 == 4'h9 ? 2'h2 : _GEN_2303; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_30 = opcode_30 == 4'h9 ? 2'h2 : _GEN_2382; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_31 = opcode_31 == 4'h9 ? 2'h2 : _GEN_2461; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_32 = opcode_32 == 4'h9 ? 2'h2 : _GEN_2540; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_33 = opcode_33 == 4'h9 ? 2'h2 : _GEN_2619; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_34 = opcode_34 == 4'h9 ? 2'h2 : _GEN_2698; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_35 = opcode_35 == 4'h9 ? 2'h2 : _GEN_2777; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_36 = opcode_36 == 4'h9 ? 2'h2 : _GEN_2856; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_37 = opcode_37 == 4'h9 ? 2'h2 : _GEN_2935; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_38 = opcode_38 == 4'h9 ? 2'h2 : _GEN_3014; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_39 = opcode_39 == 4'h9 ? 2'h2 : _GEN_3093; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_40 = opcode_40 == 4'h9 ? 2'h2 : _GEN_3172; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_41 = opcode_41 == 4'h9 ? 2'h2 : _GEN_3251; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_42 = opcode_42 == 4'h9 ? 2'h2 : _GEN_3330; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_43 = opcode_43 == 4'h9 ? 2'h2 : _GEN_3409; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_44 = opcode_44 == 4'h9 ? 2'h2 : _GEN_3488; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_45 = opcode_45 == 4'h9 ? 2'h2 : _GEN_3567; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_46 = opcode_46 == 4'h9 ? 2'h2 : _GEN_3646; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_47 = opcode_47 == 4'h9 ? 2'h2 : _GEN_3725; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_48 = opcode_48 == 4'h9 ? 2'h2 : _GEN_3804; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_49 = opcode_49 == 4'h9 ? 2'h2 : _GEN_3883; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_50 = opcode_50 == 4'h9 ? 2'h2 : _GEN_3962; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_51 = opcode_51 == 4'h9 ? 2'h2 : _GEN_4041; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_52 = opcode_52 == 4'h9 ? 2'h2 : _GEN_4120; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_53 = opcode_53 == 4'h9 ? 2'h2 : _GEN_4199; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_54 = opcode_54 == 4'h9 ? 2'h2 : _GEN_4278; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_55 = opcode_55 == 4'h9 ? 2'h2 : _GEN_4357; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_56 = opcode_56 == 4'h9 ? 2'h2 : _GEN_4436; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_57 = opcode_57 == 4'h9 ? 2'h2 : _GEN_4515; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_58 = opcode_58 == 4'h9 ? 2'h2 : _GEN_4594; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_59 = opcode_59 == 4'h9 ? 2'h2 : _GEN_4673; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_60 = opcode_60 == 4'h9 ? 2'h2 : _GEN_4752; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_61 = opcode_61 == 4'h9 ? 2'h2 : _GEN_4831; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_62 = opcode_62 == 4'h9 ? 2'h2 : _GEN_4910; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_63 = opcode_63 == 4'h9 ? 2'h2 : _GEN_4989; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_64 = opcode_64 == 4'h9 ? 2'h2 : _GEN_5077; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_65 = opcode_65 == 4'h9 ? 2'h2 : _GEN_5197; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_66 = opcode_66 == 4'h9 ? 2'h2 : _GEN_5317; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_67 = opcode_67 == 4'h9 ? 2'h2 : _GEN_5437; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_68 = opcode_68 == 4'h9 ? 2'h2 : _GEN_5557; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_69 = opcode_69 == 4'h9 ? 2'h2 : _GEN_5677; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_field_set_field8_0 = opcode == 4'h9 ? _GEN_76 : _GEN_11; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_1 = opcode_1 == 4'h9 ? _GEN_155 : _GEN_90; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_2 = opcode_2 == 4'h9 ? _GEN_234 : _GEN_169; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_3 = opcode_3 == 4'h9 ? _GEN_313 : _GEN_248; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_4 = opcode_4 == 4'h9 ? _GEN_392 : _GEN_327; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_5 = opcode_5 == 4'h9 ? _GEN_471 : _GEN_406; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_6 = opcode_6 == 4'h9 ? _GEN_550 : _GEN_485; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_7 = opcode_7 == 4'h9 ? _GEN_629 : _GEN_564; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_8 = opcode_8 == 4'h9 ? _GEN_708 : _GEN_643; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_9 = opcode_9 == 4'h9 ? _GEN_787 : _GEN_722; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_10 = opcode_10 == 4'h9 ? _GEN_866 : _GEN_801; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_11 = opcode_11 == 4'h9 ? _GEN_945 : _GEN_880; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_12 = opcode_12 == 4'h9 ? _GEN_1024 : _GEN_959; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_13 = opcode_13 == 4'h9 ? _GEN_1103 : _GEN_1038; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_14 = opcode_14 == 4'h9 ? _GEN_1182 : _GEN_1117; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_15 = opcode_15 == 4'h9 ? _GEN_1261 : _GEN_1196; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_16 = opcode_16 == 4'h9 ? _GEN_1340 : _GEN_1275; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_17 = opcode_17 == 4'h9 ? _GEN_1419 : _GEN_1354; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_18 = opcode_18 == 4'h9 ? _GEN_1498 : _GEN_1433; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_19 = opcode_19 == 4'h9 ? _GEN_1577 : _GEN_1512; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_20 = opcode_20 == 4'h9 ? _GEN_1656 : _GEN_1591; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_21 = opcode_21 == 4'h9 ? _GEN_1735 : _GEN_1670; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_22 = opcode_22 == 4'h9 ? _GEN_1814 : _GEN_1749; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_23 = opcode_23 == 4'h9 ? _GEN_1893 : _GEN_1828; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_24 = opcode_24 == 4'h9 ? _GEN_1972 : _GEN_1907; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_25 = opcode_25 == 4'h9 ? _GEN_2051 : _GEN_1986; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_26 = opcode_26 == 4'h9 ? _GEN_2130 : _GEN_2065; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_27 = opcode_27 == 4'h9 ? _GEN_2209 : _GEN_2144; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_28 = opcode_28 == 4'h9 ? _GEN_2288 : _GEN_2223; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_29 = opcode_29 == 4'h9 ? _GEN_2367 : _GEN_2302; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_30 = opcode_30 == 4'h9 ? _GEN_2446 : _GEN_2381; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_31 = opcode_31 == 4'h9 ? _GEN_2525 : _GEN_2460; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_32 = opcode_32 == 4'h9 ? _GEN_2604 : _GEN_2539; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_33 = opcode_33 == 4'h9 ? _GEN_2683 : _GEN_2618; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_34 = opcode_34 == 4'h9 ? _GEN_2762 : _GEN_2697; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_35 = opcode_35 == 4'h9 ? _GEN_2841 : _GEN_2776; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_36 = opcode_36 == 4'h9 ? _GEN_2920 : _GEN_2855; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_37 = opcode_37 == 4'h9 ? _GEN_2999 : _GEN_2934; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_38 = opcode_38 == 4'h9 ? _GEN_3078 : _GEN_3013; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_39 = opcode_39 == 4'h9 ? _GEN_3157 : _GEN_3092; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_40 = opcode_40 == 4'h9 ? _GEN_3236 : _GEN_3171; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_41 = opcode_41 == 4'h9 ? _GEN_3315 : _GEN_3250; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_42 = opcode_42 == 4'h9 ? _GEN_3394 : _GEN_3329; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_43 = opcode_43 == 4'h9 ? _GEN_3473 : _GEN_3408; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_44 = opcode_44 == 4'h9 ? _GEN_3552 : _GEN_3487; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_45 = opcode_45 == 4'h9 ? _GEN_3631 : _GEN_3566; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_46 = opcode_46 == 4'h9 ? _GEN_3710 : _GEN_3645; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_47 = opcode_47 == 4'h9 ? _GEN_3789 : _GEN_3724; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_48 = opcode_48 == 4'h9 ? _GEN_3868 : _GEN_3803; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_49 = opcode_49 == 4'h9 ? _GEN_3947 : _GEN_3882; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_50 = opcode_50 == 4'h9 ? _GEN_4026 : _GEN_3961; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_51 = opcode_51 == 4'h9 ? _GEN_4105 : _GEN_4040; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_52 = opcode_52 == 4'h9 ? _GEN_4184 : _GEN_4119; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_53 = opcode_53 == 4'h9 ? _GEN_4263 : _GEN_4198; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_54 = opcode_54 == 4'h9 ? _GEN_4342 : _GEN_4277; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_55 = opcode_55 == 4'h9 ? _GEN_4421 : _GEN_4356; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_56 = opcode_56 == 4'h9 ? _GEN_4500 : _GEN_4435; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_57 = opcode_57 == 4'h9 ? _GEN_4579 : _GEN_4514; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_58 = opcode_58 == 4'h9 ? _GEN_4658 : _GEN_4593; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_59 = opcode_59 == 4'h9 ? _GEN_4737 : _GEN_4672; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_60 = opcode_60 == 4'h9 ? _GEN_4816 : _GEN_4751; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_61 = opcode_61 == 4'h9 ? _GEN_4895 : _GEN_4830; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_62 = opcode_62 == 4'h9 ? _GEN_4974 : _GEN_4909; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_63 = opcode_63 == 4'h9 ? _GEN_5053 : _GEN_4988; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_0 = opcode_64 == 4'h9 ? _GEN_5173 : _GEN_5076; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_1 = opcode_65 == 4'h9 ? _GEN_5293 : _GEN_5196; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_2 = opcode_66 == 4'h9 ? _GEN_5413 : _GEN_5316; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_3 = opcode_67 == 4'h9 ? _GEN_5533 : _GEN_5436; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_4 = opcode_68 == 4'h9 ? _GEN_5653 : _GEN_5556; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_5 = opcode_69 == 4'h9 ? _GEN_5773 : _GEN_5676; // @[executor_pisa.scala 212:48]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[executor_pisa.scala 162:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[executor_pisa.scala 162:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[executor_pisa.scala 162:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[executor_pisa.scala 162:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[executor_pisa.scala 162:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[executor_pisa.scala 162:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[executor_pisa.scala 162:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[executor_pisa.scala 162:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[executor_pisa.scala 162:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[executor_pisa.scala 162:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[executor_pisa.scala 162:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[executor_pisa.scala 162:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[executor_pisa.scala 162:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[executor_pisa.scala 162:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[executor_pisa.scala 162:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[executor_pisa.scala 162:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[executor_pisa.scala 162:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[executor_pisa.scala 162:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[executor_pisa.scala 162:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[executor_pisa.scala 162:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[executor_pisa.scala 162:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[executor_pisa.scala 162:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[executor_pisa.scala 162:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[executor_pisa.scala 162:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[executor_pisa.scala 162:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[executor_pisa.scala 162:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[executor_pisa.scala 162:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[executor_pisa.scala 162:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[executor_pisa.scala 162:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[executor_pisa.scala 162:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[executor_pisa.scala 162:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[executor_pisa.scala 162:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[executor_pisa.scala 162:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[executor_pisa.scala 162:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[executor_pisa.scala 162:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[executor_pisa.scala 162:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[executor_pisa.scala 162:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[executor_pisa.scala 162:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[executor_pisa.scala 162:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[executor_pisa.scala 162:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[executor_pisa.scala 162:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[executor_pisa.scala 162:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[executor_pisa.scala 162:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[executor_pisa.scala 162:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[executor_pisa.scala 162:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[executor_pisa.scala 162:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[executor_pisa.scala 162:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[executor_pisa.scala 162:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[executor_pisa.scala 162:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[executor_pisa.scala 162:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[executor_pisa.scala 162:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[executor_pisa.scala 162:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[executor_pisa.scala 162:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[executor_pisa.scala 162:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[executor_pisa.scala 162:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[executor_pisa.scala 162:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[executor_pisa.scala 162:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[executor_pisa.scala 162:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[executor_pisa.scala 162:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[executor_pisa.scala 162:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[executor_pisa.scala 162:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[executor_pisa.scala 162:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[executor_pisa.scala 162:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[executor_pisa.scala 162:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[executor_pisa.scala 162:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[executor_pisa.scala 162:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[executor_pisa.scala 162:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[executor_pisa.scala 162:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[executor_pisa.scala 162:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[executor_pisa.scala 162:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[executor_pisa.scala 162:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[executor_pisa.scala 162:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[executor_pisa.scala 162:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[executor_pisa.scala 162:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[executor_pisa.scala 162:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[executor_pisa.scala 162:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[executor_pisa.scala 162:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[executor_pisa.scala 162:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[executor_pisa.scala 162:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[executor_pisa.scala 162:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[executor_pisa.scala 162:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[executor_pisa.scala 162:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[executor_pisa.scala 162:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[executor_pisa.scala 162:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[executor_pisa.scala 162:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[executor_pisa.scala 162:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[executor_pisa.scala 162:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[executor_pisa.scala 162:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[executor_pisa.scala 162:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[executor_pisa.scala 162:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[executor_pisa.scala 162:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[executor_pisa.scala 162:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[executor_pisa.scala 162:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[executor_pisa.scala 162:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[executor_pisa.scala 162:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[executor_pisa.scala 162:13]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[executor_pisa.scala 162:13]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[executor_pisa.scala 162:13]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[executor_pisa.scala 162:13]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[executor_pisa.scala 162:13]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[executor_pisa.scala 162:13]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[executor_pisa.scala 162:13]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[executor_pisa.scala 162:13]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[executor_pisa.scala 162:13]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[executor_pisa.scala 162:13]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[executor_pisa.scala 162:13]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[executor_pisa.scala 162:13]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[executor_pisa.scala 162:13]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[executor_pisa.scala 162:13]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[executor_pisa.scala 162:13]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[executor_pisa.scala 162:13]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[executor_pisa.scala 162:13]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[executor_pisa.scala 162:13]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[executor_pisa.scala 162:13]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[executor_pisa.scala 162:13]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[executor_pisa.scala 162:13]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[executor_pisa.scala 162:13]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[executor_pisa.scala 162:13]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[executor_pisa.scala 162:13]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[executor_pisa.scala 162:13]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[executor_pisa.scala 162:13]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[executor_pisa.scala 162:13]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[executor_pisa.scala 162:13]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[executor_pisa.scala 162:13]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[executor_pisa.scala 162:13]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[executor_pisa.scala 162:13]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[executor_pisa.scala 162:13]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[executor_pisa.scala 162:13]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[executor_pisa.scala 162:13]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[executor_pisa.scala 162:13]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[executor_pisa.scala 162:13]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[executor_pisa.scala 162:13]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[executor_pisa.scala 162:13]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[executor_pisa.scala 162:13]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[executor_pisa.scala 162:13]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[executor_pisa.scala 162:13]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[executor_pisa.scala 162:13]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[executor_pisa.scala 162:13]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[executor_pisa.scala 162:13]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[executor_pisa.scala 162:13]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[executor_pisa.scala 162:13]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[executor_pisa.scala 162:13]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[executor_pisa.scala 162:13]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[executor_pisa.scala 162:13]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[executor_pisa.scala 162:13]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[executor_pisa.scala 162:13]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[executor_pisa.scala 162:13]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[executor_pisa.scala 162:13]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[executor_pisa.scala 162:13]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[executor_pisa.scala 162:13]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[executor_pisa.scala 162:13]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[executor_pisa.scala 162:13]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[executor_pisa.scala 162:13]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[executor_pisa.scala 162:13]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[executor_pisa.scala 162:13]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[executor_pisa.scala 162:13]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[executor_pisa.scala 162:13]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[executor_pisa.scala 162:13]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[executor_pisa.scala 162:13]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[executor_pisa.scala 162:13]
    phv_data_160 <= io_pipe_phv_in_data_160; // @[executor_pisa.scala 162:13]
    phv_data_161 <= io_pipe_phv_in_data_161; // @[executor_pisa.scala 162:13]
    phv_data_162 <= io_pipe_phv_in_data_162; // @[executor_pisa.scala 162:13]
    phv_data_163 <= io_pipe_phv_in_data_163; // @[executor_pisa.scala 162:13]
    phv_data_164 <= io_pipe_phv_in_data_164; // @[executor_pisa.scala 162:13]
    phv_data_165 <= io_pipe_phv_in_data_165; // @[executor_pisa.scala 162:13]
    phv_data_166 <= io_pipe_phv_in_data_166; // @[executor_pisa.scala 162:13]
    phv_data_167 <= io_pipe_phv_in_data_167; // @[executor_pisa.scala 162:13]
    phv_data_168 <= io_pipe_phv_in_data_168; // @[executor_pisa.scala 162:13]
    phv_data_169 <= io_pipe_phv_in_data_169; // @[executor_pisa.scala 162:13]
    phv_data_170 <= io_pipe_phv_in_data_170; // @[executor_pisa.scala 162:13]
    phv_data_171 <= io_pipe_phv_in_data_171; // @[executor_pisa.scala 162:13]
    phv_data_172 <= io_pipe_phv_in_data_172; // @[executor_pisa.scala 162:13]
    phv_data_173 <= io_pipe_phv_in_data_173; // @[executor_pisa.scala 162:13]
    phv_data_174 <= io_pipe_phv_in_data_174; // @[executor_pisa.scala 162:13]
    phv_data_175 <= io_pipe_phv_in_data_175; // @[executor_pisa.scala 162:13]
    phv_data_176 <= io_pipe_phv_in_data_176; // @[executor_pisa.scala 162:13]
    phv_data_177 <= io_pipe_phv_in_data_177; // @[executor_pisa.scala 162:13]
    phv_data_178 <= io_pipe_phv_in_data_178; // @[executor_pisa.scala 162:13]
    phv_data_179 <= io_pipe_phv_in_data_179; // @[executor_pisa.scala 162:13]
    phv_data_180 <= io_pipe_phv_in_data_180; // @[executor_pisa.scala 162:13]
    phv_data_181 <= io_pipe_phv_in_data_181; // @[executor_pisa.scala 162:13]
    phv_data_182 <= io_pipe_phv_in_data_182; // @[executor_pisa.scala 162:13]
    phv_data_183 <= io_pipe_phv_in_data_183; // @[executor_pisa.scala 162:13]
    phv_data_184 <= io_pipe_phv_in_data_184; // @[executor_pisa.scala 162:13]
    phv_data_185 <= io_pipe_phv_in_data_185; // @[executor_pisa.scala 162:13]
    phv_data_186 <= io_pipe_phv_in_data_186; // @[executor_pisa.scala 162:13]
    phv_data_187 <= io_pipe_phv_in_data_187; // @[executor_pisa.scala 162:13]
    phv_data_188 <= io_pipe_phv_in_data_188; // @[executor_pisa.scala 162:13]
    phv_data_189 <= io_pipe_phv_in_data_189; // @[executor_pisa.scala 162:13]
    phv_data_190 <= io_pipe_phv_in_data_190; // @[executor_pisa.scala 162:13]
    phv_data_191 <= io_pipe_phv_in_data_191; // @[executor_pisa.scala 162:13]
    phv_data_192 <= io_pipe_phv_in_data_192; // @[executor_pisa.scala 162:13]
    phv_data_193 <= io_pipe_phv_in_data_193; // @[executor_pisa.scala 162:13]
    phv_data_194 <= io_pipe_phv_in_data_194; // @[executor_pisa.scala 162:13]
    phv_data_195 <= io_pipe_phv_in_data_195; // @[executor_pisa.scala 162:13]
    phv_data_196 <= io_pipe_phv_in_data_196; // @[executor_pisa.scala 162:13]
    phv_data_197 <= io_pipe_phv_in_data_197; // @[executor_pisa.scala 162:13]
    phv_data_198 <= io_pipe_phv_in_data_198; // @[executor_pisa.scala 162:13]
    phv_data_199 <= io_pipe_phv_in_data_199; // @[executor_pisa.scala 162:13]
    phv_data_200 <= io_pipe_phv_in_data_200; // @[executor_pisa.scala 162:13]
    phv_data_201 <= io_pipe_phv_in_data_201; // @[executor_pisa.scala 162:13]
    phv_data_202 <= io_pipe_phv_in_data_202; // @[executor_pisa.scala 162:13]
    phv_data_203 <= io_pipe_phv_in_data_203; // @[executor_pisa.scala 162:13]
    phv_data_204 <= io_pipe_phv_in_data_204; // @[executor_pisa.scala 162:13]
    phv_data_205 <= io_pipe_phv_in_data_205; // @[executor_pisa.scala 162:13]
    phv_data_206 <= io_pipe_phv_in_data_206; // @[executor_pisa.scala 162:13]
    phv_data_207 <= io_pipe_phv_in_data_207; // @[executor_pisa.scala 162:13]
    phv_data_208 <= io_pipe_phv_in_data_208; // @[executor_pisa.scala 162:13]
    phv_data_209 <= io_pipe_phv_in_data_209; // @[executor_pisa.scala 162:13]
    phv_data_210 <= io_pipe_phv_in_data_210; // @[executor_pisa.scala 162:13]
    phv_data_211 <= io_pipe_phv_in_data_211; // @[executor_pisa.scala 162:13]
    phv_data_212 <= io_pipe_phv_in_data_212; // @[executor_pisa.scala 162:13]
    phv_data_213 <= io_pipe_phv_in_data_213; // @[executor_pisa.scala 162:13]
    phv_data_214 <= io_pipe_phv_in_data_214; // @[executor_pisa.scala 162:13]
    phv_data_215 <= io_pipe_phv_in_data_215; // @[executor_pisa.scala 162:13]
    phv_data_216 <= io_pipe_phv_in_data_216; // @[executor_pisa.scala 162:13]
    phv_data_217 <= io_pipe_phv_in_data_217; // @[executor_pisa.scala 162:13]
    phv_data_218 <= io_pipe_phv_in_data_218; // @[executor_pisa.scala 162:13]
    phv_data_219 <= io_pipe_phv_in_data_219; // @[executor_pisa.scala 162:13]
    phv_data_220 <= io_pipe_phv_in_data_220; // @[executor_pisa.scala 162:13]
    phv_data_221 <= io_pipe_phv_in_data_221; // @[executor_pisa.scala 162:13]
    phv_data_222 <= io_pipe_phv_in_data_222; // @[executor_pisa.scala 162:13]
    phv_data_223 <= io_pipe_phv_in_data_223; // @[executor_pisa.scala 162:13]
    phv_data_224 <= io_pipe_phv_in_data_224; // @[executor_pisa.scala 162:13]
    phv_data_225 <= io_pipe_phv_in_data_225; // @[executor_pisa.scala 162:13]
    phv_data_226 <= io_pipe_phv_in_data_226; // @[executor_pisa.scala 162:13]
    phv_data_227 <= io_pipe_phv_in_data_227; // @[executor_pisa.scala 162:13]
    phv_data_228 <= io_pipe_phv_in_data_228; // @[executor_pisa.scala 162:13]
    phv_data_229 <= io_pipe_phv_in_data_229; // @[executor_pisa.scala 162:13]
    phv_data_230 <= io_pipe_phv_in_data_230; // @[executor_pisa.scala 162:13]
    phv_data_231 <= io_pipe_phv_in_data_231; // @[executor_pisa.scala 162:13]
    phv_data_232 <= io_pipe_phv_in_data_232; // @[executor_pisa.scala 162:13]
    phv_data_233 <= io_pipe_phv_in_data_233; // @[executor_pisa.scala 162:13]
    phv_data_234 <= io_pipe_phv_in_data_234; // @[executor_pisa.scala 162:13]
    phv_data_235 <= io_pipe_phv_in_data_235; // @[executor_pisa.scala 162:13]
    phv_data_236 <= io_pipe_phv_in_data_236; // @[executor_pisa.scala 162:13]
    phv_data_237 <= io_pipe_phv_in_data_237; // @[executor_pisa.scala 162:13]
    phv_data_238 <= io_pipe_phv_in_data_238; // @[executor_pisa.scala 162:13]
    phv_data_239 <= io_pipe_phv_in_data_239; // @[executor_pisa.scala 162:13]
    phv_data_240 <= io_pipe_phv_in_data_240; // @[executor_pisa.scala 162:13]
    phv_data_241 <= io_pipe_phv_in_data_241; // @[executor_pisa.scala 162:13]
    phv_data_242 <= io_pipe_phv_in_data_242; // @[executor_pisa.scala 162:13]
    phv_data_243 <= io_pipe_phv_in_data_243; // @[executor_pisa.scala 162:13]
    phv_data_244 <= io_pipe_phv_in_data_244; // @[executor_pisa.scala 162:13]
    phv_data_245 <= io_pipe_phv_in_data_245; // @[executor_pisa.scala 162:13]
    phv_data_246 <= io_pipe_phv_in_data_246; // @[executor_pisa.scala 162:13]
    phv_data_247 <= io_pipe_phv_in_data_247; // @[executor_pisa.scala 162:13]
    phv_data_248 <= io_pipe_phv_in_data_248; // @[executor_pisa.scala 162:13]
    phv_data_249 <= io_pipe_phv_in_data_249; // @[executor_pisa.scala 162:13]
    phv_data_250 <= io_pipe_phv_in_data_250; // @[executor_pisa.scala 162:13]
    phv_data_251 <= io_pipe_phv_in_data_251; // @[executor_pisa.scala 162:13]
    phv_data_252 <= io_pipe_phv_in_data_252; // @[executor_pisa.scala 162:13]
    phv_data_253 <= io_pipe_phv_in_data_253; // @[executor_pisa.scala 162:13]
    phv_data_254 <= io_pipe_phv_in_data_254; // @[executor_pisa.scala 162:13]
    phv_data_255 <= io_pipe_phv_in_data_255; // @[executor_pisa.scala 162:13]
    phv_data_256 <= io_pipe_phv_in_data_256; // @[executor_pisa.scala 162:13]
    phv_data_257 <= io_pipe_phv_in_data_257; // @[executor_pisa.scala 162:13]
    phv_data_258 <= io_pipe_phv_in_data_258; // @[executor_pisa.scala 162:13]
    phv_data_259 <= io_pipe_phv_in_data_259; // @[executor_pisa.scala 162:13]
    phv_data_260 <= io_pipe_phv_in_data_260; // @[executor_pisa.scala 162:13]
    phv_data_261 <= io_pipe_phv_in_data_261; // @[executor_pisa.scala 162:13]
    phv_data_262 <= io_pipe_phv_in_data_262; // @[executor_pisa.scala 162:13]
    phv_data_263 <= io_pipe_phv_in_data_263; // @[executor_pisa.scala 162:13]
    phv_data_264 <= io_pipe_phv_in_data_264; // @[executor_pisa.scala 162:13]
    phv_data_265 <= io_pipe_phv_in_data_265; // @[executor_pisa.scala 162:13]
    phv_data_266 <= io_pipe_phv_in_data_266; // @[executor_pisa.scala 162:13]
    phv_data_267 <= io_pipe_phv_in_data_267; // @[executor_pisa.scala 162:13]
    phv_data_268 <= io_pipe_phv_in_data_268; // @[executor_pisa.scala 162:13]
    phv_data_269 <= io_pipe_phv_in_data_269; // @[executor_pisa.scala 162:13]
    phv_data_270 <= io_pipe_phv_in_data_270; // @[executor_pisa.scala 162:13]
    phv_data_271 <= io_pipe_phv_in_data_271; // @[executor_pisa.scala 162:13]
    phv_data_272 <= io_pipe_phv_in_data_272; // @[executor_pisa.scala 162:13]
    phv_data_273 <= io_pipe_phv_in_data_273; // @[executor_pisa.scala 162:13]
    phv_data_274 <= io_pipe_phv_in_data_274; // @[executor_pisa.scala 162:13]
    phv_data_275 <= io_pipe_phv_in_data_275; // @[executor_pisa.scala 162:13]
    phv_data_276 <= io_pipe_phv_in_data_276; // @[executor_pisa.scala 162:13]
    phv_data_277 <= io_pipe_phv_in_data_277; // @[executor_pisa.scala 162:13]
    phv_data_278 <= io_pipe_phv_in_data_278; // @[executor_pisa.scala 162:13]
    phv_data_279 <= io_pipe_phv_in_data_279; // @[executor_pisa.scala 162:13]
    phv_data_280 <= io_pipe_phv_in_data_280; // @[executor_pisa.scala 162:13]
    phv_data_281 <= io_pipe_phv_in_data_281; // @[executor_pisa.scala 162:13]
    phv_data_282 <= io_pipe_phv_in_data_282; // @[executor_pisa.scala 162:13]
    phv_data_283 <= io_pipe_phv_in_data_283; // @[executor_pisa.scala 162:13]
    phv_data_284 <= io_pipe_phv_in_data_284; // @[executor_pisa.scala 162:13]
    phv_data_285 <= io_pipe_phv_in_data_285; // @[executor_pisa.scala 162:13]
    phv_data_286 <= io_pipe_phv_in_data_286; // @[executor_pisa.scala 162:13]
    phv_data_287 <= io_pipe_phv_in_data_287; // @[executor_pisa.scala 162:13]
    phv_data_288 <= io_pipe_phv_in_data_288; // @[executor_pisa.scala 162:13]
    phv_data_289 <= io_pipe_phv_in_data_289; // @[executor_pisa.scala 162:13]
    phv_data_290 <= io_pipe_phv_in_data_290; // @[executor_pisa.scala 162:13]
    phv_data_291 <= io_pipe_phv_in_data_291; // @[executor_pisa.scala 162:13]
    phv_data_292 <= io_pipe_phv_in_data_292; // @[executor_pisa.scala 162:13]
    phv_data_293 <= io_pipe_phv_in_data_293; // @[executor_pisa.scala 162:13]
    phv_data_294 <= io_pipe_phv_in_data_294; // @[executor_pisa.scala 162:13]
    phv_data_295 <= io_pipe_phv_in_data_295; // @[executor_pisa.scala 162:13]
    phv_data_296 <= io_pipe_phv_in_data_296; // @[executor_pisa.scala 162:13]
    phv_data_297 <= io_pipe_phv_in_data_297; // @[executor_pisa.scala 162:13]
    phv_data_298 <= io_pipe_phv_in_data_298; // @[executor_pisa.scala 162:13]
    phv_data_299 <= io_pipe_phv_in_data_299; // @[executor_pisa.scala 162:13]
    phv_data_300 <= io_pipe_phv_in_data_300; // @[executor_pisa.scala 162:13]
    phv_data_301 <= io_pipe_phv_in_data_301; // @[executor_pisa.scala 162:13]
    phv_data_302 <= io_pipe_phv_in_data_302; // @[executor_pisa.scala 162:13]
    phv_data_303 <= io_pipe_phv_in_data_303; // @[executor_pisa.scala 162:13]
    phv_data_304 <= io_pipe_phv_in_data_304; // @[executor_pisa.scala 162:13]
    phv_data_305 <= io_pipe_phv_in_data_305; // @[executor_pisa.scala 162:13]
    phv_data_306 <= io_pipe_phv_in_data_306; // @[executor_pisa.scala 162:13]
    phv_data_307 <= io_pipe_phv_in_data_307; // @[executor_pisa.scala 162:13]
    phv_data_308 <= io_pipe_phv_in_data_308; // @[executor_pisa.scala 162:13]
    phv_data_309 <= io_pipe_phv_in_data_309; // @[executor_pisa.scala 162:13]
    phv_data_310 <= io_pipe_phv_in_data_310; // @[executor_pisa.scala 162:13]
    phv_data_311 <= io_pipe_phv_in_data_311; // @[executor_pisa.scala 162:13]
    phv_data_312 <= io_pipe_phv_in_data_312; // @[executor_pisa.scala 162:13]
    phv_data_313 <= io_pipe_phv_in_data_313; // @[executor_pisa.scala 162:13]
    phv_data_314 <= io_pipe_phv_in_data_314; // @[executor_pisa.scala 162:13]
    phv_data_315 <= io_pipe_phv_in_data_315; // @[executor_pisa.scala 162:13]
    phv_data_316 <= io_pipe_phv_in_data_316; // @[executor_pisa.scala 162:13]
    phv_data_317 <= io_pipe_phv_in_data_317; // @[executor_pisa.scala 162:13]
    phv_data_318 <= io_pipe_phv_in_data_318; // @[executor_pisa.scala 162:13]
    phv_data_319 <= io_pipe_phv_in_data_319; // @[executor_pisa.scala 162:13]
    phv_data_320 <= io_pipe_phv_in_data_320; // @[executor_pisa.scala 162:13]
    phv_data_321 <= io_pipe_phv_in_data_321; // @[executor_pisa.scala 162:13]
    phv_data_322 <= io_pipe_phv_in_data_322; // @[executor_pisa.scala 162:13]
    phv_data_323 <= io_pipe_phv_in_data_323; // @[executor_pisa.scala 162:13]
    phv_data_324 <= io_pipe_phv_in_data_324; // @[executor_pisa.scala 162:13]
    phv_data_325 <= io_pipe_phv_in_data_325; // @[executor_pisa.scala 162:13]
    phv_data_326 <= io_pipe_phv_in_data_326; // @[executor_pisa.scala 162:13]
    phv_data_327 <= io_pipe_phv_in_data_327; // @[executor_pisa.scala 162:13]
    phv_data_328 <= io_pipe_phv_in_data_328; // @[executor_pisa.scala 162:13]
    phv_data_329 <= io_pipe_phv_in_data_329; // @[executor_pisa.scala 162:13]
    phv_data_330 <= io_pipe_phv_in_data_330; // @[executor_pisa.scala 162:13]
    phv_data_331 <= io_pipe_phv_in_data_331; // @[executor_pisa.scala 162:13]
    phv_data_332 <= io_pipe_phv_in_data_332; // @[executor_pisa.scala 162:13]
    phv_data_333 <= io_pipe_phv_in_data_333; // @[executor_pisa.scala 162:13]
    phv_data_334 <= io_pipe_phv_in_data_334; // @[executor_pisa.scala 162:13]
    phv_data_335 <= io_pipe_phv_in_data_335; // @[executor_pisa.scala 162:13]
    phv_data_336 <= io_pipe_phv_in_data_336; // @[executor_pisa.scala 162:13]
    phv_data_337 <= io_pipe_phv_in_data_337; // @[executor_pisa.scala 162:13]
    phv_data_338 <= io_pipe_phv_in_data_338; // @[executor_pisa.scala 162:13]
    phv_data_339 <= io_pipe_phv_in_data_339; // @[executor_pisa.scala 162:13]
    phv_data_340 <= io_pipe_phv_in_data_340; // @[executor_pisa.scala 162:13]
    phv_data_341 <= io_pipe_phv_in_data_341; // @[executor_pisa.scala 162:13]
    phv_data_342 <= io_pipe_phv_in_data_342; // @[executor_pisa.scala 162:13]
    phv_data_343 <= io_pipe_phv_in_data_343; // @[executor_pisa.scala 162:13]
    phv_data_344 <= io_pipe_phv_in_data_344; // @[executor_pisa.scala 162:13]
    phv_data_345 <= io_pipe_phv_in_data_345; // @[executor_pisa.scala 162:13]
    phv_data_346 <= io_pipe_phv_in_data_346; // @[executor_pisa.scala 162:13]
    phv_data_347 <= io_pipe_phv_in_data_347; // @[executor_pisa.scala 162:13]
    phv_data_348 <= io_pipe_phv_in_data_348; // @[executor_pisa.scala 162:13]
    phv_data_349 <= io_pipe_phv_in_data_349; // @[executor_pisa.scala 162:13]
    phv_data_350 <= io_pipe_phv_in_data_350; // @[executor_pisa.scala 162:13]
    phv_data_351 <= io_pipe_phv_in_data_351; // @[executor_pisa.scala 162:13]
    phv_data_352 <= io_pipe_phv_in_data_352; // @[executor_pisa.scala 162:13]
    phv_data_353 <= io_pipe_phv_in_data_353; // @[executor_pisa.scala 162:13]
    phv_data_354 <= io_pipe_phv_in_data_354; // @[executor_pisa.scala 162:13]
    phv_data_355 <= io_pipe_phv_in_data_355; // @[executor_pisa.scala 162:13]
    phv_data_356 <= io_pipe_phv_in_data_356; // @[executor_pisa.scala 162:13]
    phv_data_357 <= io_pipe_phv_in_data_357; // @[executor_pisa.scala 162:13]
    phv_data_358 <= io_pipe_phv_in_data_358; // @[executor_pisa.scala 162:13]
    phv_data_359 <= io_pipe_phv_in_data_359; // @[executor_pisa.scala 162:13]
    phv_data_360 <= io_pipe_phv_in_data_360; // @[executor_pisa.scala 162:13]
    phv_data_361 <= io_pipe_phv_in_data_361; // @[executor_pisa.scala 162:13]
    phv_data_362 <= io_pipe_phv_in_data_362; // @[executor_pisa.scala 162:13]
    phv_data_363 <= io_pipe_phv_in_data_363; // @[executor_pisa.scala 162:13]
    phv_data_364 <= io_pipe_phv_in_data_364; // @[executor_pisa.scala 162:13]
    phv_data_365 <= io_pipe_phv_in_data_365; // @[executor_pisa.scala 162:13]
    phv_data_366 <= io_pipe_phv_in_data_366; // @[executor_pisa.scala 162:13]
    phv_data_367 <= io_pipe_phv_in_data_367; // @[executor_pisa.scala 162:13]
    phv_data_368 <= io_pipe_phv_in_data_368; // @[executor_pisa.scala 162:13]
    phv_data_369 <= io_pipe_phv_in_data_369; // @[executor_pisa.scala 162:13]
    phv_data_370 <= io_pipe_phv_in_data_370; // @[executor_pisa.scala 162:13]
    phv_data_371 <= io_pipe_phv_in_data_371; // @[executor_pisa.scala 162:13]
    phv_data_372 <= io_pipe_phv_in_data_372; // @[executor_pisa.scala 162:13]
    phv_data_373 <= io_pipe_phv_in_data_373; // @[executor_pisa.scala 162:13]
    phv_data_374 <= io_pipe_phv_in_data_374; // @[executor_pisa.scala 162:13]
    phv_data_375 <= io_pipe_phv_in_data_375; // @[executor_pisa.scala 162:13]
    phv_data_376 <= io_pipe_phv_in_data_376; // @[executor_pisa.scala 162:13]
    phv_data_377 <= io_pipe_phv_in_data_377; // @[executor_pisa.scala 162:13]
    phv_data_378 <= io_pipe_phv_in_data_378; // @[executor_pisa.scala 162:13]
    phv_data_379 <= io_pipe_phv_in_data_379; // @[executor_pisa.scala 162:13]
    phv_data_380 <= io_pipe_phv_in_data_380; // @[executor_pisa.scala 162:13]
    phv_data_381 <= io_pipe_phv_in_data_381; // @[executor_pisa.scala 162:13]
    phv_data_382 <= io_pipe_phv_in_data_382; // @[executor_pisa.scala 162:13]
    phv_data_383 <= io_pipe_phv_in_data_383; // @[executor_pisa.scala 162:13]
    phv_data_384 <= io_pipe_phv_in_data_384; // @[executor_pisa.scala 162:13]
    phv_data_385 <= io_pipe_phv_in_data_385; // @[executor_pisa.scala 162:13]
    phv_data_386 <= io_pipe_phv_in_data_386; // @[executor_pisa.scala 162:13]
    phv_data_387 <= io_pipe_phv_in_data_387; // @[executor_pisa.scala 162:13]
    phv_data_388 <= io_pipe_phv_in_data_388; // @[executor_pisa.scala 162:13]
    phv_data_389 <= io_pipe_phv_in_data_389; // @[executor_pisa.scala 162:13]
    phv_data_390 <= io_pipe_phv_in_data_390; // @[executor_pisa.scala 162:13]
    phv_data_391 <= io_pipe_phv_in_data_391; // @[executor_pisa.scala 162:13]
    phv_data_392 <= io_pipe_phv_in_data_392; // @[executor_pisa.scala 162:13]
    phv_data_393 <= io_pipe_phv_in_data_393; // @[executor_pisa.scala 162:13]
    phv_data_394 <= io_pipe_phv_in_data_394; // @[executor_pisa.scala 162:13]
    phv_data_395 <= io_pipe_phv_in_data_395; // @[executor_pisa.scala 162:13]
    phv_data_396 <= io_pipe_phv_in_data_396; // @[executor_pisa.scala 162:13]
    phv_data_397 <= io_pipe_phv_in_data_397; // @[executor_pisa.scala 162:13]
    phv_data_398 <= io_pipe_phv_in_data_398; // @[executor_pisa.scala 162:13]
    phv_data_399 <= io_pipe_phv_in_data_399; // @[executor_pisa.scala 162:13]
    phv_data_400 <= io_pipe_phv_in_data_400; // @[executor_pisa.scala 162:13]
    phv_data_401 <= io_pipe_phv_in_data_401; // @[executor_pisa.scala 162:13]
    phv_data_402 <= io_pipe_phv_in_data_402; // @[executor_pisa.scala 162:13]
    phv_data_403 <= io_pipe_phv_in_data_403; // @[executor_pisa.scala 162:13]
    phv_data_404 <= io_pipe_phv_in_data_404; // @[executor_pisa.scala 162:13]
    phv_data_405 <= io_pipe_phv_in_data_405; // @[executor_pisa.scala 162:13]
    phv_data_406 <= io_pipe_phv_in_data_406; // @[executor_pisa.scala 162:13]
    phv_data_407 <= io_pipe_phv_in_data_407; // @[executor_pisa.scala 162:13]
    phv_data_408 <= io_pipe_phv_in_data_408; // @[executor_pisa.scala 162:13]
    phv_data_409 <= io_pipe_phv_in_data_409; // @[executor_pisa.scala 162:13]
    phv_data_410 <= io_pipe_phv_in_data_410; // @[executor_pisa.scala 162:13]
    phv_data_411 <= io_pipe_phv_in_data_411; // @[executor_pisa.scala 162:13]
    phv_data_412 <= io_pipe_phv_in_data_412; // @[executor_pisa.scala 162:13]
    phv_data_413 <= io_pipe_phv_in_data_413; // @[executor_pisa.scala 162:13]
    phv_data_414 <= io_pipe_phv_in_data_414; // @[executor_pisa.scala 162:13]
    phv_data_415 <= io_pipe_phv_in_data_415; // @[executor_pisa.scala 162:13]
    phv_data_416 <= io_pipe_phv_in_data_416; // @[executor_pisa.scala 162:13]
    phv_data_417 <= io_pipe_phv_in_data_417; // @[executor_pisa.scala 162:13]
    phv_data_418 <= io_pipe_phv_in_data_418; // @[executor_pisa.scala 162:13]
    phv_data_419 <= io_pipe_phv_in_data_419; // @[executor_pisa.scala 162:13]
    phv_data_420 <= io_pipe_phv_in_data_420; // @[executor_pisa.scala 162:13]
    phv_data_421 <= io_pipe_phv_in_data_421; // @[executor_pisa.scala 162:13]
    phv_data_422 <= io_pipe_phv_in_data_422; // @[executor_pisa.scala 162:13]
    phv_data_423 <= io_pipe_phv_in_data_423; // @[executor_pisa.scala 162:13]
    phv_data_424 <= io_pipe_phv_in_data_424; // @[executor_pisa.scala 162:13]
    phv_data_425 <= io_pipe_phv_in_data_425; // @[executor_pisa.scala 162:13]
    phv_data_426 <= io_pipe_phv_in_data_426; // @[executor_pisa.scala 162:13]
    phv_data_427 <= io_pipe_phv_in_data_427; // @[executor_pisa.scala 162:13]
    phv_data_428 <= io_pipe_phv_in_data_428; // @[executor_pisa.scala 162:13]
    phv_data_429 <= io_pipe_phv_in_data_429; // @[executor_pisa.scala 162:13]
    phv_data_430 <= io_pipe_phv_in_data_430; // @[executor_pisa.scala 162:13]
    phv_data_431 <= io_pipe_phv_in_data_431; // @[executor_pisa.scala 162:13]
    phv_data_432 <= io_pipe_phv_in_data_432; // @[executor_pisa.scala 162:13]
    phv_data_433 <= io_pipe_phv_in_data_433; // @[executor_pisa.scala 162:13]
    phv_data_434 <= io_pipe_phv_in_data_434; // @[executor_pisa.scala 162:13]
    phv_data_435 <= io_pipe_phv_in_data_435; // @[executor_pisa.scala 162:13]
    phv_data_436 <= io_pipe_phv_in_data_436; // @[executor_pisa.scala 162:13]
    phv_data_437 <= io_pipe_phv_in_data_437; // @[executor_pisa.scala 162:13]
    phv_data_438 <= io_pipe_phv_in_data_438; // @[executor_pisa.scala 162:13]
    phv_data_439 <= io_pipe_phv_in_data_439; // @[executor_pisa.scala 162:13]
    phv_data_440 <= io_pipe_phv_in_data_440; // @[executor_pisa.scala 162:13]
    phv_data_441 <= io_pipe_phv_in_data_441; // @[executor_pisa.scala 162:13]
    phv_data_442 <= io_pipe_phv_in_data_442; // @[executor_pisa.scala 162:13]
    phv_data_443 <= io_pipe_phv_in_data_443; // @[executor_pisa.scala 162:13]
    phv_data_444 <= io_pipe_phv_in_data_444; // @[executor_pisa.scala 162:13]
    phv_data_445 <= io_pipe_phv_in_data_445; // @[executor_pisa.scala 162:13]
    phv_data_446 <= io_pipe_phv_in_data_446; // @[executor_pisa.scala 162:13]
    phv_data_447 <= io_pipe_phv_in_data_447; // @[executor_pisa.scala 162:13]
    phv_data_448 <= io_pipe_phv_in_data_448; // @[executor_pisa.scala 162:13]
    phv_data_449 <= io_pipe_phv_in_data_449; // @[executor_pisa.scala 162:13]
    phv_data_450 <= io_pipe_phv_in_data_450; // @[executor_pisa.scala 162:13]
    phv_data_451 <= io_pipe_phv_in_data_451; // @[executor_pisa.scala 162:13]
    phv_data_452 <= io_pipe_phv_in_data_452; // @[executor_pisa.scala 162:13]
    phv_data_453 <= io_pipe_phv_in_data_453; // @[executor_pisa.scala 162:13]
    phv_data_454 <= io_pipe_phv_in_data_454; // @[executor_pisa.scala 162:13]
    phv_data_455 <= io_pipe_phv_in_data_455; // @[executor_pisa.scala 162:13]
    phv_data_456 <= io_pipe_phv_in_data_456; // @[executor_pisa.scala 162:13]
    phv_data_457 <= io_pipe_phv_in_data_457; // @[executor_pisa.scala 162:13]
    phv_data_458 <= io_pipe_phv_in_data_458; // @[executor_pisa.scala 162:13]
    phv_data_459 <= io_pipe_phv_in_data_459; // @[executor_pisa.scala 162:13]
    phv_data_460 <= io_pipe_phv_in_data_460; // @[executor_pisa.scala 162:13]
    phv_data_461 <= io_pipe_phv_in_data_461; // @[executor_pisa.scala 162:13]
    phv_data_462 <= io_pipe_phv_in_data_462; // @[executor_pisa.scala 162:13]
    phv_data_463 <= io_pipe_phv_in_data_463; // @[executor_pisa.scala 162:13]
    phv_data_464 <= io_pipe_phv_in_data_464; // @[executor_pisa.scala 162:13]
    phv_data_465 <= io_pipe_phv_in_data_465; // @[executor_pisa.scala 162:13]
    phv_data_466 <= io_pipe_phv_in_data_466; // @[executor_pisa.scala 162:13]
    phv_data_467 <= io_pipe_phv_in_data_467; // @[executor_pisa.scala 162:13]
    phv_data_468 <= io_pipe_phv_in_data_468; // @[executor_pisa.scala 162:13]
    phv_data_469 <= io_pipe_phv_in_data_469; // @[executor_pisa.scala 162:13]
    phv_data_470 <= io_pipe_phv_in_data_470; // @[executor_pisa.scala 162:13]
    phv_data_471 <= io_pipe_phv_in_data_471; // @[executor_pisa.scala 162:13]
    phv_data_472 <= io_pipe_phv_in_data_472; // @[executor_pisa.scala 162:13]
    phv_data_473 <= io_pipe_phv_in_data_473; // @[executor_pisa.scala 162:13]
    phv_data_474 <= io_pipe_phv_in_data_474; // @[executor_pisa.scala 162:13]
    phv_data_475 <= io_pipe_phv_in_data_475; // @[executor_pisa.scala 162:13]
    phv_data_476 <= io_pipe_phv_in_data_476; // @[executor_pisa.scala 162:13]
    phv_data_477 <= io_pipe_phv_in_data_477; // @[executor_pisa.scala 162:13]
    phv_data_478 <= io_pipe_phv_in_data_478; // @[executor_pisa.scala 162:13]
    phv_data_479 <= io_pipe_phv_in_data_479; // @[executor_pisa.scala 162:13]
    phv_data_480 <= io_pipe_phv_in_data_480; // @[executor_pisa.scala 162:13]
    phv_data_481 <= io_pipe_phv_in_data_481; // @[executor_pisa.scala 162:13]
    phv_data_482 <= io_pipe_phv_in_data_482; // @[executor_pisa.scala 162:13]
    phv_data_483 <= io_pipe_phv_in_data_483; // @[executor_pisa.scala 162:13]
    phv_data_484 <= io_pipe_phv_in_data_484; // @[executor_pisa.scala 162:13]
    phv_data_485 <= io_pipe_phv_in_data_485; // @[executor_pisa.scala 162:13]
    phv_data_486 <= io_pipe_phv_in_data_486; // @[executor_pisa.scala 162:13]
    phv_data_487 <= io_pipe_phv_in_data_487; // @[executor_pisa.scala 162:13]
    phv_data_488 <= io_pipe_phv_in_data_488; // @[executor_pisa.scala 162:13]
    phv_data_489 <= io_pipe_phv_in_data_489; // @[executor_pisa.scala 162:13]
    phv_data_490 <= io_pipe_phv_in_data_490; // @[executor_pisa.scala 162:13]
    phv_data_491 <= io_pipe_phv_in_data_491; // @[executor_pisa.scala 162:13]
    phv_data_492 <= io_pipe_phv_in_data_492; // @[executor_pisa.scala 162:13]
    phv_data_493 <= io_pipe_phv_in_data_493; // @[executor_pisa.scala 162:13]
    phv_data_494 <= io_pipe_phv_in_data_494; // @[executor_pisa.scala 162:13]
    phv_data_495 <= io_pipe_phv_in_data_495; // @[executor_pisa.scala 162:13]
    phv_data_496 <= io_pipe_phv_in_data_496; // @[executor_pisa.scala 162:13]
    phv_data_497 <= io_pipe_phv_in_data_497; // @[executor_pisa.scala 162:13]
    phv_data_498 <= io_pipe_phv_in_data_498; // @[executor_pisa.scala 162:13]
    phv_data_499 <= io_pipe_phv_in_data_499; // @[executor_pisa.scala 162:13]
    phv_data_500 <= io_pipe_phv_in_data_500; // @[executor_pisa.scala 162:13]
    phv_data_501 <= io_pipe_phv_in_data_501; // @[executor_pisa.scala 162:13]
    phv_data_502 <= io_pipe_phv_in_data_502; // @[executor_pisa.scala 162:13]
    phv_data_503 <= io_pipe_phv_in_data_503; // @[executor_pisa.scala 162:13]
    phv_data_504 <= io_pipe_phv_in_data_504; // @[executor_pisa.scala 162:13]
    phv_data_505 <= io_pipe_phv_in_data_505; // @[executor_pisa.scala 162:13]
    phv_data_506 <= io_pipe_phv_in_data_506; // @[executor_pisa.scala 162:13]
    phv_data_507 <= io_pipe_phv_in_data_507; // @[executor_pisa.scala 162:13]
    phv_data_508 <= io_pipe_phv_in_data_508; // @[executor_pisa.scala 162:13]
    phv_data_509 <= io_pipe_phv_in_data_509; // @[executor_pisa.scala 162:13]
    phv_data_510 <= io_pipe_phv_in_data_510; // @[executor_pisa.scala 162:13]
    phv_data_511 <= io_pipe_phv_in_data_511; // @[executor_pisa.scala 162:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[executor_pisa.scala 162:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[executor_pisa.scala 162:13]
    args_0 <= io_args_in_0; // @[executor_pisa.scala 166:14]
    args_1 <= io_args_in_1; // @[executor_pisa.scala 166:14]
    args_2 <= io_args_in_2; // @[executor_pisa.scala 166:14]
    args_3 <= io_args_in_3; // @[executor_pisa.scala 166:14]
    args_4 <= io_args_in_4; // @[executor_pisa.scala 166:14]
    args_5 <= io_args_in_5; // @[executor_pisa.scala 166:14]
    args_6 <= io_args_in_6; // @[executor_pisa.scala 166:14]
    vliw_0 <= io_vliw_in_0; // @[executor_pisa.scala 169:14]
    vliw_1 <= io_vliw_in_1; // @[executor_pisa.scala 169:14]
    vliw_2 <= io_vliw_in_2; // @[executor_pisa.scala 169:14]
    vliw_3 <= io_vliw_in_3; // @[executor_pisa.scala 169:14]
    vliw_4 <= io_vliw_in_4; // @[executor_pisa.scala 169:14]
    vliw_5 <= io_vliw_in_5; // @[executor_pisa.scala 169:14]
    vliw_6 <= io_vliw_in_6; // @[executor_pisa.scala 169:14]
    vliw_7 <= io_vliw_in_7; // @[executor_pisa.scala 169:14]
    vliw_8 <= io_vliw_in_8; // @[executor_pisa.scala 169:14]
    vliw_9 <= io_vliw_in_9; // @[executor_pisa.scala 169:14]
    vliw_10 <= io_vliw_in_10; // @[executor_pisa.scala 169:14]
    vliw_11 <= io_vliw_in_11; // @[executor_pisa.scala 169:14]
    vliw_12 <= io_vliw_in_12; // @[executor_pisa.scala 169:14]
    vliw_13 <= io_vliw_in_13; // @[executor_pisa.scala 169:14]
    vliw_14 <= io_vliw_in_14; // @[executor_pisa.scala 169:14]
    vliw_15 <= io_vliw_in_15; // @[executor_pisa.scala 169:14]
    vliw_16 <= io_vliw_in_16; // @[executor_pisa.scala 169:14]
    vliw_17 <= io_vliw_in_17; // @[executor_pisa.scala 169:14]
    vliw_18 <= io_vliw_in_18; // @[executor_pisa.scala 169:14]
    vliw_19 <= io_vliw_in_19; // @[executor_pisa.scala 169:14]
    vliw_20 <= io_vliw_in_20; // @[executor_pisa.scala 169:14]
    vliw_21 <= io_vliw_in_21; // @[executor_pisa.scala 169:14]
    vliw_22 <= io_vliw_in_22; // @[executor_pisa.scala 169:14]
    vliw_23 <= io_vliw_in_23; // @[executor_pisa.scala 169:14]
    vliw_24 <= io_vliw_in_24; // @[executor_pisa.scala 169:14]
    vliw_25 <= io_vliw_in_25; // @[executor_pisa.scala 169:14]
    vliw_26 <= io_vliw_in_26; // @[executor_pisa.scala 169:14]
    vliw_27 <= io_vliw_in_27; // @[executor_pisa.scala 169:14]
    vliw_28 <= io_vliw_in_28; // @[executor_pisa.scala 169:14]
    vliw_29 <= io_vliw_in_29; // @[executor_pisa.scala 169:14]
    vliw_30 <= io_vliw_in_30; // @[executor_pisa.scala 169:14]
    vliw_31 <= io_vliw_in_31; // @[executor_pisa.scala 169:14]
    vliw_32 <= io_vliw_in_32; // @[executor_pisa.scala 169:14]
    vliw_33 <= io_vliw_in_33; // @[executor_pisa.scala 169:14]
    vliw_34 <= io_vliw_in_34; // @[executor_pisa.scala 169:14]
    vliw_35 <= io_vliw_in_35; // @[executor_pisa.scala 169:14]
    vliw_36 <= io_vliw_in_36; // @[executor_pisa.scala 169:14]
    vliw_37 <= io_vliw_in_37; // @[executor_pisa.scala 169:14]
    vliw_38 <= io_vliw_in_38; // @[executor_pisa.scala 169:14]
    vliw_39 <= io_vliw_in_39; // @[executor_pisa.scala 169:14]
    vliw_40 <= io_vliw_in_40; // @[executor_pisa.scala 169:14]
    vliw_41 <= io_vliw_in_41; // @[executor_pisa.scala 169:14]
    vliw_42 <= io_vliw_in_42; // @[executor_pisa.scala 169:14]
    vliw_43 <= io_vliw_in_43; // @[executor_pisa.scala 169:14]
    vliw_44 <= io_vliw_in_44; // @[executor_pisa.scala 169:14]
    vliw_45 <= io_vliw_in_45; // @[executor_pisa.scala 169:14]
    vliw_46 <= io_vliw_in_46; // @[executor_pisa.scala 169:14]
    vliw_47 <= io_vliw_in_47; // @[executor_pisa.scala 169:14]
    vliw_48 <= io_vliw_in_48; // @[executor_pisa.scala 169:14]
    vliw_49 <= io_vliw_in_49; // @[executor_pisa.scala 169:14]
    vliw_50 <= io_vliw_in_50; // @[executor_pisa.scala 169:14]
    vliw_51 <= io_vliw_in_51; // @[executor_pisa.scala 169:14]
    vliw_52 <= io_vliw_in_52; // @[executor_pisa.scala 169:14]
    vliw_53 <= io_vliw_in_53; // @[executor_pisa.scala 169:14]
    vliw_54 <= io_vliw_in_54; // @[executor_pisa.scala 169:14]
    vliw_55 <= io_vliw_in_55; // @[executor_pisa.scala 169:14]
    vliw_56 <= io_vliw_in_56; // @[executor_pisa.scala 169:14]
    vliw_57 <= io_vliw_in_57; // @[executor_pisa.scala 169:14]
    vliw_58 <= io_vliw_in_58; // @[executor_pisa.scala 169:14]
    vliw_59 <= io_vliw_in_59; // @[executor_pisa.scala 169:14]
    vliw_60 <= io_vliw_in_60; // @[executor_pisa.scala 169:14]
    vliw_61 <= io_vliw_in_61; // @[executor_pisa.scala 169:14]
    vliw_62 <= io_vliw_in_62; // @[executor_pisa.scala 169:14]
    vliw_63 <= io_vliw_in_63; // @[executor_pisa.scala 169:14]
    vliw_64 <= io_vliw_in_64; // @[executor_pisa.scala 169:14]
    vliw_65 <= io_vliw_in_65; // @[executor_pisa.scala 169:14]
    vliw_66 <= io_vliw_in_66; // @[executor_pisa.scala 169:14]
    vliw_67 <= io_vliw_in_67; // @[executor_pisa.scala 169:14]
    vliw_68 <= io_vliw_in_68; // @[executor_pisa.scala 169:14]
    vliw_69 <= io_vliw_in_69; // @[executor_pisa.scala 169:14]
    nid <= io_nid_in; // @[executor_pisa.scala 172:13]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_data_160 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  phv_data_161 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  phv_data_162 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  phv_data_163 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  phv_data_164 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  phv_data_165 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  phv_data_166 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  phv_data_167 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  phv_data_168 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  phv_data_169 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  phv_data_170 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  phv_data_171 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  phv_data_172 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  phv_data_173 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  phv_data_174 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  phv_data_175 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  phv_data_176 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_data_177 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_data_178 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  phv_data_179 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  phv_data_180 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  phv_data_181 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  phv_data_182 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  phv_data_183 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  phv_data_184 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  phv_data_185 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  phv_data_186 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  phv_data_187 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  phv_data_188 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  phv_data_189 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  phv_data_190 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  phv_data_191 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  phv_data_192 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  phv_data_193 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  phv_data_194 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  phv_data_195 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  phv_data_196 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  phv_data_197 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  phv_data_198 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  phv_data_199 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  phv_data_200 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  phv_data_201 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  phv_data_202 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  phv_data_203 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  phv_data_204 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  phv_data_205 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  phv_data_206 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  phv_data_207 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  phv_data_208 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  phv_data_209 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  phv_data_210 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  phv_data_211 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  phv_data_212 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  phv_data_213 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  phv_data_214 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  phv_data_215 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  phv_data_216 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  phv_data_217 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  phv_data_218 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  phv_data_219 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  phv_data_220 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  phv_data_221 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  phv_data_222 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  phv_data_223 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  phv_data_224 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  phv_data_225 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  phv_data_226 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  phv_data_227 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  phv_data_228 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  phv_data_229 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  phv_data_230 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  phv_data_231 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  phv_data_232 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  phv_data_233 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  phv_data_234 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  phv_data_235 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  phv_data_236 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  phv_data_237 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  phv_data_238 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  phv_data_239 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  phv_data_240 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  phv_data_241 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  phv_data_242 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  phv_data_243 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  phv_data_244 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  phv_data_245 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  phv_data_246 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  phv_data_247 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  phv_data_248 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  phv_data_249 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  phv_data_250 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  phv_data_251 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  phv_data_252 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  phv_data_253 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  phv_data_254 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  phv_data_255 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  phv_data_256 = _RAND_256[7:0];
  _RAND_257 = {1{`RANDOM}};
  phv_data_257 = _RAND_257[7:0];
  _RAND_258 = {1{`RANDOM}};
  phv_data_258 = _RAND_258[7:0];
  _RAND_259 = {1{`RANDOM}};
  phv_data_259 = _RAND_259[7:0];
  _RAND_260 = {1{`RANDOM}};
  phv_data_260 = _RAND_260[7:0];
  _RAND_261 = {1{`RANDOM}};
  phv_data_261 = _RAND_261[7:0];
  _RAND_262 = {1{`RANDOM}};
  phv_data_262 = _RAND_262[7:0];
  _RAND_263 = {1{`RANDOM}};
  phv_data_263 = _RAND_263[7:0];
  _RAND_264 = {1{`RANDOM}};
  phv_data_264 = _RAND_264[7:0];
  _RAND_265 = {1{`RANDOM}};
  phv_data_265 = _RAND_265[7:0];
  _RAND_266 = {1{`RANDOM}};
  phv_data_266 = _RAND_266[7:0];
  _RAND_267 = {1{`RANDOM}};
  phv_data_267 = _RAND_267[7:0];
  _RAND_268 = {1{`RANDOM}};
  phv_data_268 = _RAND_268[7:0];
  _RAND_269 = {1{`RANDOM}};
  phv_data_269 = _RAND_269[7:0];
  _RAND_270 = {1{`RANDOM}};
  phv_data_270 = _RAND_270[7:0];
  _RAND_271 = {1{`RANDOM}};
  phv_data_271 = _RAND_271[7:0];
  _RAND_272 = {1{`RANDOM}};
  phv_data_272 = _RAND_272[7:0];
  _RAND_273 = {1{`RANDOM}};
  phv_data_273 = _RAND_273[7:0];
  _RAND_274 = {1{`RANDOM}};
  phv_data_274 = _RAND_274[7:0];
  _RAND_275 = {1{`RANDOM}};
  phv_data_275 = _RAND_275[7:0];
  _RAND_276 = {1{`RANDOM}};
  phv_data_276 = _RAND_276[7:0];
  _RAND_277 = {1{`RANDOM}};
  phv_data_277 = _RAND_277[7:0];
  _RAND_278 = {1{`RANDOM}};
  phv_data_278 = _RAND_278[7:0];
  _RAND_279 = {1{`RANDOM}};
  phv_data_279 = _RAND_279[7:0];
  _RAND_280 = {1{`RANDOM}};
  phv_data_280 = _RAND_280[7:0];
  _RAND_281 = {1{`RANDOM}};
  phv_data_281 = _RAND_281[7:0];
  _RAND_282 = {1{`RANDOM}};
  phv_data_282 = _RAND_282[7:0];
  _RAND_283 = {1{`RANDOM}};
  phv_data_283 = _RAND_283[7:0];
  _RAND_284 = {1{`RANDOM}};
  phv_data_284 = _RAND_284[7:0];
  _RAND_285 = {1{`RANDOM}};
  phv_data_285 = _RAND_285[7:0];
  _RAND_286 = {1{`RANDOM}};
  phv_data_286 = _RAND_286[7:0];
  _RAND_287 = {1{`RANDOM}};
  phv_data_287 = _RAND_287[7:0];
  _RAND_288 = {1{`RANDOM}};
  phv_data_288 = _RAND_288[7:0];
  _RAND_289 = {1{`RANDOM}};
  phv_data_289 = _RAND_289[7:0];
  _RAND_290 = {1{`RANDOM}};
  phv_data_290 = _RAND_290[7:0];
  _RAND_291 = {1{`RANDOM}};
  phv_data_291 = _RAND_291[7:0];
  _RAND_292 = {1{`RANDOM}};
  phv_data_292 = _RAND_292[7:0];
  _RAND_293 = {1{`RANDOM}};
  phv_data_293 = _RAND_293[7:0];
  _RAND_294 = {1{`RANDOM}};
  phv_data_294 = _RAND_294[7:0];
  _RAND_295 = {1{`RANDOM}};
  phv_data_295 = _RAND_295[7:0];
  _RAND_296 = {1{`RANDOM}};
  phv_data_296 = _RAND_296[7:0];
  _RAND_297 = {1{`RANDOM}};
  phv_data_297 = _RAND_297[7:0];
  _RAND_298 = {1{`RANDOM}};
  phv_data_298 = _RAND_298[7:0];
  _RAND_299 = {1{`RANDOM}};
  phv_data_299 = _RAND_299[7:0];
  _RAND_300 = {1{`RANDOM}};
  phv_data_300 = _RAND_300[7:0];
  _RAND_301 = {1{`RANDOM}};
  phv_data_301 = _RAND_301[7:0];
  _RAND_302 = {1{`RANDOM}};
  phv_data_302 = _RAND_302[7:0];
  _RAND_303 = {1{`RANDOM}};
  phv_data_303 = _RAND_303[7:0];
  _RAND_304 = {1{`RANDOM}};
  phv_data_304 = _RAND_304[7:0];
  _RAND_305 = {1{`RANDOM}};
  phv_data_305 = _RAND_305[7:0];
  _RAND_306 = {1{`RANDOM}};
  phv_data_306 = _RAND_306[7:0];
  _RAND_307 = {1{`RANDOM}};
  phv_data_307 = _RAND_307[7:0];
  _RAND_308 = {1{`RANDOM}};
  phv_data_308 = _RAND_308[7:0];
  _RAND_309 = {1{`RANDOM}};
  phv_data_309 = _RAND_309[7:0];
  _RAND_310 = {1{`RANDOM}};
  phv_data_310 = _RAND_310[7:0];
  _RAND_311 = {1{`RANDOM}};
  phv_data_311 = _RAND_311[7:0];
  _RAND_312 = {1{`RANDOM}};
  phv_data_312 = _RAND_312[7:0];
  _RAND_313 = {1{`RANDOM}};
  phv_data_313 = _RAND_313[7:0];
  _RAND_314 = {1{`RANDOM}};
  phv_data_314 = _RAND_314[7:0];
  _RAND_315 = {1{`RANDOM}};
  phv_data_315 = _RAND_315[7:0];
  _RAND_316 = {1{`RANDOM}};
  phv_data_316 = _RAND_316[7:0];
  _RAND_317 = {1{`RANDOM}};
  phv_data_317 = _RAND_317[7:0];
  _RAND_318 = {1{`RANDOM}};
  phv_data_318 = _RAND_318[7:0];
  _RAND_319 = {1{`RANDOM}};
  phv_data_319 = _RAND_319[7:0];
  _RAND_320 = {1{`RANDOM}};
  phv_data_320 = _RAND_320[7:0];
  _RAND_321 = {1{`RANDOM}};
  phv_data_321 = _RAND_321[7:0];
  _RAND_322 = {1{`RANDOM}};
  phv_data_322 = _RAND_322[7:0];
  _RAND_323 = {1{`RANDOM}};
  phv_data_323 = _RAND_323[7:0];
  _RAND_324 = {1{`RANDOM}};
  phv_data_324 = _RAND_324[7:0];
  _RAND_325 = {1{`RANDOM}};
  phv_data_325 = _RAND_325[7:0];
  _RAND_326 = {1{`RANDOM}};
  phv_data_326 = _RAND_326[7:0];
  _RAND_327 = {1{`RANDOM}};
  phv_data_327 = _RAND_327[7:0];
  _RAND_328 = {1{`RANDOM}};
  phv_data_328 = _RAND_328[7:0];
  _RAND_329 = {1{`RANDOM}};
  phv_data_329 = _RAND_329[7:0];
  _RAND_330 = {1{`RANDOM}};
  phv_data_330 = _RAND_330[7:0];
  _RAND_331 = {1{`RANDOM}};
  phv_data_331 = _RAND_331[7:0];
  _RAND_332 = {1{`RANDOM}};
  phv_data_332 = _RAND_332[7:0];
  _RAND_333 = {1{`RANDOM}};
  phv_data_333 = _RAND_333[7:0];
  _RAND_334 = {1{`RANDOM}};
  phv_data_334 = _RAND_334[7:0];
  _RAND_335 = {1{`RANDOM}};
  phv_data_335 = _RAND_335[7:0];
  _RAND_336 = {1{`RANDOM}};
  phv_data_336 = _RAND_336[7:0];
  _RAND_337 = {1{`RANDOM}};
  phv_data_337 = _RAND_337[7:0];
  _RAND_338 = {1{`RANDOM}};
  phv_data_338 = _RAND_338[7:0];
  _RAND_339 = {1{`RANDOM}};
  phv_data_339 = _RAND_339[7:0];
  _RAND_340 = {1{`RANDOM}};
  phv_data_340 = _RAND_340[7:0];
  _RAND_341 = {1{`RANDOM}};
  phv_data_341 = _RAND_341[7:0];
  _RAND_342 = {1{`RANDOM}};
  phv_data_342 = _RAND_342[7:0];
  _RAND_343 = {1{`RANDOM}};
  phv_data_343 = _RAND_343[7:0];
  _RAND_344 = {1{`RANDOM}};
  phv_data_344 = _RAND_344[7:0];
  _RAND_345 = {1{`RANDOM}};
  phv_data_345 = _RAND_345[7:0];
  _RAND_346 = {1{`RANDOM}};
  phv_data_346 = _RAND_346[7:0];
  _RAND_347 = {1{`RANDOM}};
  phv_data_347 = _RAND_347[7:0];
  _RAND_348 = {1{`RANDOM}};
  phv_data_348 = _RAND_348[7:0];
  _RAND_349 = {1{`RANDOM}};
  phv_data_349 = _RAND_349[7:0];
  _RAND_350 = {1{`RANDOM}};
  phv_data_350 = _RAND_350[7:0];
  _RAND_351 = {1{`RANDOM}};
  phv_data_351 = _RAND_351[7:0];
  _RAND_352 = {1{`RANDOM}};
  phv_data_352 = _RAND_352[7:0];
  _RAND_353 = {1{`RANDOM}};
  phv_data_353 = _RAND_353[7:0];
  _RAND_354 = {1{`RANDOM}};
  phv_data_354 = _RAND_354[7:0];
  _RAND_355 = {1{`RANDOM}};
  phv_data_355 = _RAND_355[7:0];
  _RAND_356 = {1{`RANDOM}};
  phv_data_356 = _RAND_356[7:0];
  _RAND_357 = {1{`RANDOM}};
  phv_data_357 = _RAND_357[7:0];
  _RAND_358 = {1{`RANDOM}};
  phv_data_358 = _RAND_358[7:0];
  _RAND_359 = {1{`RANDOM}};
  phv_data_359 = _RAND_359[7:0];
  _RAND_360 = {1{`RANDOM}};
  phv_data_360 = _RAND_360[7:0];
  _RAND_361 = {1{`RANDOM}};
  phv_data_361 = _RAND_361[7:0];
  _RAND_362 = {1{`RANDOM}};
  phv_data_362 = _RAND_362[7:0];
  _RAND_363 = {1{`RANDOM}};
  phv_data_363 = _RAND_363[7:0];
  _RAND_364 = {1{`RANDOM}};
  phv_data_364 = _RAND_364[7:0];
  _RAND_365 = {1{`RANDOM}};
  phv_data_365 = _RAND_365[7:0];
  _RAND_366 = {1{`RANDOM}};
  phv_data_366 = _RAND_366[7:0];
  _RAND_367 = {1{`RANDOM}};
  phv_data_367 = _RAND_367[7:0];
  _RAND_368 = {1{`RANDOM}};
  phv_data_368 = _RAND_368[7:0];
  _RAND_369 = {1{`RANDOM}};
  phv_data_369 = _RAND_369[7:0];
  _RAND_370 = {1{`RANDOM}};
  phv_data_370 = _RAND_370[7:0];
  _RAND_371 = {1{`RANDOM}};
  phv_data_371 = _RAND_371[7:0];
  _RAND_372 = {1{`RANDOM}};
  phv_data_372 = _RAND_372[7:0];
  _RAND_373 = {1{`RANDOM}};
  phv_data_373 = _RAND_373[7:0];
  _RAND_374 = {1{`RANDOM}};
  phv_data_374 = _RAND_374[7:0];
  _RAND_375 = {1{`RANDOM}};
  phv_data_375 = _RAND_375[7:0];
  _RAND_376 = {1{`RANDOM}};
  phv_data_376 = _RAND_376[7:0];
  _RAND_377 = {1{`RANDOM}};
  phv_data_377 = _RAND_377[7:0];
  _RAND_378 = {1{`RANDOM}};
  phv_data_378 = _RAND_378[7:0];
  _RAND_379 = {1{`RANDOM}};
  phv_data_379 = _RAND_379[7:0];
  _RAND_380 = {1{`RANDOM}};
  phv_data_380 = _RAND_380[7:0];
  _RAND_381 = {1{`RANDOM}};
  phv_data_381 = _RAND_381[7:0];
  _RAND_382 = {1{`RANDOM}};
  phv_data_382 = _RAND_382[7:0];
  _RAND_383 = {1{`RANDOM}};
  phv_data_383 = _RAND_383[7:0];
  _RAND_384 = {1{`RANDOM}};
  phv_data_384 = _RAND_384[7:0];
  _RAND_385 = {1{`RANDOM}};
  phv_data_385 = _RAND_385[7:0];
  _RAND_386 = {1{`RANDOM}};
  phv_data_386 = _RAND_386[7:0];
  _RAND_387 = {1{`RANDOM}};
  phv_data_387 = _RAND_387[7:0];
  _RAND_388 = {1{`RANDOM}};
  phv_data_388 = _RAND_388[7:0];
  _RAND_389 = {1{`RANDOM}};
  phv_data_389 = _RAND_389[7:0];
  _RAND_390 = {1{`RANDOM}};
  phv_data_390 = _RAND_390[7:0];
  _RAND_391 = {1{`RANDOM}};
  phv_data_391 = _RAND_391[7:0];
  _RAND_392 = {1{`RANDOM}};
  phv_data_392 = _RAND_392[7:0];
  _RAND_393 = {1{`RANDOM}};
  phv_data_393 = _RAND_393[7:0];
  _RAND_394 = {1{`RANDOM}};
  phv_data_394 = _RAND_394[7:0];
  _RAND_395 = {1{`RANDOM}};
  phv_data_395 = _RAND_395[7:0];
  _RAND_396 = {1{`RANDOM}};
  phv_data_396 = _RAND_396[7:0];
  _RAND_397 = {1{`RANDOM}};
  phv_data_397 = _RAND_397[7:0];
  _RAND_398 = {1{`RANDOM}};
  phv_data_398 = _RAND_398[7:0];
  _RAND_399 = {1{`RANDOM}};
  phv_data_399 = _RAND_399[7:0];
  _RAND_400 = {1{`RANDOM}};
  phv_data_400 = _RAND_400[7:0];
  _RAND_401 = {1{`RANDOM}};
  phv_data_401 = _RAND_401[7:0];
  _RAND_402 = {1{`RANDOM}};
  phv_data_402 = _RAND_402[7:0];
  _RAND_403 = {1{`RANDOM}};
  phv_data_403 = _RAND_403[7:0];
  _RAND_404 = {1{`RANDOM}};
  phv_data_404 = _RAND_404[7:0];
  _RAND_405 = {1{`RANDOM}};
  phv_data_405 = _RAND_405[7:0];
  _RAND_406 = {1{`RANDOM}};
  phv_data_406 = _RAND_406[7:0];
  _RAND_407 = {1{`RANDOM}};
  phv_data_407 = _RAND_407[7:0];
  _RAND_408 = {1{`RANDOM}};
  phv_data_408 = _RAND_408[7:0];
  _RAND_409 = {1{`RANDOM}};
  phv_data_409 = _RAND_409[7:0];
  _RAND_410 = {1{`RANDOM}};
  phv_data_410 = _RAND_410[7:0];
  _RAND_411 = {1{`RANDOM}};
  phv_data_411 = _RAND_411[7:0];
  _RAND_412 = {1{`RANDOM}};
  phv_data_412 = _RAND_412[7:0];
  _RAND_413 = {1{`RANDOM}};
  phv_data_413 = _RAND_413[7:0];
  _RAND_414 = {1{`RANDOM}};
  phv_data_414 = _RAND_414[7:0];
  _RAND_415 = {1{`RANDOM}};
  phv_data_415 = _RAND_415[7:0];
  _RAND_416 = {1{`RANDOM}};
  phv_data_416 = _RAND_416[7:0];
  _RAND_417 = {1{`RANDOM}};
  phv_data_417 = _RAND_417[7:0];
  _RAND_418 = {1{`RANDOM}};
  phv_data_418 = _RAND_418[7:0];
  _RAND_419 = {1{`RANDOM}};
  phv_data_419 = _RAND_419[7:0];
  _RAND_420 = {1{`RANDOM}};
  phv_data_420 = _RAND_420[7:0];
  _RAND_421 = {1{`RANDOM}};
  phv_data_421 = _RAND_421[7:0];
  _RAND_422 = {1{`RANDOM}};
  phv_data_422 = _RAND_422[7:0];
  _RAND_423 = {1{`RANDOM}};
  phv_data_423 = _RAND_423[7:0];
  _RAND_424 = {1{`RANDOM}};
  phv_data_424 = _RAND_424[7:0];
  _RAND_425 = {1{`RANDOM}};
  phv_data_425 = _RAND_425[7:0];
  _RAND_426 = {1{`RANDOM}};
  phv_data_426 = _RAND_426[7:0];
  _RAND_427 = {1{`RANDOM}};
  phv_data_427 = _RAND_427[7:0];
  _RAND_428 = {1{`RANDOM}};
  phv_data_428 = _RAND_428[7:0];
  _RAND_429 = {1{`RANDOM}};
  phv_data_429 = _RAND_429[7:0];
  _RAND_430 = {1{`RANDOM}};
  phv_data_430 = _RAND_430[7:0];
  _RAND_431 = {1{`RANDOM}};
  phv_data_431 = _RAND_431[7:0];
  _RAND_432 = {1{`RANDOM}};
  phv_data_432 = _RAND_432[7:0];
  _RAND_433 = {1{`RANDOM}};
  phv_data_433 = _RAND_433[7:0];
  _RAND_434 = {1{`RANDOM}};
  phv_data_434 = _RAND_434[7:0];
  _RAND_435 = {1{`RANDOM}};
  phv_data_435 = _RAND_435[7:0];
  _RAND_436 = {1{`RANDOM}};
  phv_data_436 = _RAND_436[7:0];
  _RAND_437 = {1{`RANDOM}};
  phv_data_437 = _RAND_437[7:0];
  _RAND_438 = {1{`RANDOM}};
  phv_data_438 = _RAND_438[7:0];
  _RAND_439 = {1{`RANDOM}};
  phv_data_439 = _RAND_439[7:0];
  _RAND_440 = {1{`RANDOM}};
  phv_data_440 = _RAND_440[7:0];
  _RAND_441 = {1{`RANDOM}};
  phv_data_441 = _RAND_441[7:0];
  _RAND_442 = {1{`RANDOM}};
  phv_data_442 = _RAND_442[7:0];
  _RAND_443 = {1{`RANDOM}};
  phv_data_443 = _RAND_443[7:0];
  _RAND_444 = {1{`RANDOM}};
  phv_data_444 = _RAND_444[7:0];
  _RAND_445 = {1{`RANDOM}};
  phv_data_445 = _RAND_445[7:0];
  _RAND_446 = {1{`RANDOM}};
  phv_data_446 = _RAND_446[7:0];
  _RAND_447 = {1{`RANDOM}};
  phv_data_447 = _RAND_447[7:0];
  _RAND_448 = {1{`RANDOM}};
  phv_data_448 = _RAND_448[7:0];
  _RAND_449 = {1{`RANDOM}};
  phv_data_449 = _RAND_449[7:0];
  _RAND_450 = {1{`RANDOM}};
  phv_data_450 = _RAND_450[7:0];
  _RAND_451 = {1{`RANDOM}};
  phv_data_451 = _RAND_451[7:0];
  _RAND_452 = {1{`RANDOM}};
  phv_data_452 = _RAND_452[7:0];
  _RAND_453 = {1{`RANDOM}};
  phv_data_453 = _RAND_453[7:0];
  _RAND_454 = {1{`RANDOM}};
  phv_data_454 = _RAND_454[7:0];
  _RAND_455 = {1{`RANDOM}};
  phv_data_455 = _RAND_455[7:0];
  _RAND_456 = {1{`RANDOM}};
  phv_data_456 = _RAND_456[7:0];
  _RAND_457 = {1{`RANDOM}};
  phv_data_457 = _RAND_457[7:0];
  _RAND_458 = {1{`RANDOM}};
  phv_data_458 = _RAND_458[7:0];
  _RAND_459 = {1{`RANDOM}};
  phv_data_459 = _RAND_459[7:0];
  _RAND_460 = {1{`RANDOM}};
  phv_data_460 = _RAND_460[7:0];
  _RAND_461 = {1{`RANDOM}};
  phv_data_461 = _RAND_461[7:0];
  _RAND_462 = {1{`RANDOM}};
  phv_data_462 = _RAND_462[7:0];
  _RAND_463 = {1{`RANDOM}};
  phv_data_463 = _RAND_463[7:0];
  _RAND_464 = {1{`RANDOM}};
  phv_data_464 = _RAND_464[7:0];
  _RAND_465 = {1{`RANDOM}};
  phv_data_465 = _RAND_465[7:0];
  _RAND_466 = {1{`RANDOM}};
  phv_data_466 = _RAND_466[7:0];
  _RAND_467 = {1{`RANDOM}};
  phv_data_467 = _RAND_467[7:0];
  _RAND_468 = {1{`RANDOM}};
  phv_data_468 = _RAND_468[7:0];
  _RAND_469 = {1{`RANDOM}};
  phv_data_469 = _RAND_469[7:0];
  _RAND_470 = {1{`RANDOM}};
  phv_data_470 = _RAND_470[7:0];
  _RAND_471 = {1{`RANDOM}};
  phv_data_471 = _RAND_471[7:0];
  _RAND_472 = {1{`RANDOM}};
  phv_data_472 = _RAND_472[7:0];
  _RAND_473 = {1{`RANDOM}};
  phv_data_473 = _RAND_473[7:0];
  _RAND_474 = {1{`RANDOM}};
  phv_data_474 = _RAND_474[7:0];
  _RAND_475 = {1{`RANDOM}};
  phv_data_475 = _RAND_475[7:0];
  _RAND_476 = {1{`RANDOM}};
  phv_data_476 = _RAND_476[7:0];
  _RAND_477 = {1{`RANDOM}};
  phv_data_477 = _RAND_477[7:0];
  _RAND_478 = {1{`RANDOM}};
  phv_data_478 = _RAND_478[7:0];
  _RAND_479 = {1{`RANDOM}};
  phv_data_479 = _RAND_479[7:0];
  _RAND_480 = {1{`RANDOM}};
  phv_data_480 = _RAND_480[7:0];
  _RAND_481 = {1{`RANDOM}};
  phv_data_481 = _RAND_481[7:0];
  _RAND_482 = {1{`RANDOM}};
  phv_data_482 = _RAND_482[7:0];
  _RAND_483 = {1{`RANDOM}};
  phv_data_483 = _RAND_483[7:0];
  _RAND_484 = {1{`RANDOM}};
  phv_data_484 = _RAND_484[7:0];
  _RAND_485 = {1{`RANDOM}};
  phv_data_485 = _RAND_485[7:0];
  _RAND_486 = {1{`RANDOM}};
  phv_data_486 = _RAND_486[7:0];
  _RAND_487 = {1{`RANDOM}};
  phv_data_487 = _RAND_487[7:0];
  _RAND_488 = {1{`RANDOM}};
  phv_data_488 = _RAND_488[7:0];
  _RAND_489 = {1{`RANDOM}};
  phv_data_489 = _RAND_489[7:0];
  _RAND_490 = {1{`RANDOM}};
  phv_data_490 = _RAND_490[7:0];
  _RAND_491 = {1{`RANDOM}};
  phv_data_491 = _RAND_491[7:0];
  _RAND_492 = {1{`RANDOM}};
  phv_data_492 = _RAND_492[7:0];
  _RAND_493 = {1{`RANDOM}};
  phv_data_493 = _RAND_493[7:0];
  _RAND_494 = {1{`RANDOM}};
  phv_data_494 = _RAND_494[7:0];
  _RAND_495 = {1{`RANDOM}};
  phv_data_495 = _RAND_495[7:0];
  _RAND_496 = {1{`RANDOM}};
  phv_data_496 = _RAND_496[7:0];
  _RAND_497 = {1{`RANDOM}};
  phv_data_497 = _RAND_497[7:0];
  _RAND_498 = {1{`RANDOM}};
  phv_data_498 = _RAND_498[7:0];
  _RAND_499 = {1{`RANDOM}};
  phv_data_499 = _RAND_499[7:0];
  _RAND_500 = {1{`RANDOM}};
  phv_data_500 = _RAND_500[7:0];
  _RAND_501 = {1{`RANDOM}};
  phv_data_501 = _RAND_501[7:0];
  _RAND_502 = {1{`RANDOM}};
  phv_data_502 = _RAND_502[7:0];
  _RAND_503 = {1{`RANDOM}};
  phv_data_503 = _RAND_503[7:0];
  _RAND_504 = {1{`RANDOM}};
  phv_data_504 = _RAND_504[7:0];
  _RAND_505 = {1{`RANDOM}};
  phv_data_505 = _RAND_505[7:0];
  _RAND_506 = {1{`RANDOM}};
  phv_data_506 = _RAND_506[7:0];
  _RAND_507 = {1{`RANDOM}};
  phv_data_507 = _RAND_507[7:0];
  _RAND_508 = {1{`RANDOM}};
  phv_data_508 = _RAND_508[7:0];
  _RAND_509 = {1{`RANDOM}};
  phv_data_509 = _RAND_509[7:0];
  _RAND_510 = {1{`RANDOM}};
  phv_data_510 = _RAND_510[7:0];
  _RAND_511 = {1{`RANDOM}};
  phv_data_511 = _RAND_511[7:0];
  _RAND_512 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_512[3:0];
  _RAND_513 = {1{`RANDOM}};
  phv_next_config_id = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  args_0 = _RAND_514[7:0];
  _RAND_515 = {1{`RANDOM}};
  args_1 = _RAND_515[7:0];
  _RAND_516 = {1{`RANDOM}};
  args_2 = _RAND_516[7:0];
  _RAND_517 = {1{`RANDOM}};
  args_3 = _RAND_517[7:0];
  _RAND_518 = {1{`RANDOM}};
  args_4 = _RAND_518[7:0];
  _RAND_519 = {1{`RANDOM}};
  args_5 = _RAND_519[7:0];
  _RAND_520 = {1{`RANDOM}};
  args_6 = _RAND_520[7:0];
  _RAND_521 = {1{`RANDOM}};
  vliw_0 = _RAND_521[17:0];
  _RAND_522 = {1{`RANDOM}};
  vliw_1 = _RAND_522[17:0];
  _RAND_523 = {1{`RANDOM}};
  vliw_2 = _RAND_523[17:0];
  _RAND_524 = {1{`RANDOM}};
  vliw_3 = _RAND_524[17:0];
  _RAND_525 = {1{`RANDOM}};
  vliw_4 = _RAND_525[17:0];
  _RAND_526 = {1{`RANDOM}};
  vliw_5 = _RAND_526[17:0];
  _RAND_527 = {1{`RANDOM}};
  vliw_6 = _RAND_527[17:0];
  _RAND_528 = {1{`RANDOM}};
  vliw_7 = _RAND_528[17:0];
  _RAND_529 = {1{`RANDOM}};
  vliw_8 = _RAND_529[17:0];
  _RAND_530 = {1{`RANDOM}};
  vliw_9 = _RAND_530[17:0];
  _RAND_531 = {1{`RANDOM}};
  vliw_10 = _RAND_531[17:0];
  _RAND_532 = {1{`RANDOM}};
  vliw_11 = _RAND_532[17:0];
  _RAND_533 = {1{`RANDOM}};
  vliw_12 = _RAND_533[17:0];
  _RAND_534 = {1{`RANDOM}};
  vliw_13 = _RAND_534[17:0];
  _RAND_535 = {1{`RANDOM}};
  vliw_14 = _RAND_535[17:0];
  _RAND_536 = {1{`RANDOM}};
  vliw_15 = _RAND_536[17:0];
  _RAND_537 = {1{`RANDOM}};
  vliw_16 = _RAND_537[17:0];
  _RAND_538 = {1{`RANDOM}};
  vliw_17 = _RAND_538[17:0];
  _RAND_539 = {1{`RANDOM}};
  vliw_18 = _RAND_539[17:0];
  _RAND_540 = {1{`RANDOM}};
  vliw_19 = _RAND_540[17:0];
  _RAND_541 = {1{`RANDOM}};
  vliw_20 = _RAND_541[17:0];
  _RAND_542 = {1{`RANDOM}};
  vliw_21 = _RAND_542[17:0];
  _RAND_543 = {1{`RANDOM}};
  vliw_22 = _RAND_543[17:0];
  _RAND_544 = {1{`RANDOM}};
  vliw_23 = _RAND_544[17:0];
  _RAND_545 = {1{`RANDOM}};
  vliw_24 = _RAND_545[17:0];
  _RAND_546 = {1{`RANDOM}};
  vliw_25 = _RAND_546[17:0];
  _RAND_547 = {1{`RANDOM}};
  vliw_26 = _RAND_547[17:0];
  _RAND_548 = {1{`RANDOM}};
  vliw_27 = _RAND_548[17:0];
  _RAND_549 = {1{`RANDOM}};
  vliw_28 = _RAND_549[17:0];
  _RAND_550 = {1{`RANDOM}};
  vliw_29 = _RAND_550[17:0];
  _RAND_551 = {1{`RANDOM}};
  vliw_30 = _RAND_551[17:0];
  _RAND_552 = {1{`RANDOM}};
  vliw_31 = _RAND_552[17:0];
  _RAND_553 = {1{`RANDOM}};
  vliw_32 = _RAND_553[17:0];
  _RAND_554 = {1{`RANDOM}};
  vliw_33 = _RAND_554[17:0];
  _RAND_555 = {1{`RANDOM}};
  vliw_34 = _RAND_555[17:0];
  _RAND_556 = {1{`RANDOM}};
  vliw_35 = _RAND_556[17:0];
  _RAND_557 = {1{`RANDOM}};
  vliw_36 = _RAND_557[17:0];
  _RAND_558 = {1{`RANDOM}};
  vliw_37 = _RAND_558[17:0];
  _RAND_559 = {1{`RANDOM}};
  vliw_38 = _RAND_559[17:0];
  _RAND_560 = {1{`RANDOM}};
  vliw_39 = _RAND_560[17:0];
  _RAND_561 = {1{`RANDOM}};
  vliw_40 = _RAND_561[17:0];
  _RAND_562 = {1{`RANDOM}};
  vliw_41 = _RAND_562[17:0];
  _RAND_563 = {1{`RANDOM}};
  vliw_42 = _RAND_563[17:0];
  _RAND_564 = {1{`RANDOM}};
  vliw_43 = _RAND_564[17:0];
  _RAND_565 = {1{`RANDOM}};
  vliw_44 = _RAND_565[17:0];
  _RAND_566 = {1{`RANDOM}};
  vliw_45 = _RAND_566[17:0];
  _RAND_567 = {1{`RANDOM}};
  vliw_46 = _RAND_567[17:0];
  _RAND_568 = {1{`RANDOM}};
  vliw_47 = _RAND_568[17:0];
  _RAND_569 = {1{`RANDOM}};
  vliw_48 = _RAND_569[17:0];
  _RAND_570 = {1{`RANDOM}};
  vliw_49 = _RAND_570[17:0];
  _RAND_571 = {1{`RANDOM}};
  vliw_50 = _RAND_571[17:0];
  _RAND_572 = {1{`RANDOM}};
  vliw_51 = _RAND_572[17:0];
  _RAND_573 = {1{`RANDOM}};
  vliw_52 = _RAND_573[17:0];
  _RAND_574 = {1{`RANDOM}};
  vliw_53 = _RAND_574[17:0];
  _RAND_575 = {1{`RANDOM}};
  vliw_54 = _RAND_575[17:0];
  _RAND_576 = {1{`RANDOM}};
  vliw_55 = _RAND_576[17:0];
  _RAND_577 = {1{`RANDOM}};
  vliw_56 = _RAND_577[17:0];
  _RAND_578 = {1{`RANDOM}};
  vliw_57 = _RAND_578[17:0];
  _RAND_579 = {1{`RANDOM}};
  vliw_58 = _RAND_579[17:0];
  _RAND_580 = {1{`RANDOM}};
  vliw_59 = _RAND_580[17:0];
  _RAND_581 = {1{`RANDOM}};
  vliw_60 = _RAND_581[17:0];
  _RAND_582 = {1{`RANDOM}};
  vliw_61 = _RAND_582[17:0];
  _RAND_583 = {1{`RANDOM}};
  vliw_62 = _RAND_583[17:0];
  _RAND_584 = {1{`RANDOM}};
  vliw_63 = _RAND_584[17:0];
  _RAND_585 = {1{`RANDOM}};
  vliw_64 = _RAND_585[17:0];
  _RAND_586 = {1{`RANDOM}};
  vliw_65 = _RAND_586[17:0];
  _RAND_587 = {1{`RANDOM}};
  vliw_66 = _RAND_587[17:0];
  _RAND_588 = {1{`RANDOM}};
  vliw_67 = _RAND_588[17:0];
  _RAND_589 = {1{`RANDOM}};
  vliw_68 = _RAND_589[17:0];
  _RAND_590 = {1{`RANDOM}};
  vliw_69 = _RAND_590[17:0];
  _RAND_591 = {1{`RANDOM}};
  nid = _RAND_591[14:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
